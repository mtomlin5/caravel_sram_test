magic
tech sky130A
magscale 1 2
timestamp 1636725489
<< obsli1 >>
rect 673 901 49099 47345
<< obsm1 >>
rect 14 892 49850 47376
<< metal2 >>
rect 202 49200 258 50000
rect 570 49200 626 50000
rect 1030 49200 1086 50000
rect 1398 49200 1454 50000
rect 1858 49200 1914 50000
rect 2226 49200 2282 50000
rect 2686 49200 2742 50000
rect 3054 49200 3110 50000
rect 3514 49200 3570 50000
rect 3882 49200 3938 50000
rect 4342 49200 4398 50000
rect 4710 49200 4766 50000
rect 5170 49200 5226 50000
rect 5538 49200 5594 50000
rect 5998 49200 6054 50000
rect 6366 49200 6422 50000
rect 6826 49200 6882 50000
rect 7194 49200 7250 50000
rect 7654 49200 7710 50000
rect 8022 49200 8078 50000
rect 8482 49200 8538 50000
rect 8942 49200 8998 50000
rect 9310 49200 9366 50000
rect 9770 49200 9826 50000
rect 10138 49200 10194 50000
rect 10598 49200 10654 50000
rect 10966 49200 11022 50000
rect 11426 49200 11482 50000
rect 11794 49200 11850 50000
rect 12254 49200 12310 50000
rect 12622 49200 12678 50000
rect 13082 49200 13138 50000
rect 13450 49200 13506 50000
rect 13910 49200 13966 50000
rect 14278 49200 14334 50000
rect 14738 49200 14794 50000
rect 15106 49200 15162 50000
rect 15566 49200 15622 50000
rect 15934 49200 15990 50000
rect 16394 49200 16450 50000
rect 16854 49200 16910 50000
rect 17222 49200 17278 50000
rect 17682 49200 17738 50000
rect 18050 49200 18106 50000
rect 18510 49200 18566 50000
rect 18878 49200 18934 50000
rect 19338 49200 19394 50000
rect 19706 49200 19762 50000
rect 20166 49200 20222 50000
rect 20534 49200 20590 50000
rect 20994 49200 21050 50000
rect 21362 49200 21418 50000
rect 21822 49200 21878 50000
rect 22190 49200 22246 50000
rect 22650 49200 22706 50000
rect 23018 49200 23074 50000
rect 23478 49200 23534 50000
rect 23846 49200 23902 50000
rect 24306 49200 24362 50000
rect 24674 49200 24730 50000
rect 25134 49200 25190 50000
rect 25594 49200 25650 50000
rect 25962 49200 26018 50000
rect 26422 49200 26478 50000
rect 26790 49200 26846 50000
rect 27250 49200 27306 50000
rect 27618 49200 27674 50000
rect 28078 49200 28134 50000
rect 28446 49200 28502 50000
rect 28906 49200 28962 50000
rect 29274 49200 29330 50000
rect 29734 49200 29790 50000
rect 30102 49200 30158 50000
rect 30562 49200 30618 50000
rect 30930 49200 30986 50000
rect 31390 49200 31446 50000
rect 31758 49200 31814 50000
rect 32218 49200 32274 50000
rect 32586 49200 32642 50000
rect 33046 49200 33102 50000
rect 33506 49200 33562 50000
rect 33874 49200 33930 50000
rect 34334 49200 34390 50000
rect 34702 49200 34758 50000
rect 35162 49200 35218 50000
rect 35530 49200 35586 50000
rect 35990 49200 36046 50000
rect 36358 49200 36414 50000
rect 36818 49200 36874 50000
rect 37186 49200 37242 50000
rect 37646 49200 37702 50000
rect 38014 49200 38070 50000
rect 38474 49200 38530 50000
rect 38842 49200 38898 50000
rect 39302 49200 39358 50000
rect 39670 49200 39726 50000
rect 40130 49200 40186 50000
rect 40498 49200 40554 50000
rect 40958 49200 41014 50000
rect 41326 49200 41382 50000
rect 41786 49200 41842 50000
rect 42246 49200 42302 50000
rect 42614 49200 42670 50000
rect 43074 49200 43130 50000
rect 43442 49200 43498 50000
rect 43902 49200 43958 50000
rect 44270 49200 44326 50000
rect 44730 49200 44786 50000
rect 45098 49200 45154 50000
rect 45558 49200 45614 50000
rect 45926 49200 45982 50000
rect 46386 49200 46442 50000
rect 46754 49200 46810 50000
rect 47214 49200 47270 50000
rect 47582 49200 47638 50000
rect 48042 49200 48098 50000
rect 48410 49200 48466 50000
rect 48870 49200 48926 50000
rect 49238 49200 49294 50000
rect 49698 49200 49754 50000
rect 18 0 74 800
rect 110 0 166 800
rect 202 0 258 800
rect 294 0 350 800
rect 386 0 442 800
rect 478 0 534 800
rect 570 0 626 800
rect 662 0 718 800
rect 754 0 810 800
rect 846 0 902 800
rect 938 0 994 800
rect 1030 0 1086 800
rect 1214 0 1270 800
rect 1306 0 1362 800
rect 1398 0 1454 800
rect 1490 0 1546 800
rect 1582 0 1638 800
rect 1674 0 1730 800
rect 1766 0 1822 800
rect 1858 0 1914 800
rect 1950 0 2006 800
rect 2042 0 2098 800
rect 2134 0 2190 800
rect 2226 0 2282 800
rect 2410 0 2466 800
rect 2502 0 2558 800
rect 2594 0 2650 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2870 0 2926 800
rect 2962 0 3018 800
rect 3054 0 3110 800
rect 3146 0 3202 800
rect 3238 0 3294 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3606 0 3662 800
rect 3698 0 3754 800
rect 3790 0 3846 800
rect 3882 0 3938 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4158 0 4214 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4434 0 4490 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4802 0 4858 800
rect 4894 0 4950 800
rect 4986 0 5042 800
rect 5078 0 5134 800
rect 5170 0 5226 800
rect 5262 0 5318 800
rect 5354 0 5410 800
rect 5446 0 5502 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 7010 0 7066 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
<< obsm2 >>
rect 20 49144 146 49745
rect 314 49144 514 49745
rect 682 49144 974 49745
rect 1142 49144 1342 49745
rect 1510 49144 1802 49745
rect 1970 49144 2170 49745
rect 2338 49144 2630 49745
rect 2798 49144 2998 49745
rect 3166 49144 3458 49745
rect 3626 49144 3826 49745
rect 3994 49144 4286 49745
rect 4454 49144 4654 49745
rect 4822 49144 5114 49745
rect 5282 49144 5482 49745
rect 5650 49144 5942 49745
rect 6110 49144 6310 49745
rect 6478 49144 6770 49745
rect 6938 49144 7138 49745
rect 7306 49144 7598 49745
rect 7766 49144 7966 49745
rect 8134 49144 8426 49745
rect 8594 49144 8886 49745
rect 9054 49144 9254 49745
rect 9422 49144 9714 49745
rect 9882 49144 10082 49745
rect 10250 49144 10542 49745
rect 10710 49144 10910 49745
rect 11078 49144 11370 49745
rect 11538 49144 11738 49745
rect 11906 49144 12198 49745
rect 12366 49144 12566 49745
rect 12734 49144 13026 49745
rect 13194 49144 13394 49745
rect 13562 49144 13854 49745
rect 14022 49144 14222 49745
rect 14390 49144 14682 49745
rect 14850 49144 15050 49745
rect 15218 49144 15510 49745
rect 15678 49144 15878 49745
rect 16046 49144 16338 49745
rect 16506 49144 16798 49745
rect 16966 49144 17166 49745
rect 17334 49144 17626 49745
rect 17794 49144 17994 49745
rect 18162 49144 18454 49745
rect 18622 49144 18822 49745
rect 18990 49144 19282 49745
rect 19450 49144 19650 49745
rect 19818 49144 20110 49745
rect 20278 49144 20478 49745
rect 20646 49144 20938 49745
rect 21106 49144 21306 49745
rect 21474 49144 21766 49745
rect 21934 49144 22134 49745
rect 22302 49144 22594 49745
rect 22762 49144 22962 49745
rect 23130 49144 23422 49745
rect 23590 49144 23790 49745
rect 23958 49144 24250 49745
rect 24418 49144 24618 49745
rect 24786 49144 25078 49745
rect 25246 49144 25538 49745
rect 25706 49144 25906 49745
rect 26074 49144 26366 49745
rect 26534 49144 26734 49745
rect 26902 49144 27194 49745
rect 27362 49144 27562 49745
rect 27730 49144 28022 49745
rect 28190 49144 28390 49745
rect 28558 49144 28850 49745
rect 29018 49144 29218 49745
rect 29386 49144 29678 49745
rect 29846 49144 30046 49745
rect 30214 49144 30506 49745
rect 30674 49144 30874 49745
rect 31042 49144 31334 49745
rect 31502 49144 31702 49745
rect 31870 49144 32162 49745
rect 32330 49144 32530 49745
rect 32698 49144 32990 49745
rect 33158 49144 33450 49745
rect 33618 49144 33818 49745
rect 33986 49144 34278 49745
rect 34446 49144 34646 49745
rect 34814 49144 35106 49745
rect 35274 49144 35474 49745
rect 35642 49144 35934 49745
rect 36102 49144 36302 49745
rect 36470 49144 36762 49745
rect 36930 49144 37130 49745
rect 37298 49144 37590 49745
rect 37758 49144 37958 49745
rect 38126 49144 38418 49745
rect 38586 49144 38786 49745
rect 38954 49144 39246 49745
rect 39414 49144 39614 49745
rect 39782 49144 40074 49745
rect 40242 49144 40442 49745
rect 40610 49144 40902 49745
rect 41070 49144 41270 49745
rect 41438 49144 41730 49745
rect 41898 49144 42190 49745
rect 42358 49144 42558 49745
rect 42726 49144 43018 49745
rect 43186 49144 43386 49745
rect 43554 49144 43846 49745
rect 44014 49144 44214 49745
rect 44382 49144 44674 49745
rect 44842 49144 45042 49745
rect 45210 49144 45502 49745
rect 45670 49144 45870 49745
rect 46038 49144 46330 49745
rect 46498 49144 46698 49745
rect 46866 49144 47158 49745
rect 47326 49144 47526 49745
rect 47694 49144 47986 49745
rect 48154 49144 48354 49745
rect 48522 49144 48814 49745
rect 48982 49144 49182 49745
rect 49350 49144 49642 49745
rect 49810 49144 49844 49745
rect 20 856 49844 49144
rect 1142 303 1158 856
rect 2338 303 2354 856
rect 3442 303 3458 856
rect 4638 303 4654 856
rect 5834 303 5850 856
rect 6938 303 6954 856
rect 8134 303 8150 856
rect 9330 303 9346 856
rect 10434 303 10450 856
rect 11630 303 11646 856
rect 12734 303 12750 856
rect 13930 303 13946 856
rect 15126 303 15142 856
rect 16230 303 16246 856
rect 17426 303 17442 856
rect 18622 303 18638 856
rect 19726 303 19742 856
rect 20922 303 20938 856
rect 22026 303 22042 856
rect 23222 303 23238 856
rect 24418 303 24434 856
rect 25522 303 25538 856
rect 26718 303 26734 856
rect 27914 303 27930 856
rect 29018 303 29034 856
rect 30214 303 30230 856
rect 31318 303 31334 856
rect 32514 303 32530 856
rect 33710 303 33726 856
rect 34814 303 34830 856
rect 36010 303 36026 856
rect 37206 303 37222 856
rect 38310 303 38326 856
rect 39506 303 39522 856
rect 40610 303 40626 856
rect 41806 303 41822 856
rect 43002 303 43018 856
rect 44106 303 44122 856
rect 45302 303 45318 856
rect 46498 303 46514 856
rect 47602 303 47618 856
rect 48798 303 48814 856
<< metal3 >>
rect 49200 49648 50000 49768
rect 49200 48968 50000 49088
rect 49200 48288 50000 48408
rect 49200 47608 50000 47728
rect 0 47200 800 47320
rect 49200 47064 50000 47184
rect 49200 46384 50000 46504
rect 49200 45704 50000 45824
rect 49200 45024 50000 45144
rect 49200 44344 50000 44464
rect 49200 43800 50000 43920
rect 49200 43120 50000 43240
rect 49200 42440 50000 42560
rect 0 41624 800 41744
rect 49200 41760 50000 41880
rect 49200 41216 50000 41336
rect 49200 40536 50000 40656
rect 49200 39856 50000 39976
rect 49200 39176 50000 39296
rect 49200 38496 50000 38616
rect 49200 37952 50000 38072
rect 49200 37272 50000 37392
rect 49200 36592 50000 36712
rect 0 36048 800 36168
rect 49200 35912 50000 36032
rect 49200 35368 50000 35488
rect 49200 34688 50000 34808
rect 49200 34008 50000 34128
rect 49200 33328 50000 33448
rect 49200 32648 50000 32768
rect 49200 32104 50000 32224
rect 49200 31424 50000 31544
rect 49200 30744 50000 30864
rect 0 30472 800 30592
rect 49200 30064 50000 30184
rect 49200 29520 50000 29640
rect 49200 28840 50000 28960
rect 49200 28160 50000 28280
rect 49200 27480 50000 27600
rect 49200 26800 50000 26920
rect 49200 26256 50000 26376
rect 49200 25576 50000 25696
rect 0 24896 800 25016
rect 49200 24896 50000 25016
rect 49200 24216 50000 24336
rect 49200 23672 50000 23792
rect 49200 22992 50000 23112
rect 49200 22312 50000 22432
rect 49200 21632 50000 21752
rect 49200 20952 50000 21072
rect 49200 20408 50000 20528
rect 49200 19728 50000 19848
rect 0 19320 800 19440
rect 49200 19048 50000 19168
rect 49200 18368 50000 18488
rect 49200 17824 50000 17944
rect 49200 17144 50000 17264
rect 49200 16464 50000 16584
rect 49200 15784 50000 15904
rect 49200 15104 50000 15224
rect 49200 14560 50000 14680
rect 0 13744 800 13864
rect 49200 13880 50000 14000
rect 49200 13200 50000 13320
rect 49200 12520 50000 12640
rect 49200 11976 50000 12096
rect 49200 11296 50000 11416
rect 49200 10616 50000 10736
rect 49200 9936 50000 10056
rect 49200 9256 50000 9376
rect 49200 8712 50000 8832
rect 0 8168 800 8288
rect 49200 8032 50000 8152
rect 49200 7352 50000 7472
rect 49200 6672 50000 6792
rect 49200 6128 50000 6248
rect 49200 5448 50000 5568
rect 49200 4768 50000 4888
rect 49200 4088 50000 4208
rect 49200 3408 50000 3528
rect 0 2728 800 2848
rect 49200 2864 50000 2984
rect 49200 2184 50000 2304
rect 49200 1504 50000 1624
rect 49200 824 50000 944
rect 49200 280 50000 400
<< obsm3 >>
rect 800 49568 49120 49741
rect 800 49168 49200 49568
rect 800 48888 49120 49168
rect 800 48488 49200 48888
rect 800 48208 49120 48488
rect 800 47808 49200 48208
rect 800 47528 49120 47808
rect 800 47400 49200 47528
rect 880 47264 49200 47400
rect 880 47120 49120 47264
rect 800 46984 49120 47120
rect 800 46584 49200 46984
rect 800 46304 49120 46584
rect 800 45904 49200 46304
rect 800 45624 49120 45904
rect 800 45224 49200 45624
rect 800 44944 49120 45224
rect 800 44544 49200 44944
rect 800 44264 49120 44544
rect 800 44000 49200 44264
rect 800 43720 49120 44000
rect 800 43320 49200 43720
rect 800 43040 49120 43320
rect 800 42640 49200 43040
rect 800 42360 49120 42640
rect 800 41960 49200 42360
rect 800 41824 49120 41960
rect 880 41680 49120 41824
rect 880 41544 49200 41680
rect 800 41416 49200 41544
rect 800 41136 49120 41416
rect 800 40736 49200 41136
rect 800 40456 49120 40736
rect 800 40056 49200 40456
rect 800 39776 49120 40056
rect 800 39376 49200 39776
rect 800 39096 49120 39376
rect 800 38696 49200 39096
rect 800 38416 49120 38696
rect 800 38152 49200 38416
rect 800 37872 49120 38152
rect 800 37472 49200 37872
rect 800 37192 49120 37472
rect 800 36792 49200 37192
rect 800 36512 49120 36792
rect 800 36248 49200 36512
rect 880 36112 49200 36248
rect 880 35968 49120 36112
rect 800 35832 49120 35968
rect 800 35568 49200 35832
rect 800 35288 49120 35568
rect 800 34888 49200 35288
rect 800 34608 49120 34888
rect 800 34208 49200 34608
rect 800 33928 49120 34208
rect 800 33528 49200 33928
rect 800 33248 49120 33528
rect 800 32848 49200 33248
rect 800 32568 49120 32848
rect 800 32304 49200 32568
rect 800 32024 49120 32304
rect 800 31624 49200 32024
rect 800 31344 49120 31624
rect 800 30944 49200 31344
rect 800 30672 49120 30944
rect 880 30664 49120 30672
rect 880 30392 49200 30664
rect 800 30264 49200 30392
rect 800 29984 49120 30264
rect 800 29720 49200 29984
rect 800 29440 49120 29720
rect 800 29040 49200 29440
rect 800 28760 49120 29040
rect 800 28360 49200 28760
rect 800 28080 49120 28360
rect 800 27680 49200 28080
rect 800 27400 49120 27680
rect 800 27000 49200 27400
rect 800 26720 49120 27000
rect 800 26456 49200 26720
rect 800 26176 49120 26456
rect 800 25776 49200 26176
rect 800 25496 49120 25776
rect 800 25096 49200 25496
rect 880 24816 49120 25096
rect 800 24416 49200 24816
rect 800 24136 49120 24416
rect 800 23872 49200 24136
rect 800 23592 49120 23872
rect 800 23192 49200 23592
rect 800 22912 49120 23192
rect 800 22512 49200 22912
rect 800 22232 49120 22512
rect 800 21832 49200 22232
rect 800 21552 49120 21832
rect 800 21152 49200 21552
rect 800 20872 49120 21152
rect 800 20608 49200 20872
rect 800 20328 49120 20608
rect 800 19928 49200 20328
rect 800 19648 49120 19928
rect 800 19520 49200 19648
rect 880 19248 49200 19520
rect 880 19240 49120 19248
rect 800 18968 49120 19240
rect 800 18568 49200 18968
rect 800 18288 49120 18568
rect 800 18024 49200 18288
rect 800 17744 49120 18024
rect 800 17344 49200 17744
rect 800 17064 49120 17344
rect 800 16664 49200 17064
rect 800 16384 49120 16664
rect 800 15984 49200 16384
rect 800 15704 49120 15984
rect 800 15304 49200 15704
rect 800 15024 49120 15304
rect 800 14760 49200 15024
rect 800 14480 49120 14760
rect 800 14080 49200 14480
rect 800 13944 49120 14080
rect 880 13800 49120 13944
rect 880 13664 49200 13800
rect 800 13400 49200 13664
rect 800 13120 49120 13400
rect 800 12720 49200 13120
rect 800 12440 49120 12720
rect 800 12176 49200 12440
rect 800 11896 49120 12176
rect 800 11496 49200 11896
rect 800 11216 49120 11496
rect 800 10816 49200 11216
rect 800 10536 49120 10816
rect 800 10136 49200 10536
rect 800 9856 49120 10136
rect 800 9456 49200 9856
rect 800 9176 49120 9456
rect 800 8912 49200 9176
rect 800 8632 49120 8912
rect 800 8368 49200 8632
rect 880 8232 49200 8368
rect 880 8088 49120 8232
rect 800 7952 49120 8088
rect 800 7552 49200 7952
rect 800 7272 49120 7552
rect 800 6872 49200 7272
rect 800 6592 49120 6872
rect 800 6328 49200 6592
rect 800 6048 49120 6328
rect 800 5648 49200 6048
rect 800 5368 49120 5648
rect 800 4968 49200 5368
rect 800 4688 49120 4968
rect 800 4288 49200 4688
rect 800 4008 49120 4288
rect 800 3608 49200 4008
rect 800 3328 49120 3608
rect 800 3064 49200 3328
rect 800 2928 49120 3064
rect 880 2784 49120 2928
rect 880 2648 49200 2784
rect 800 2384 49200 2648
rect 800 2104 49120 2384
rect 800 1704 49200 2104
rect 800 1424 49120 1704
rect 800 1024 49200 1424
rect 800 744 49120 1024
rect 800 480 49200 744
rect 800 307 49120 480
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
<< obsm4 >>
rect 1163 2048 4128 42533
rect 4608 2048 19488 42533
rect 19968 2048 34848 42533
rect 35328 2048 48149 42533
rect 1163 851 48149 2048
<< labels >>
rlabel metal3 s 49200 41760 50000 41880 6 csb0
port 1 nsew signal output
rlabel metal3 s 49200 43120 50000 43240 6 csb1
port 2 nsew signal output
rlabel metal3 s 49200 43800 50000 43920 6 din0[0]
port 3 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 din0[10]
port 4 nsew signal output
rlabel metal2 s 48410 49200 48466 50000 6 din0[11]
port 5 nsew signal output
rlabel metal3 s 49200 45704 50000 45824 6 din0[12]
port 6 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 din0[13]
port 7 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 din0[14]
port 8 nsew signal output
rlabel metal3 s 49200 46384 50000 46504 6 din0[15]
port 9 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 din0[16]
port 10 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 din0[17]
port 11 nsew signal output
rlabel metal3 s 49200 47064 50000 47184 6 din0[18]
port 12 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 din0[19]
port 13 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 din0[1]
port 14 nsew signal output
rlabel metal2 s 48870 49200 48926 50000 6 din0[20]
port 15 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 din0[21]
port 16 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 din0[22]
port 17 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 din0[23]
port 18 nsew signal output
rlabel metal2 s 49238 49200 49294 50000 6 din0[24]
port 19 nsew signal output
rlabel metal2 s 49698 49200 49754 50000 6 din0[25]
port 20 nsew signal output
rlabel metal3 s 49200 47608 50000 47728 6 din0[26]
port 21 nsew signal output
rlabel metal3 s 49200 48288 50000 48408 6 din0[27]
port 22 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 din0[28]
port 23 nsew signal output
rlabel metal3 s 49200 48968 50000 49088 6 din0[29]
port 24 nsew signal output
rlabel metal2 s 47582 49200 47638 50000 6 din0[2]
port 25 nsew signal output
rlabel metal3 s 49200 49648 50000 49768 6 din0[30]
port 26 nsew signal output
rlabel metal3 s 0 47200 800 47320 6 din0[31]
port 27 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 din0[3]
port 28 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 din0[4]
port 29 nsew signal output
rlabel metal3 s 49200 44344 50000 44464 6 din0[5]
port 30 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 din0[6]
port 31 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 din0[7]
port 32 nsew signal output
rlabel metal3 s 49200 45024 50000 45144 6 din0[8]
port 33 nsew signal output
rlabel metal2 s 48042 49200 48098 50000 6 din0[9]
port 34 nsew signal output
rlabel metal3 s 49200 280 50000 400 6 dout0[0]
port 35 nsew signal input
rlabel metal3 s 49200 6672 50000 6792 6 dout0[10]
port 36 nsew signal input
rlabel metal3 s 49200 7352 50000 7472 6 dout0[11]
port 37 nsew signal input
rlabel metal3 s 49200 8032 50000 8152 6 dout0[12]
port 38 nsew signal input
rlabel metal3 s 49200 8712 50000 8832 6 dout0[13]
port 39 nsew signal input
rlabel metal3 s 49200 9256 50000 9376 6 dout0[14]
port 40 nsew signal input
rlabel metal3 s 49200 9936 50000 10056 6 dout0[15]
port 41 nsew signal input
rlabel metal3 s 49200 10616 50000 10736 6 dout0[16]
port 42 nsew signal input
rlabel metal3 s 49200 11296 50000 11416 6 dout0[17]
port 43 nsew signal input
rlabel metal3 s 49200 11976 50000 12096 6 dout0[18]
port 44 nsew signal input
rlabel metal3 s 49200 12520 50000 12640 6 dout0[19]
port 45 nsew signal input
rlabel metal3 s 49200 824 50000 944 6 dout0[1]
port 46 nsew signal input
rlabel metal3 s 49200 13200 50000 13320 6 dout0[20]
port 47 nsew signal input
rlabel metal3 s 49200 13880 50000 14000 6 dout0[21]
port 48 nsew signal input
rlabel metal3 s 49200 14560 50000 14680 6 dout0[22]
port 49 nsew signal input
rlabel metal3 s 49200 15104 50000 15224 6 dout0[23]
port 50 nsew signal input
rlabel metal3 s 49200 15784 50000 15904 6 dout0[24]
port 51 nsew signal input
rlabel metal3 s 49200 16464 50000 16584 6 dout0[25]
port 52 nsew signal input
rlabel metal3 s 49200 17144 50000 17264 6 dout0[26]
port 53 nsew signal input
rlabel metal3 s 49200 17824 50000 17944 6 dout0[27]
port 54 nsew signal input
rlabel metal3 s 49200 18368 50000 18488 6 dout0[28]
port 55 nsew signal input
rlabel metal3 s 49200 19048 50000 19168 6 dout0[29]
port 56 nsew signal input
rlabel metal3 s 49200 1504 50000 1624 6 dout0[2]
port 57 nsew signal input
rlabel metal3 s 49200 19728 50000 19848 6 dout0[30]
port 58 nsew signal input
rlabel metal3 s 49200 20408 50000 20528 6 dout0[31]
port 59 nsew signal input
rlabel metal3 s 49200 2184 50000 2304 6 dout0[3]
port 60 nsew signal input
rlabel metal3 s 49200 2864 50000 2984 6 dout0[4]
port 61 nsew signal input
rlabel metal3 s 49200 3408 50000 3528 6 dout0[5]
port 62 nsew signal input
rlabel metal3 s 49200 4088 50000 4208 6 dout0[6]
port 63 nsew signal input
rlabel metal3 s 49200 4768 50000 4888 6 dout0[7]
port 64 nsew signal input
rlabel metal3 s 49200 5448 50000 5568 6 dout0[8]
port 65 nsew signal input
rlabel metal3 s 49200 6128 50000 6248 6 dout0[9]
port 66 nsew signal input
rlabel metal3 s 49200 20952 50000 21072 6 dout1[0]
port 67 nsew signal input
rlabel metal3 s 49200 27480 50000 27600 6 dout1[10]
port 68 nsew signal input
rlabel metal3 s 49200 28160 50000 28280 6 dout1[11]
port 69 nsew signal input
rlabel metal3 s 49200 28840 50000 28960 6 dout1[12]
port 70 nsew signal input
rlabel metal3 s 49200 29520 50000 29640 6 dout1[13]
port 71 nsew signal input
rlabel metal3 s 49200 30064 50000 30184 6 dout1[14]
port 72 nsew signal input
rlabel metal3 s 49200 30744 50000 30864 6 dout1[15]
port 73 nsew signal input
rlabel metal3 s 49200 31424 50000 31544 6 dout1[16]
port 74 nsew signal input
rlabel metal3 s 49200 32104 50000 32224 6 dout1[17]
port 75 nsew signal input
rlabel metal3 s 49200 32648 50000 32768 6 dout1[18]
port 76 nsew signal input
rlabel metal3 s 49200 33328 50000 33448 6 dout1[19]
port 77 nsew signal input
rlabel metal3 s 49200 21632 50000 21752 6 dout1[1]
port 78 nsew signal input
rlabel metal3 s 49200 34008 50000 34128 6 dout1[20]
port 79 nsew signal input
rlabel metal3 s 49200 34688 50000 34808 6 dout1[21]
port 80 nsew signal input
rlabel metal3 s 49200 35368 50000 35488 6 dout1[22]
port 81 nsew signal input
rlabel metal3 s 49200 35912 50000 36032 6 dout1[23]
port 82 nsew signal input
rlabel metal3 s 49200 36592 50000 36712 6 dout1[24]
port 83 nsew signal input
rlabel metal3 s 49200 37272 50000 37392 6 dout1[25]
port 84 nsew signal input
rlabel metal3 s 49200 37952 50000 38072 6 dout1[26]
port 85 nsew signal input
rlabel metal3 s 49200 38496 50000 38616 6 dout1[27]
port 86 nsew signal input
rlabel metal3 s 49200 39176 50000 39296 6 dout1[28]
port 87 nsew signal input
rlabel metal3 s 49200 39856 50000 39976 6 dout1[29]
port 88 nsew signal input
rlabel metal3 s 49200 22312 50000 22432 6 dout1[2]
port 89 nsew signal input
rlabel metal3 s 49200 40536 50000 40656 6 dout1[30]
port 90 nsew signal input
rlabel metal3 s 49200 41216 50000 41336 6 dout1[31]
port 91 nsew signal input
rlabel metal3 s 49200 22992 50000 23112 6 dout1[3]
port 92 nsew signal input
rlabel metal3 s 49200 23672 50000 23792 6 dout1[4]
port 93 nsew signal input
rlabel metal3 s 49200 24216 50000 24336 6 dout1[5]
port 94 nsew signal input
rlabel metal3 s 49200 24896 50000 25016 6 dout1[6]
port 95 nsew signal input
rlabel metal3 s 49200 25576 50000 25696 6 dout1[7]
port 96 nsew signal input
rlabel metal3 s 49200 26256 50000 26376 6 dout1[8]
port 97 nsew signal input
rlabel metal3 s 49200 26800 50000 26920 6 dout1[9]
port 98 nsew signal input
rlabel metal2 s 202 49200 258 50000 6 io_in[0]
port 99 nsew signal input
rlabel metal2 s 12622 49200 12678 50000 6 io_in[10]
port 100 nsew signal input
rlabel metal2 s 13910 49200 13966 50000 6 io_in[11]
port 101 nsew signal input
rlabel metal2 s 15106 49200 15162 50000 6 io_in[12]
port 102 nsew signal input
rlabel metal2 s 16394 49200 16450 50000 6 io_in[13]
port 103 nsew signal input
rlabel metal2 s 17682 49200 17738 50000 6 io_in[14]
port 104 nsew signal input
rlabel metal2 s 18878 49200 18934 50000 6 io_in[15]
port 105 nsew signal input
rlabel metal2 s 20166 49200 20222 50000 6 io_in[16]
port 106 nsew signal input
rlabel metal2 s 21362 49200 21418 50000 6 io_in[17]
port 107 nsew signal input
rlabel metal2 s 22650 49200 22706 50000 6 io_in[18]
port 108 nsew signal input
rlabel metal2 s 23846 49200 23902 50000 6 io_in[19]
port 109 nsew signal input
rlabel metal2 s 1398 49200 1454 50000 6 io_in[1]
port 110 nsew signal input
rlabel metal2 s 25134 49200 25190 50000 6 io_in[20]
port 111 nsew signal input
rlabel metal2 s 26422 49200 26478 50000 6 io_in[21]
port 112 nsew signal input
rlabel metal2 s 27618 49200 27674 50000 6 io_in[22]
port 113 nsew signal input
rlabel metal2 s 28906 49200 28962 50000 6 io_in[23]
port 114 nsew signal input
rlabel metal2 s 30102 49200 30158 50000 6 io_in[24]
port 115 nsew signal input
rlabel metal2 s 31390 49200 31446 50000 6 io_in[25]
port 116 nsew signal input
rlabel metal2 s 32586 49200 32642 50000 6 io_in[26]
port 117 nsew signal input
rlabel metal2 s 33874 49200 33930 50000 6 io_in[27]
port 118 nsew signal input
rlabel metal2 s 35162 49200 35218 50000 6 io_in[28]
port 119 nsew signal input
rlabel metal2 s 36358 49200 36414 50000 6 io_in[29]
port 120 nsew signal input
rlabel metal2 s 2686 49200 2742 50000 6 io_in[2]
port 121 nsew signal input
rlabel metal2 s 37646 49200 37702 50000 6 io_in[30]
port 122 nsew signal input
rlabel metal2 s 38842 49200 38898 50000 6 io_in[31]
port 123 nsew signal input
rlabel metal2 s 40130 49200 40186 50000 6 io_in[32]
port 124 nsew signal input
rlabel metal2 s 41326 49200 41382 50000 6 io_in[33]
port 125 nsew signal input
rlabel metal2 s 42614 49200 42670 50000 6 io_in[34]
port 126 nsew signal input
rlabel metal2 s 43902 49200 43958 50000 6 io_in[35]
port 127 nsew signal input
rlabel metal2 s 45098 49200 45154 50000 6 io_in[36]
port 128 nsew signal input
rlabel metal2 s 46386 49200 46442 50000 6 io_in[37]
port 129 nsew signal input
rlabel metal2 s 3882 49200 3938 50000 6 io_in[3]
port 130 nsew signal input
rlabel metal2 s 5170 49200 5226 50000 6 io_in[4]
port 131 nsew signal input
rlabel metal2 s 6366 49200 6422 50000 6 io_in[5]
port 132 nsew signal input
rlabel metal2 s 7654 49200 7710 50000 6 io_in[6]
port 133 nsew signal input
rlabel metal2 s 8942 49200 8998 50000 6 io_in[7]
port 134 nsew signal input
rlabel metal2 s 10138 49200 10194 50000 6 io_in[8]
port 135 nsew signal input
rlabel metal2 s 11426 49200 11482 50000 6 io_in[9]
port 136 nsew signal input
rlabel metal2 s 570 49200 626 50000 6 io_oeb[0]
port 137 nsew signal output
rlabel metal2 s 13082 49200 13138 50000 6 io_oeb[10]
port 138 nsew signal output
rlabel metal2 s 14278 49200 14334 50000 6 io_oeb[11]
port 139 nsew signal output
rlabel metal2 s 15566 49200 15622 50000 6 io_oeb[12]
port 140 nsew signal output
rlabel metal2 s 16854 49200 16910 50000 6 io_oeb[13]
port 141 nsew signal output
rlabel metal2 s 18050 49200 18106 50000 6 io_oeb[14]
port 142 nsew signal output
rlabel metal2 s 19338 49200 19394 50000 6 io_oeb[15]
port 143 nsew signal output
rlabel metal2 s 20534 49200 20590 50000 6 io_oeb[16]
port 144 nsew signal output
rlabel metal2 s 21822 49200 21878 50000 6 io_oeb[17]
port 145 nsew signal output
rlabel metal2 s 23018 49200 23074 50000 6 io_oeb[18]
port 146 nsew signal output
rlabel metal2 s 24306 49200 24362 50000 6 io_oeb[19]
port 147 nsew signal output
rlabel metal2 s 1858 49200 1914 50000 6 io_oeb[1]
port 148 nsew signal output
rlabel metal2 s 25594 49200 25650 50000 6 io_oeb[20]
port 149 nsew signal output
rlabel metal2 s 26790 49200 26846 50000 6 io_oeb[21]
port 150 nsew signal output
rlabel metal2 s 28078 49200 28134 50000 6 io_oeb[22]
port 151 nsew signal output
rlabel metal2 s 29274 49200 29330 50000 6 io_oeb[23]
port 152 nsew signal output
rlabel metal2 s 30562 49200 30618 50000 6 io_oeb[24]
port 153 nsew signal output
rlabel metal2 s 31758 49200 31814 50000 6 io_oeb[25]
port 154 nsew signal output
rlabel metal2 s 33046 49200 33102 50000 6 io_oeb[26]
port 155 nsew signal output
rlabel metal2 s 34334 49200 34390 50000 6 io_oeb[27]
port 156 nsew signal output
rlabel metal2 s 35530 49200 35586 50000 6 io_oeb[28]
port 157 nsew signal output
rlabel metal2 s 36818 49200 36874 50000 6 io_oeb[29]
port 158 nsew signal output
rlabel metal2 s 3054 49200 3110 50000 6 io_oeb[2]
port 159 nsew signal output
rlabel metal2 s 38014 49200 38070 50000 6 io_oeb[30]
port 160 nsew signal output
rlabel metal2 s 39302 49200 39358 50000 6 io_oeb[31]
port 161 nsew signal output
rlabel metal2 s 40498 49200 40554 50000 6 io_oeb[32]
port 162 nsew signal output
rlabel metal2 s 41786 49200 41842 50000 6 io_oeb[33]
port 163 nsew signal output
rlabel metal2 s 43074 49200 43130 50000 6 io_oeb[34]
port 164 nsew signal output
rlabel metal2 s 44270 49200 44326 50000 6 io_oeb[35]
port 165 nsew signal output
rlabel metal2 s 45558 49200 45614 50000 6 io_oeb[36]
port 166 nsew signal output
rlabel metal2 s 46754 49200 46810 50000 6 io_oeb[37]
port 167 nsew signal output
rlabel metal2 s 4342 49200 4398 50000 6 io_oeb[3]
port 168 nsew signal output
rlabel metal2 s 5538 49200 5594 50000 6 io_oeb[4]
port 169 nsew signal output
rlabel metal2 s 6826 49200 6882 50000 6 io_oeb[5]
port 170 nsew signal output
rlabel metal2 s 8022 49200 8078 50000 6 io_oeb[6]
port 171 nsew signal output
rlabel metal2 s 9310 49200 9366 50000 6 io_oeb[7]
port 172 nsew signal output
rlabel metal2 s 10598 49200 10654 50000 6 io_oeb[8]
port 173 nsew signal output
rlabel metal2 s 11794 49200 11850 50000 6 io_oeb[9]
port 174 nsew signal output
rlabel metal2 s 1030 49200 1086 50000 6 io_out[0]
port 175 nsew signal output
rlabel metal2 s 13450 49200 13506 50000 6 io_out[10]
port 176 nsew signal output
rlabel metal2 s 14738 49200 14794 50000 6 io_out[11]
port 177 nsew signal output
rlabel metal2 s 15934 49200 15990 50000 6 io_out[12]
port 178 nsew signal output
rlabel metal2 s 17222 49200 17278 50000 6 io_out[13]
port 179 nsew signal output
rlabel metal2 s 18510 49200 18566 50000 6 io_out[14]
port 180 nsew signal output
rlabel metal2 s 19706 49200 19762 50000 6 io_out[15]
port 181 nsew signal output
rlabel metal2 s 20994 49200 21050 50000 6 io_out[16]
port 182 nsew signal output
rlabel metal2 s 22190 49200 22246 50000 6 io_out[17]
port 183 nsew signal output
rlabel metal2 s 23478 49200 23534 50000 6 io_out[18]
port 184 nsew signal output
rlabel metal2 s 24674 49200 24730 50000 6 io_out[19]
port 185 nsew signal output
rlabel metal2 s 2226 49200 2282 50000 6 io_out[1]
port 186 nsew signal output
rlabel metal2 s 25962 49200 26018 50000 6 io_out[20]
port 187 nsew signal output
rlabel metal2 s 27250 49200 27306 50000 6 io_out[21]
port 188 nsew signal output
rlabel metal2 s 28446 49200 28502 50000 6 io_out[22]
port 189 nsew signal output
rlabel metal2 s 29734 49200 29790 50000 6 io_out[23]
port 190 nsew signal output
rlabel metal2 s 30930 49200 30986 50000 6 io_out[24]
port 191 nsew signal output
rlabel metal2 s 32218 49200 32274 50000 6 io_out[25]
port 192 nsew signal output
rlabel metal2 s 33506 49200 33562 50000 6 io_out[26]
port 193 nsew signal output
rlabel metal2 s 34702 49200 34758 50000 6 io_out[27]
port 194 nsew signal output
rlabel metal2 s 35990 49200 36046 50000 6 io_out[28]
port 195 nsew signal output
rlabel metal2 s 37186 49200 37242 50000 6 io_out[29]
port 196 nsew signal output
rlabel metal2 s 3514 49200 3570 50000 6 io_out[2]
port 197 nsew signal output
rlabel metal2 s 38474 49200 38530 50000 6 io_out[30]
port 198 nsew signal output
rlabel metal2 s 39670 49200 39726 50000 6 io_out[31]
port 199 nsew signal output
rlabel metal2 s 40958 49200 41014 50000 6 io_out[32]
port 200 nsew signal output
rlabel metal2 s 42246 49200 42302 50000 6 io_out[33]
port 201 nsew signal output
rlabel metal2 s 43442 49200 43498 50000 6 io_out[34]
port 202 nsew signal output
rlabel metal2 s 44730 49200 44786 50000 6 io_out[35]
port 203 nsew signal output
rlabel metal2 s 45926 49200 45982 50000 6 io_out[36]
port 204 nsew signal output
rlabel metal2 s 47214 49200 47270 50000 6 io_out[37]
port 205 nsew signal output
rlabel metal2 s 4710 49200 4766 50000 6 io_out[3]
port 206 nsew signal output
rlabel metal2 s 5998 49200 6054 50000 6 io_out[4]
port 207 nsew signal output
rlabel metal2 s 7194 49200 7250 50000 6 io_out[5]
port 208 nsew signal output
rlabel metal2 s 8482 49200 8538 50000 6 io_out[6]
port 209 nsew signal output
rlabel metal2 s 9770 49200 9826 50000 6 io_out[7]
port 210 nsew signal output
rlabel metal2 s 10966 49200 11022 50000 6 io_out[8]
port 211 nsew signal output
rlabel metal2 s 12254 49200 12310 50000 6 io_out[9]
port 212 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 irq[0]
port 213 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 irq[1]
port 214 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 irq[2]
port 215 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 la_data_in[0]
port 216 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[100]
port 217 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[101]
port 218 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[102]
port 219 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[103]
port 220 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[104]
port 221 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_data_in[105]
port 222 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[106]
port 223 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_data_in[107]
port 224 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_data_in[108]
port 225 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_data_in[109]
port 226 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 la_data_in[10]
port 227 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[110]
port 228 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_data_in[111]
port 229 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[112]
port 230 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[113]
port 231 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[114]
port 232 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[115]
port 233 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_data_in[116]
port 234 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[117]
port 235 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_data_in[118]
port 236 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_data_in[119]
port 237 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 la_data_in[11]
port 238 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[120]
port 239 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[121]
port 240 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_data_in[122]
port 241 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_data_in[123]
port 242 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[124]
port 243 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[125]
port 244 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[126]
port 245 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[127]
port 246 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 la_data_in[12]
port 247 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 la_data_in[13]
port 248 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 la_data_in[14]
port 249 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 la_data_in[15]
port 250 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 la_data_in[16]
port 251 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 la_data_in[17]
port 252 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 la_data_in[18]
port 253 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 la_data_in[19]
port 254 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 la_data_in[1]
port 255 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 la_data_in[20]
port 256 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 la_data_in[21]
port 257 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 la_data_in[22]
port 258 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 la_data_in[23]
port 259 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 la_data_in[24]
port 260 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 la_data_in[25]
port 261 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 la_data_in[26]
port 262 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 la_data_in[27]
port 263 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 la_data_in[28]
port 264 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 la_data_in[29]
port 265 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 la_data_in[2]
port 266 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 la_data_in[30]
port 267 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 la_data_in[31]
port 268 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 la_data_in[32]
port 269 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 la_data_in[33]
port 270 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 la_data_in[34]
port 271 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 la_data_in[35]
port 272 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 la_data_in[36]
port 273 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_data_in[37]
port 274 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 la_data_in[38]
port 275 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 la_data_in[39]
port 276 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 la_data_in[3]
port 277 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_data_in[40]
port 278 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 la_data_in[41]
port 279 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 la_data_in[42]
port 280 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[43]
port 281 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 la_data_in[44]
port 282 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_data_in[45]
port 283 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 la_data_in[46]
port 284 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 la_data_in[47]
port 285 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 la_data_in[48]
port 286 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[49]
port 287 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 la_data_in[4]
port 288 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 la_data_in[50]
port 289 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_data_in[51]
port 290 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 la_data_in[52]
port 291 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_data_in[53]
port 292 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_data_in[54]
port 293 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[55]
port 294 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_data_in[56]
port 295 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[57]
port 296 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 la_data_in[58]
port 297 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 la_data_in[59]
port 298 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 la_data_in[5]
port 299 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 la_data_in[60]
port 300 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 la_data_in[61]
port 301 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 la_data_in[62]
port 302 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 la_data_in[63]
port 303 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_data_in[64]
port 304 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_data_in[65]
port 305 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 la_data_in[66]
port 306 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_data_in[67]
port 307 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_data_in[68]
port 308 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_data_in[69]
port 309 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 la_data_in[6]
port 310 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_data_in[70]
port 311 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_data_in[71]
port 312 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_data_in[72]
port 313 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_data_in[73]
port 314 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 la_data_in[74]
port 315 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 la_data_in[75]
port 316 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_data_in[76]
port 317 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in[77]
port 318 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_data_in[78]
port 319 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_data_in[79]
port 320 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 la_data_in[7]
port 321 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[80]
port 322 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_data_in[81]
port 323 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 la_data_in[82]
port 324 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[83]
port 325 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 la_data_in[84]
port 326 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_data_in[85]
port 327 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_data_in[86]
port 328 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_data_in[87]
port 329 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_data_in[88]
port 330 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_data_in[89]
port 331 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 la_data_in[8]
port 332 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_data_in[90]
port 333 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_data_in[91]
port 334 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[92]
port 335 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_data_in[93]
port 336 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_data_in[94]
port 337 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_data_in[95]
port 338 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_in[96]
port 339 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[97]
port 340 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[98]
port 341 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[99]
port 342 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 la_data_in[9]
port 343 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 la_data_out[0]
port 344 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 la_data_out[100]
port 345 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[101]
port 346 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 la_data_out[102]
port 347 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 la_data_out[103]
port 348 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[104]
port 349 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 la_data_out[105]
port 350 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 la_data_out[106]
port 351 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 la_data_out[107]
port 352 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 la_data_out[108]
port 353 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 la_data_out[109]
port 354 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 la_data_out[10]
port 355 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 la_data_out[110]
port 356 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 la_data_out[111]
port 357 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 la_data_out[112]
port 358 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 la_data_out[113]
port 359 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[114]
port 360 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 la_data_out[115]
port 361 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[116]
port 362 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 la_data_out[117]
port 363 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 la_data_out[118]
port 364 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 la_data_out[119]
port 365 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 la_data_out[11]
port 366 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 la_data_out[120]
port 367 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 la_data_out[121]
port 368 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_data_out[122]
port 369 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 la_data_out[123]
port 370 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 la_data_out[124]
port 371 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[125]
port 372 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[126]
port 373 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[127]
port 374 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 la_data_out[12]
port 375 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 la_data_out[13]
port 376 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 la_data_out[14]
port 377 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 la_data_out[15]
port 378 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 la_data_out[16]
port 379 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 la_data_out[17]
port 380 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 la_data_out[18]
port 381 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 la_data_out[19]
port 382 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 la_data_out[1]
port 383 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 la_data_out[20]
port 384 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 la_data_out[21]
port 385 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 la_data_out[22]
port 386 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 la_data_out[23]
port 387 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 la_data_out[24]
port 388 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 la_data_out[25]
port 389 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 la_data_out[26]
port 390 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 la_data_out[27]
port 391 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 la_data_out[28]
port 392 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 la_data_out[29]
port 393 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 la_data_out[2]
port 394 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 la_data_out[30]
port 395 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 la_data_out[31]
port 396 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 la_data_out[32]
port 397 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 la_data_out[33]
port 398 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 la_data_out[34]
port 399 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 la_data_out[35]
port 400 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 la_data_out[36]
port 401 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 la_data_out[37]
port 402 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 la_data_out[38]
port 403 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 la_data_out[39]
port 404 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 la_data_out[3]
port 405 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 la_data_out[40]
port 406 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 la_data_out[41]
port 407 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 la_data_out[42]
port 408 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 la_data_out[43]
port 409 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 la_data_out[44]
port 410 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 la_data_out[45]
port 411 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 la_data_out[46]
port 412 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 la_data_out[47]
port 413 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 la_data_out[48]
port 414 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 la_data_out[49]
port 415 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 la_data_out[4]
port 416 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 la_data_out[50]
port 417 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 la_data_out[51]
port 418 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 la_data_out[52]
port 419 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 la_data_out[53]
port 420 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 la_data_out[54]
port 421 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 la_data_out[55]
port 422 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 la_data_out[56]
port 423 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 la_data_out[57]
port 424 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 la_data_out[58]
port 425 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 la_data_out[59]
port 426 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 la_data_out[5]
port 427 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 la_data_out[60]
port 428 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 la_data_out[61]
port 429 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 la_data_out[62]
port 430 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 la_data_out[63]
port 431 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 la_data_out[64]
port 432 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 la_data_out[65]
port 433 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 la_data_out[66]
port 434 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 la_data_out[67]
port 435 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 la_data_out[68]
port 436 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 la_data_out[69]
port 437 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 la_data_out[6]
port 438 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 la_data_out[70]
port 439 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 la_data_out[71]
port 440 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 la_data_out[72]
port 441 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 la_data_out[73]
port 442 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 la_data_out[74]
port 443 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 la_data_out[75]
port 444 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 la_data_out[76]
port 445 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 la_data_out[77]
port 446 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 la_data_out[78]
port 447 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 la_data_out[79]
port 448 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 la_data_out[7]
port 449 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 la_data_out[80]
port 450 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 la_data_out[81]
port 451 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 la_data_out[82]
port 452 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 la_data_out[83]
port 453 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[84]
port 454 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 la_data_out[85]
port 455 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 la_data_out[86]
port 456 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 la_data_out[87]
port 457 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 la_data_out[88]
port 458 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 la_data_out[89]
port 459 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 la_data_out[8]
port 460 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[90]
port 461 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 la_data_out[91]
port 462 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[92]
port 463 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 la_data_out[93]
port 464 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 la_data_out[94]
port 465 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 la_data_out[95]
port 466 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 la_data_out[96]
port 467 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 la_data_out[97]
port 468 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 la_data_out[98]
port 469 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 la_data_out[99]
port 470 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 la_data_out[9]
port 471 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 la_oenb[0]
port 472 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_oenb[100]
port 473 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_oenb[101]
port 474 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_oenb[102]
port 475 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_oenb[103]
port 476 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_oenb[104]
port 477 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_oenb[105]
port 478 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_oenb[106]
port 479 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_oenb[107]
port 480 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[108]
port 481 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_oenb[109]
port 482 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 la_oenb[10]
port 483 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_oenb[110]
port 484 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_oenb[111]
port 485 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_oenb[112]
port 486 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_oenb[113]
port 487 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_oenb[114]
port 488 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[115]
port 489 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_oenb[116]
port 490 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[117]
port 491 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_oenb[118]
port 492 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[119]
port 493 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 la_oenb[11]
port 494 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_oenb[120]
port 495 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[121]
port 496 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_oenb[122]
port 497 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_oenb[123]
port 498 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_oenb[124]
port 499 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[125]
port 500 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[126]
port 501 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[127]
port 502 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 la_oenb[12]
port 503 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 la_oenb[13]
port 504 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 la_oenb[14]
port 505 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 la_oenb[15]
port 506 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 la_oenb[16]
port 507 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 la_oenb[17]
port 508 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_oenb[18]
port 509 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 la_oenb[19]
port 510 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 la_oenb[1]
port 511 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 la_oenb[20]
port 512 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 la_oenb[21]
port 513 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 la_oenb[22]
port 514 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 la_oenb[23]
port 515 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 la_oenb[24]
port 516 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 la_oenb[25]
port 517 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 la_oenb[26]
port 518 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 la_oenb[27]
port 519 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 la_oenb[28]
port 520 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 la_oenb[29]
port 521 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 la_oenb[2]
port 522 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 la_oenb[30]
port 523 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 la_oenb[31]
port 524 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 la_oenb[32]
port 525 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 la_oenb[33]
port 526 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 la_oenb[34]
port 527 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_oenb[35]
port 528 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 la_oenb[36]
port 529 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_oenb[37]
port 530 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_oenb[38]
port 531 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 la_oenb[39]
port 532 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 la_oenb[3]
port 533 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 la_oenb[40]
port 534 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 la_oenb[41]
port 535 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 la_oenb[42]
port 536 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 la_oenb[43]
port 537 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_oenb[44]
port 538 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 la_oenb[45]
port 539 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_oenb[46]
port 540 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 la_oenb[47]
port 541 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_oenb[48]
port 542 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 la_oenb[49]
port 543 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 la_oenb[4]
port 544 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_oenb[50]
port 545 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 la_oenb[51]
port 546 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_oenb[52]
port 547 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 la_oenb[53]
port 548 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_oenb[54]
port 549 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 la_oenb[55]
port 550 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_oenb[56]
port 551 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 la_oenb[57]
port 552 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_oenb[58]
port 553 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_oenb[59]
port 554 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_oenb[5]
port 555 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_oenb[60]
port 556 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 la_oenb[61]
port 557 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_oenb[62]
port 558 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la_oenb[63]
port 559 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[64]
port 560 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_oenb[65]
port 561 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_oenb[66]
port 562 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 la_oenb[67]
port 563 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_oenb[68]
port 564 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 la_oenb[69]
port 565 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 la_oenb[6]
port 566 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_oenb[70]
port 567 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 la_oenb[71]
port 568 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_oenb[72]
port 569 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_oenb[73]
port 570 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_oenb[74]
port 571 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_oenb[75]
port 572 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_oenb[76]
port 573 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 la_oenb[77]
port 574 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_oenb[78]
port 575 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_oenb[79]
port 576 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 la_oenb[7]
port 577 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_oenb[80]
port 578 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_oenb[81]
port 579 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_oenb[82]
port 580 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_oenb[83]
port 581 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_oenb[84]
port 582 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_oenb[85]
port 583 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[86]
port 584 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_oenb[87]
port 585 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_oenb[88]
port 586 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_oenb[89]
port 587 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 la_oenb[8]
port 588 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_oenb[90]
port 589 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_oenb[91]
port 590 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_oenb[92]
port 591 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_oenb[93]
port 592 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_oenb[94]
port 593 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_oenb[95]
port 594 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_oenb[96]
port 595 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_oenb[97]
port 596 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 la_oenb[98]
port 597 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[99]
port 598 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 la_oenb[9]
port 599 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 600 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 600 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 601 nsew ground input
rlabel metal2 s 18 0 74 800 6 wb_clk_i
port 602 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_rst_i
port 603 nsew signal input
rlabel metal2 s 202 0 258 800 6 wbs_ack_o
port 604 nsew signal output
rlabel metal2 s 570 0 626 800 6 wbs_adr_i[0]
port 605 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_adr_i[10]
port 606 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[11]
port 607 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[12]
port 608 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_adr_i[13]
port 609 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[14]
port 610 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[15]
port 611 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[16]
port 612 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_adr_i[17]
port 613 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[18]
port 614 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[19]
port 615 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_adr_i[1]
port 616 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_adr_i[20]
port 617 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wbs_adr_i[21]
port 618 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[22]
port 619 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_adr_i[23]
port 620 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[24]
port 621 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[25]
port 622 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[26]
port 623 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[27]
port 624 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[28]
port 625 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_adr_i[29]
port 626 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_adr_i[2]
port 627 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[30]
port 628 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[31]
port 629 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_adr_i[3]
port 630 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[4]
port 631 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_adr_i[5]
port 632 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_adr_i[6]
port 633 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_adr_i[7]
port 634 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_adr_i[8]
port 635 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[9]
port 636 nsew signal input
rlabel metal2 s 294 0 350 800 6 wbs_cyc_i
port 637 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_dat_i[0]
port 638 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[10]
port 639 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_i[11]
port 640 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[12]
port 641 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_i[13]
port 642 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_i[14]
port 643 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[15]
port 644 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[16]
port 645 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_i[17]
port 646 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_i[18]
port 647 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[19]
port 648 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_dat_i[1]
port 649 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[20]
port 650 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_i[21]
port 651 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_i[22]
port 652 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_i[23]
port 653 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[24]
port 654 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_i[25]
port 655 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_i[26]
port 656 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_i[27]
port 657 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[28]
port 658 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_i[29]
port 659 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[2]
port 660 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_i[30]
port 661 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_i[31]
port 662 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_dat_i[3]
port 663 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_dat_i[4]
port 664 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[5]
port 665 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_dat_i[6]
port 666 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_i[7]
port 667 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_dat_i[8]
port 668 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_dat_i[9]
port 669 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_dat_o[0]
port 670 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_o[10]
port 671 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[11]
port 672 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 wbs_dat_o[12]
port 673 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[13]
port 674 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_o[14]
port 675 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 wbs_dat_o[15]
port 676 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_o[16]
port 677 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_o[17]
port 678 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[18]
port 679 nsew signal output
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_o[19]
port 680 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 wbs_dat_o[1]
port 681 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[20]
port 682 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_o[21]
port 683 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_o[22]
port 684 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[23]
port 685 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_o[24]
port 686 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[25]
port 687 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_o[26]
port 688 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[27]
port 689 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[28]
port 690 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[29]
port 691 nsew signal output
rlabel metal2 s 1582 0 1638 800 6 wbs_dat_o[2]
port 692 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[30]
port 693 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_o[31]
port 694 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_o[3]
port 695 nsew signal output
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_o[4]
port 696 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_o[5]
port 697 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[6]
port 698 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_o[7]
port 699 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_o[8]
port 700 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[9]
port 701 nsew signal output
rlabel metal2 s 846 0 902 800 6 wbs_sel_i[0]
port 702 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_sel_i[1]
port 703 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_sel_i[2]
port 704 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_sel_i[3]
port 705 nsew signal input
rlabel metal2 s 386 0 442 800 6 wbs_stb_i
port 706 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_we_i
port 707 nsew signal input
rlabel metal3 s 49200 42440 50000 42560 6 web0
port 708 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 50000 50000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 2443324
string GDS_START 209526
<< end >>

