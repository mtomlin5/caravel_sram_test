magic
tech sky130A
magscale 1 2
timestamp 1636669832
<< locali >>
rect 262597 391527 262631 391765
rect 249073 389283 249107 389929
rect 256617 389351 256651 390405
rect 281089 390031 281123 390133
rect 284953 390133 285229 390167
rect 284953 390099 284987 390133
rect 237297 386971 237331 387277
rect 238033 386495 238067 387277
rect 239137 386631 239171 387277
rect 239965 386563 239999 387277
rect 241069 386699 241103 387277
rect 242173 386767 242207 387277
rect 244289 386835 244323 387277
rect 244841 386903 244875 387277
rect 269129 387039 269163 387277
rect 274741 387107 274775 387277
rect 283849 386427 283883 387277
rect 234721 335359 234755 337841
rect 235457 337603 235491 337977
rect 235641 337603 235675 337773
rect 234813 335427 234847 335529
rect 235917 335427 235951 337841
rect 236193 337263 236227 337909
rect 234663 334577 234755 334611
rect 234721 334135 234755 334577
rect 234813 334577 235641 334611
rect 234629 334067 234663 334101
rect 234813 334067 234847 334577
rect 234629 334033 234847 334067
rect 236469 329851 236503 337773
rect 236653 331347 236687 337773
rect 236929 331959 236963 337841
rect 237481 337535 237515 337773
rect 237757 337603 237791 337909
rect 237849 337263 237883 337909
rect 238033 337603 238067 337841
rect 238493 337603 238527 337841
rect 238585 336379 238619 337909
rect 237297 336039 237331 336277
rect 237205 335631 237239 336005
rect 238677 331959 238711 338045
rect 238769 336515 238803 337909
rect 238861 336175 238895 337909
rect 239229 337603 239263 337909
rect 239413 337331 239447 337569
rect 238953 336447 238987 336685
rect 239505 336379 239539 337909
rect 238953 335937 239171 335971
rect 238953 335835 238987 335937
rect 239045 335631 239079 335869
rect 239137 335767 239171 335937
rect 239229 335699 239263 336141
rect 239413 335835 239447 336209
rect 239321 335631 239355 335665
rect 239045 335597 239355 335631
rect 239873 335359 239907 337841
rect 240333 334611 240367 334713
rect 240425 334611 240459 337841
rect 240701 337535 240735 337841
rect 239045 334135 239079 334577
rect 239505 329307 239539 331789
rect 241069 331347 241103 337909
rect 241253 336515 241287 337909
rect 241713 336991 241747 337841
rect 241345 336379 241379 336481
rect 241621 335495 241655 336753
rect 241805 329647 241839 337841
rect 242173 336583 242207 337977
rect 242265 336583 242299 336821
rect 242357 335563 242391 335801
rect 242541 328967 242575 337773
rect 242817 331959 242851 337909
rect 242909 334951 242943 337977
rect 243001 334135 243035 337841
rect 243277 330667 243311 337841
rect 243369 337535 243403 337841
rect 244013 337535 244047 337841
rect 243737 335767 243771 336889
rect 243921 336039 243955 336549
rect 243829 335767 243863 336005
rect 244381 335903 244415 337841
rect 244565 335631 244599 335937
rect 244507 335597 244599 335631
rect 244749 333591 244783 335801
rect 244841 335427 244875 335869
rect 244933 328695 244967 337773
rect 245117 336379 245151 337841
rect 245209 334135 245243 337909
rect 245301 332095 245335 337773
rect 245485 334951 245519 337909
rect 245577 335495 245611 335665
rect 245393 333387 245427 333489
rect 245669 332639 245703 333285
rect 245761 332163 245795 337773
rect 246129 337535 246163 337841
rect 246865 337535 246899 337841
rect 247049 337535 247083 337841
rect 247325 333999 247359 337841
rect 248337 331891 248371 337909
rect 248429 330463 248463 337841
rect 248521 333659 248555 337909
rect 248797 333727 248831 337841
rect 248521 332707 248555 333217
rect 248981 331143 249015 337841
rect 249073 337535 249107 337841
rect 249625 333931 249659 337841
rect 249993 330327 250027 337773
rect 250085 334883 250119 337841
rect 250545 335087 250579 337909
rect 250821 337331 250855 337773
rect 251005 337331 251039 337909
rect 251373 332911 251407 337909
rect 251465 335223 251499 337773
rect 251557 330259 251591 337909
rect 251649 332843 251683 337909
rect 252017 336107 252051 337841
rect 252477 334407 252511 337909
rect 252661 329987 252695 337909
rect 253121 337535 253155 337841
rect 253305 337535 253339 337773
rect 253397 329919 253431 337909
rect 253581 332027 253615 337773
rect 253765 337535 253799 337909
rect 254041 331279 254075 337501
rect 254225 337331 254259 337841
rect 254317 334611 254351 337773
rect 254501 337331 254535 337977
rect 254961 337195 254995 337977
rect 272659 337977 272751 338011
rect 255145 337331 255179 337773
rect 255237 333251 255271 337909
rect 255789 337331 255823 337909
rect 256341 337535 256375 337841
rect 256525 331279 256559 337909
rect 256893 333251 256927 337841
rect 257169 337535 257203 337909
rect 257353 336039 257387 337909
rect 257445 333183 257479 337909
rect 257629 334679 257663 337909
rect 257905 335631 257939 337773
rect 257997 336243 258031 337909
rect 258089 333319 258123 337841
rect 258365 334883 258399 337773
rect 258549 333931 258583 337841
rect 258641 331551 258675 337909
rect 258917 335223 258951 337909
rect 259101 337535 259135 337909
rect 259469 333115 259503 337909
rect 259653 336515 259687 337909
rect 259837 336719 259871 337841
rect 260205 337535 260239 337909
rect 260481 332911 260515 337909
rect 260573 333183 260607 337841
rect 261125 333047 261159 337841
rect 261401 328831 261435 336617
rect 261769 335087 261803 337909
rect 262045 335971 262079 337841
rect 262137 333183 262171 337841
rect 262413 337535 262447 337909
rect 262689 332979 262723 337841
rect 262873 335563 262907 337841
rect 262965 337535 262999 337841
rect 263241 336787 263275 337909
rect 263057 336039 263091 336481
rect 263241 335631 263275 336549
rect 263425 335835 263459 335937
rect 263425 335801 263551 335835
rect 263517 335767 263551 335801
rect 263701 332571 263735 337841
rect 264253 330327 264287 337909
rect 264529 333183 264563 337841
rect 264621 330531 264655 337909
rect 265081 331755 265115 337909
rect 265265 337331 265299 337909
rect 265449 337535 265483 337909
rect 265725 337263 265759 337773
rect 266369 333863 266403 337841
rect 266553 331007 266587 337909
rect 266645 333659 266679 337909
rect 266829 330939 266863 337909
rect 266921 333523 266955 337841
rect 267381 330803 267415 337909
rect 267749 333455 267783 337841
rect 268025 337535 268059 337841
rect 268025 336651 268059 337025
rect 268025 335767 268059 336073
rect 268117 333319 268151 337841
rect 268209 335971 268243 336957
rect 268393 336175 268427 337909
rect 268979 337841 269071 337875
rect 268519 337773 268611 337807
rect 268335 335597 268519 335631
rect 268485 335495 268519 335597
rect 268301 335291 268335 335461
rect 268209 331143 268243 334509
rect 268577 333251 268611 337773
rect 268853 337535 268887 337841
rect 268761 336311 268795 337161
rect 268853 335563 268887 337229
rect 268393 332707 268427 333081
rect 268761 332979 268795 335393
rect 268945 334951 268979 337297
rect 269037 334339 269071 337841
rect 269221 337195 269255 337909
rect 269163 336685 269255 336719
rect 269221 336583 269255 336685
rect 269497 335767 269531 337977
rect 269773 337535 269807 337841
rect 268669 332911 268703 332945
rect 268853 332911 268887 333081
rect 268669 332877 268887 332911
rect 269589 328967 269623 337501
rect 270049 337263 270083 337909
rect 270325 337535 270359 337841
rect 270417 332571 270451 337909
rect 271061 332367 271095 337841
rect 271337 337535 271371 337841
rect 271521 332639 271555 337841
rect 271797 334815 271831 337841
rect 271889 337535 271923 337841
rect 271981 337127 272015 337909
rect 272073 329783 272107 337909
rect 272199 336141 272441 336175
rect 272625 336107 272659 336413
rect 272717 329647 272751 337977
rect 272993 337535 273027 337909
rect 272809 336651 272843 336957
rect 272993 336651 273027 336889
rect 273085 336719 273119 337025
rect 273177 336651 273211 336753
rect 273085 336617 273211 336651
rect 273085 336515 273119 336617
rect 273027 336481 273119 336515
rect 272809 335427 272843 336345
rect 273085 335495 273119 335937
rect 273177 335903 273211 336549
rect 273269 336107 273303 336821
rect 273821 336787 273855 337841
rect 273729 336311 273763 336753
rect 272809 335393 272993 335427
rect 273729 335019 273763 335529
rect 273821 335495 273855 336005
rect 272901 329103 272935 334101
rect 273913 332027 273947 337841
rect 274189 336243 274223 336481
rect 274281 336243 274315 336957
rect 274373 331347 274407 337841
rect 274465 335835 274499 337909
rect 274925 334271 274959 337909
rect 275477 335359 275511 337909
rect 275661 337535 275695 337841
rect 275753 335495 275787 337297
rect 276213 332231 276247 338181
rect 276397 337841 276581 337875
rect 276305 334815 276339 334985
rect 276397 332095 276431 337841
rect 276581 334271 276615 337501
rect 276765 334883 276799 337909
rect 276857 332435 276891 336957
rect 276949 334135 276983 337501
rect 277593 337127 277627 337909
rect 277041 335087 277075 336821
rect 277317 332435 277351 337093
rect 277409 334475 277443 336821
rect 277869 335359 277903 337841
rect 278145 337331 278179 337909
rect 278237 336107 278271 337841
rect 278329 337535 278363 337909
rect 277961 335971 277995 336073
rect 277961 335937 278363 335971
rect 278329 335903 278363 335937
rect 278329 335869 278697 335903
rect 278789 335835 278823 337773
rect 277961 334067 277995 334849
rect 278053 334339 278087 334781
rect 278329 333999 278363 335461
rect 278513 335427 278547 335733
rect 278881 334067 278915 338249
rect 279249 331959 279283 337977
rect 279709 336855 279743 337841
rect 279525 335903 279559 336073
rect 279801 331959 279835 337841
rect 279893 332571 279927 337025
rect 279985 334407 280019 336889
rect 280169 332673 280387 332707
rect 280169 332639 280203 332673
rect 280353 332639 280387 332673
rect 280123 332605 280203 332639
rect 280123 332571 280157 332605
rect 279893 332537 280157 332571
rect 280261 331891 280295 332605
rect 274281 330531 274315 330633
rect 277317 329715 277351 330633
rect 277259 329681 277351 329715
rect 280445 328695 280479 337841
rect 280721 336855 280755 337841
rect 281181 336991 281215 337909
rect 281365 335495 281399 337909
rect 281733 329239 281767 337909
rect 281825 334611 281859 335869
rect 282009 335495 282043 337909
rect 282193 332163 282227 337909
rect 282285 337535 282319 337909
rect 282561 335291 282595 337501
rect 282929 337059 282963 338113
rect 282745 335291 282779 335801
rect 283481 335563 283515 337501
rect 284401 335903 284435 337841
rect 287529 336923 287563 337093
rect 285229 335767 285263 336889
rect 287713 336787 287747 338045
rect 288081 337127 288115 337773
rect 292773 337195 292807 337297
rect 282929 335189 285229 335223
rect 282929 335155 282963 335189
rect 283113 334543 283147 335053
rect 282285 334067 282319 334373
rect 282285 334033 282469 334067
rect 282745 333999 282779 334441
rect 283791 334373 284527 334407
rect 284033 334135 284067 334237
rect 284493 333999 284527 334373
rect 283113 331483 283147 332061
rect 286609 331415 286643 332061
rect 286701 331891 286735 332061
rect 287805 331279 287839 332197
rect 291761 328695 291795 329545
rect 291853 328763 291887 329477
rect 272717 322507 272751 326417
rect 474749 322643 474783 322881
rect 435925 239683 435959 239989
rect 445619 239853 445861 239887
rect 445711 239785 445953 239819
rect 456165 239547 456199 239649
rect 456015 239513 456199 239547
rect 464721 239581 465031 239615
rect 464721 239547 464755 239581
rect 464813 239411 464847 239513
rect 464997 239479 465031 239581
rect 272441 4879 272475 5457
rect 272533 5219 272567 5457
rect 276121 4675 276155 4845
rect 276213 4199 276247 4641
rect 169585 3077 169769 3111
rect 169585 2975 169619 3077
rect 173081 3043 173115 3893
rect 208409 3043 208443 3893
rect 227729 3655 227763 3825
rect 233893 3791 233927 4097
rect 212825 2975 212859 3621
rect 478245 3383 478279 4029
rect 229569 2975 229603 3349
rect 465733 3247 465767 3349
rect 344201 2941 344845 2975
rect 344201 2907 344235 2941
rect 365637 2771 365671 2941
rect 367109 2771 367143 2941
rect 398205 2941 398389 2975
rect 398205 2839 398239 2941
rect 405565 2839 405599 2941
rect 418721 2771 418755 2941
rect 420285 2839 420319 2941
rect 420227 2805 420319 2839
rect 583401 2839 583435 4777
<< viali >>
rect 262597 391765 262631 391799
rect 262597 391493 262631 391527
rect 256617 390405 256651 390439
rect 249073 389929 249107 389963
rect 281089 390133 281123 390167
rect 285229 390133 285263 390167
rect 284953 390065 284987 390099
rect 281089 389997 281123 390031
rect 256617 389317 256651 389351
rect 249073 389249 249107 389283
rect 237297 387277 237331 387311
rect 237297 386937 237331 386971
rect 238033 387277 238067 387311
rect 239137 387277 239171 387311
rect 239137 386597 239171 386631
rect 239965 387277 239999 387311
rect 241069 387277 241103 387311
rect 242173 387277 242207 387311
rect 244289 387277 244323 387311
rect 244841 387277 244875 387311
rect 269129 387277 269163 387311
rect 274741 387277 274775 387311
rect 274741 387073 274775 387107
rect 283849 387277 283883 387311
rect 269129 387005 269163 387039
rect 244841 386869 244875 386903
rect 244289 386801 244323 386835
rect 242173 386733 242207 386767
rect 241069 386665 241103 386699
rect 239965 386529 239999 386563
rect 238033 386461 238067 386495
rect 283849 386393 283883 386427
rect 278881 338249 278915 338283
rect 276213 338181 276247 338215
rect 238677 338045 238711 338079
rect 235457 337977 235491 338011
rect 234721 337841 234755 337875
rect 236193 337909 236227 337943
rect 235917 337841 235951 337875
rect 235457 337569 235491 337603
rect 235641 337773 235675 337807
rect 235641 337569 235675 337603
rect 234813 335529 234847 335563
rect 234813 335393 234847 335427
rect 237757 337909 237791 337943
rect 236929 337841 236963 337875
rect 236193 337229 236227 337263
rect 236469 337773 236503 337807
rect 235917 335393 235951 335427
rect 234721 335325 234755 335359
rect 234629 334577 234663 334611
rect 234629 334101 234663 334135
rect 234721 334101 234755 334135
rect 235641 334577 235675 334611
rect 236653 337773 236687 337807
rect 237481 337773 237515 337807
rect 237757 337569 237791 337603
rect 237849 337909 237883 337943
rect 237481 337501 237515 337535
rect 238585 337909 238619 337943
rect 238033 337841 238067 337875
rect 238033 337569 238067 337603
rect 238493 337841 238527 337875
rect 238493 337569 238527 337603
rect 237849 337229 237883 337263
rect 238585 336345 238619 336379
rect 237297 336277 237331 336311
rect 237205 336005 237239 336039
rect 237297 336005 237331 336039
rect 237205 335597 237239 335631
rect 236929 331925 236963 331959
rect 242173 337977 242207 338011
rect 238769 337909 238803 337943
rect 238769 336481 238803 336515
rect 238861 337909 238895 337943
rect 239229 337909 239263 337943
rect 239505 337909 239539 337943
rect 239229 337569 239263 337603
rect 239413 337569 239447 337603
rect 239413 337297 239447 337331
rect 238953 336685 238987 336719
rect 238953 336413 238987 336447
rect 241069 337909 241103 337943
rect 239505 336345 239539 336379
rect 239873 337841 239907 337875
rect 239413 336209 239447 336243
rect 238861 336141 238895 336175
rect 239229 336141 239263 336175
rect 238953 335801 238987 335835
rect 239045 335869 239079 335903
rect 239137 335733 239171 335767
rect 239413 335801 239447 335835
rect 239229 335665 239263 335699
rect 239321 335665 239355 335699
rect 239873 335325 239907 335359
rect 240425 337841 240459 337875
rect 240333 334713 240367 334747
rect 239045 334577 239079 334611
rect 240333 334577 240367 334611
rect 240701 337841 240735 337875
rect 240701 337501 240735 337535
rect 240425 334577 240459 334611
rect 239045 334101 239079 334135
rect 238677 331925 238711 331959
rect 236653 331313 236687 331347
rect 239505 331789 239539 331823
rect 236469 329817 236503 329851
rect 241253 337909 241287 337943
rect 241713 337841 241747 337875
rect 241713 336957 241747 336991
rect 241805 337841 241839 337875
rect 241621 336753 241655 336787
rect 241253 336481 241287 336515
rect 241345 336481 241379 336515
rect 241345 336345 241379 336379
rect 241621 335461 241655 335495
rect 241069 331313 241103 331347
rect 242909 337977 242943 338011
rect 242817 337909 242851 337943
rect 242541 337773 242575 337807
rect 242173 336549 242207 336583
rect 242265 336821 242299 336855
rect 242265 336549 242299 336583
rect 242357 335801 242391 335835
rect 242357 335529 242391 335563
rect 241805 329613 241839 329647
rect 239505 329273 239539 329307
rect 254501 337977 254535 338011
rect 245209 337909 245243 337943
rect 242909 334917 242943 334951
rect 243001 337841 243035 337875
rect 243001 334101 243035 334135
rect 243277 337841 243311 337875
rect 242817 331925 242851 331959
rect 243369 337841 243403 337875
rect 243369 337501 243403 337535
rect 244013 337841 244047 337875
rect 244013 337501 244047 337535
rect 244381 337841 244415 337875
rect 243737 336889 243771 336923
rect 243921 336549 243955 336583
rect 243737 335733 243771 335767
rect 243829 336005 243863 336039
rect 243921 336005 243955 336039
rect 245117 337841 245151 337875
rect 244933 337773 244967 337807
rect 244381 335869 244415 335903
rect 244565 335937 244599 335971
rect 243829 335733 243863 335767
rect 244841 335869 244875 335903
rect 244473 335597 244507 335631
rect 244749 335801 244783 335835
rect 244841 335393 244875 335427
rect 244749 333557 244783 333591
rect 243277 330633 243311 330667
rect 242541 328933 242575 328967
rect 245117 336345 245151 336379
rect 245485 337909 245519 337943
rect 245209 334101 245243 334135
rect 245301 337773 245335 337807
rect 248337 337909 248371 337943
rect 246129 337841 246163 337875
rect 245761 337773 245795 337807
rect 245577 335665 245611 335699
rect 245577 335461 245611 335495
rect 245485 334917 245519 334951
rect 245393 333489 245427 333523
rect 245393 333353 245427 333387
rect 245669 333285 245703 333319
rect 245669 332605 245703 332639
rect 246129 337501 246163 337535
rect 246865 337841 246899 337875
rect 246865 337501 246899 337535
rect 247049 337841 247083 337875
rect 247049 337501 247083 337535
rect 247325 337841 247359 337875
rect 247325 333965 247359 333999
rect 245761 332129 245795 332163
rect 245301 332061 245335 332095
rect 248521 337909 248555 337943
rect 248337 331857 248371 331891
rect 248429 337841 248463 337875
rect 250545 337909 250579 337943
rect 248797 337841 248831 337875
rect 248797 333693 248831 333727
rect 248981 337841 249015 337875
rect 248521 333625 248555 333659
rect 248521 333217 248555 333251
rect 248521 332673 248555 332707
rect 249073 337841 249107 337875
rect 249073 337501 249107 337535
rect 249625 337841 249659 337875
rect 250085 337841 250119 337875
rect 249625 333897 249659 333931
rect 249993 337773 250027 337807
rect 248981 331109 249015 331143
rect 248429 330429 248463 330463
rect 251005 337909 251039 337943
rect 250821 337773 250855 337807
rect 250821 337297 250855 337331
rect 251005 337297 251039 337331
rect 251373 337909 251407 337943
rect 250545 335053 250579 335087
rect 250085 334849 250119 334883
rect 251557 337909 251591 337943
rect 251465 337773 251499 337807
rect 251465 335189 251499 335223
rect 251373 332877 251407 332911
rect 249993 330293 250027 330327
rect 251649 337909 251683 337943
rect 252477 337909 252511 337943
rect 252017 337841 252051 337875
rect 252017 336073 252051 336107
rect 252477 334373 252511 334407
rect 252661 337909 252695 337943
rect 251649 332809 251683 332843
rect 251557 330225 251591 330259
rect 253397 337909 253431 337943
rect 253121 337841 253155 337875
rect 253121 337501 253155 337535
rect 253305 337773 253339 337807
rect 253305 337501 253339 337535
rect 252661 329953 252695 329987
rect 253765 337909 253799 337943
rect 253581 337773 253615 337807
rect 254225 337841 254259 337875
rect 253765 337501 253799 337535
rect 254041 337501 254075 337535
rect 253581 331993 253615 332027
rect 254225 337297 254259 337331
rect 254317 337773 254351 337807
rect 254501 337297 254535 337331
rect 254961 337977 254995 338011
rect 269497 337977 269531 338011
rect 272625 337977 272659 338011
rect 255237 337909 255271 337943
rect 255145 337773 255179 337807
rect 255145 337297 255179 337331
rect 254961 337161 254995 337195
rect 254317 334577 254351 334611
rect 255789 337909 255823 337943
rect 256525 337909 256559 337943
rect 256341 337841 256375 337875
rect 256341 337501 256375 337535
rect 255789 337297 255823 337331
rect 255237 333217 255271 333251
rect 254041 331245 254075 331279
rect 257169 337909 257203 337943
rect 256893 337841 256927 337875
rect 257169 337501 257203 337535
rect 257353 337909 257387 337943
rect 257353 336005 257387 336039
rect 257445 337909 257479 337943
rect 256893 333217 256927 333251
rect 257629 337909 257663 337943
rect 257997 337909 258031 337943
rect 257905 337773 257939 337807
rect 258641 337909 258675 337943
rect 257997 336209 258031 336243
rect 258089 337841 258123 337875
rect 257905 335597 257939 335631
rect 257629 334645 257663 334679
rect 258549 337841 258583 337875
rect 258365 337773 258399 337807
rect 258365 334849 258399 334883
rect 258549 333897 258583 333931
rect 258089 333285 258123 333319
rect 257445 333149 257479 333183
rect 258917 337909 258951 337943
rect 259101 337909 259135 337943
rect 259101 337501 259135 337535
rect 259469 337909 259503 337943
rect 258917 335189 258951 335223
rect 259653 337909 259687 337943
rect 260205 337909 260239 337943
rect 259837 337841 259871 337875
rect 260205 337501 260239 337535
rect 260481 337909 260515 337943
rect 259837 336685 259871 336719
rect 259653 336481 259687 336515
rect 259469 333081 259503 333115
rect 261769 337909 261803 337943
rect 260573 337841 260607 337875
rect 260573 333149 260607 333183
rect 261125 337841 261159 337875
rect 261125 333013 261159 333047
rect 261401 336617 261435 336651
rect 260481 332877 260515 332911
rect 258641 331517 258675 331551
rect 256525 331245 256559 331279
rect 253397 329885 253431 329919
rect 262413 337909 262447 337943
rect 262045 337841 262079 337875
rect 262045 335937 262079 335971
rect 262137 337841 262171 337875
rect 261769 335053 261803 335087
rect 263241 337909 263275 337943
rect 262413 337501 262447 337535
rect 262689 337841 262723 337875
rect 262137 333149 262171 333183
rect 262873 337841 262907 337875
rect 262965 337841 262999 337875
rect 262965 337501 262999 337535
rect 264253 337909 264287 337943
rect 263241 336753 263275 336787
rect 263701 337841 263735 337875
rect 263241 336549 263275 336583
rect 263057 336481 263091 336515
rect 263057 336005 263091 336039
rect 263425 335937 263459 335971
rect 263517 335733 263551 335767
rect 263241 335597 263275 335631
rect 262873 335529 262907 335563
rect 262689 332945 262723 332979
rect 263701 332537 263735 332571
rect 264621 337909 264655 337943
rect 264529 337841 264563 337875
rect 264529 333149 264563 333183
rect 265081 337909 265115 337943
rect 265265 337909 265299 337943
rect 265449 337909 265483 337943
rect 266553 337909 266587 337943
rect 266369 337841 266403 337875
rect 265449 337501 265483 337535
rect 265725 337773 265759 337807
rect 265265 337297 265299 337331
rect 265725 337229 265759 337263
rect 266369 333829 266403 333863
rect 265081 331721 265115 331755
rect 266645 337909 266679 337943
rect 266645 333625 266679 333659
rect 266829 337909 266863 337943
rect 266553 330973 266587 331007
rect 267381 337909 267415 337943
rect 266921 337841 266955 337875
rect 266921 333489 266955 333523
rect 266829 330905 266863 330939
rect 268393 337909 268427 337943
rect 267749 337841 267783 337875
rect 268025 337841 268059 337875
rect 268025 337501 268059 337535
rect 268117 337841 268151 337875
rect 268025 337025 268059 337059
rect 268025 336617 268059 336651
rect 268025 336073 268059 336107
rect 268025 335733 268059 335767
rect 267749 333421 267783 333455
rect 268209 336957 268243 336991
rect 269221 337909 269255 337943
rect 268853 337841 268887 337875
rect 268945 337841 268979 337875
rect 268485 337773 268519 337807
rect 268393 336141 268427 336175
rect 268209 335937 268243 335971
rect 268301 335597 268335 335631
rect 268301 335461 268335 335495
rect 268485 335461 268519 335495
rect 268301 335257 268335 335291
rect 268117 333285 268151 333319
rect 268209 334509 268243 334543
rect 268853 337501 268887 337535
rect 268945 337297 268979 337331
rect 268853 337229 268887 337263
rect 268761 337161 268795 337195
rect 268761 336277 268795 336311
rect 268853 335529 268887 335563
rect 268577 333217 268611 333251
rect 268761 335393 268795 335427
rect 268393 333081 268427 333115
rect 268945 334917 268979 334951
rect 269221 337161 269255 337195
rect 269129 336685 269163 336719
rect 269221 336549 269255 336583
rect 270049 337909 270083 337943
rect 269773 337841 269807 337875
rect 269497 335733 269531 335767
rect 269589 337501 269623 337535
rect 269773 337501 269807 337535
rect 269037 334305 269071 334339
rect 268669 332945 268703 332979
rect 268761 332945 268795 332979
rect 268853 333081 268887 333115
rect 268393 332673 268427 332707
rect 268209 331109 268243 331143
rect 267381 330769 267415 330803
rect 264621 330497 264655 330531
rect 264253 330293 264287 330327
rect 270417 337909 270451 337943
rect 270325 337841 270359 337875
rect 270325 337501 270359 337535
rect 270049 337229 270083 337263
rect 271981 337909 272015 337943
rect 270417 332537 270451 332571
rect 271061 337841 271095 337875
rect 271337 337841 271371 337875
rect 271337 337501 271371 337535
rect 271521 337841 271555 337875
rect 271797 337841 271831 337875
rect 271889 337841 271923 337875
rect 271889 337501 271923 337535
rect 271981 337093 272015 337127
rect 272073 337909 272107 337943
rect 271797 334781 271831 334815
rect 271521 332605 271555 332639
rect 271061 332333 271095 332367
rect 272625 336413 272659 336447
rect 272165 336141 272199 336175
rect 272441 336141 272475 336175
rect 272625 336073 272659 336107
rect 272073 329749 272107 329783
rect 272993 337909 273027 337943
rect 274465 337909 274499 337943
rect 272993 337501 273027 337535
rect 273821 337841 273855 337875
rect 273085 337025 273119 337059
rect 272809 336957 272843 336991
rect 272809 336617 272843 336651
rect 272993 336889 273027 336923
rect 273269 336821 273303 336855
rect 273085 336685 273119 336719
rect 273177 336753 273211 336787
rect 272993 336617 273027 336651
rect 272993 336481 273027 336515
rect 273177 336549 273211 336583
rect 272809 336345 272843 336379
rect 273085 335937 273119 335971
rect 273729 336753 273763 336787
rect 273821 336753 273855 336787
rect 273913 337841 273947 337875
rect 273729 336277 273763 336311
rect 273269 336073 273303 336107
rect 273177 335869 273211 335903
rect 273821 336005 273855 336039
rect 273085 335461 273119 335495
rect 273729 335529 273763 335563
rect 272993 335393 273027 335427
rect 273821 335461 273855 335495
rect 273729 334985 273763 335019
rect 272717 329613 272751 329647
rect 272901 334101 272935 334135
rect 274373 337841 274407 337875
rect 274281 336957 274315 336991
rect 274189 336481 274223 336515
rect 274189 336209 274223 336243
rect 274281 336209 274315 336243
rect 273913 331993 273947 332027
rect 274465 335801 274499 335835
rect 274925 337909 274959 337943
rect 275477 337909 275511 337943
rect 275661 337841 275695 337875
rect 275661 337501 275695 337535
rect 275753 337297 275787 337331
rect 275753 335461 275787 335495
rect 275477 335325 275511 335359
rect 274925 334237 274959 334271
rect 276765 337909 276799 337943
rect 276581 337841 276615 337875
rect 276305 334985 276339 335019
rect 276305 334781 276339 334815
rect 276213 332197 276247 332231
rect 276581 337501 276615 337535
rect 277593 337909 277627 337943
rect 276949 337501 276983 337535
rect 276765 334849 276799 334883
rect 276857 336957 276891 336991
rect 276581 334237 276615 334271
rect 278145 337909 278179 337943
rect 277317 337093 277351 337127
rect 277593 337093 277627 337127
rect 277869 337841 277903 337875
rect 277041 336821 277075 336855
rect 277041 335053 277075 335087
rect 276949 334101 276983 334135
rect 276857 332401 276891 332435
rect 277409 336821 277443 336855
rect 278329 337909 278363 337943
rect 278145 337297 278179 337331
rect 278237 337841 278271 337875
rect 278329 337501 278363 337535
rect 278789 337773 278823 337807
rect 277961 336073 277995 336107
rect 278237 336073 278271 336107
rect 278697 335869 278731 335903
rect 278789 335801 278823 335835
rect 278513 335733 278547 335767
rect 277869 335325 277903 335359
rect 278329 335461 278363 335495
rect 277409 334441 277443 334475
rect 277961 334849 277995 334883
rect 278053 334781 278087 334815
rect 278053 334305 278087 334339
rect 277961 334033 277995 334067
rect 278513 335393 278547 335427
rect 282929 338113 282963 338147
rect 278881 334033 278915 334067
rect 279249 337977 279283 338011
rect 278329 333965 278363 333999
rect 277317 332401 277351 332435
rect 276397 332061 276431 332095
rect 281181 337909 281215 337943
rect 279709 337841 279743 337875
rect 279709 336821 279743 336855
rect 279801 337841 279835 337875
rect 279525 336073 279559 336107
rect 279525 335869 279559 335903
rect 279249 331925 279283 331959
rect 280445 337841 280479 337875
rect 279893 337025 279927 337059
rect 279985 336889 280019 336923
rect 279985 334373 280019 334407
rect 280261 332605 280295 332639
rect 280353 332605 280387 332639
rect 279801 331925 279835 331959
rect 280261 331857 280295 331891
rect 274373 331313 274407 331347
rect 274281 330633 274315 330667
rect 274281 330497 274315 330531
rect 277317 330633 277351 330667
rect 277225 329681 277259 329715
rect 272901 329069 272935 329103
rect 269589 328933 269623 328967
rect 261401 328797 261435 328831
rect 244933 328661 244967 328695
rect 280721 337841 280755 337875
rect 281181 336957 281215 336991
rect 281365 337909 281399 337943
rect 280721 336821 280755 336855
rect 281365 335461 281399 335495
rect 281733 337909 281767 337943
rect 282009 337909 282043 337943
rect 281825 335869 281859 335903
rect 282009 335461 282043 335495
rect 282193 337909 282227 337943
rect 281825 334577 281859 334611
rect 282285 337909 282319 337943
rect 282285 337501 282319 337535
rect 282561 337501 282595 337535
rect 287713 338045 287747 338079
rect 284401 337841 284435 337875
rect 282929 337025 282963 337059
rect 283481 337501 283515 337535
rect 282561 335257 282595 335291
rect 282745 335801 282779 335835
rect 287529 337093 287563 337127
rect 284401 335869 284435 335903
rect 285229 336889 285263 336923
rect 287529 336889 287563 336923
rect 288081 337773 288115 337807
rect 292773 337297 292807 337331
rect 292773 337161 292807 337195
rect 288081 337093 288115 337127
rect 287713 336753 287747 336787
rect 285229 335733 285263 335767
rect 283481 335529 283515 335563
rect 282745 335257 282779 335291
rect 285229 335189 285263 335223
rect 282929 335121 282963 335155
rect 283113 335053 283147 335087
rect 283113 334509 283147 334543
rect 282745 334441 282779 334475
rect 282285 334373 282319 334407
rect 282469 334033 282503 334067
rect 283757 334373 283791 334407
rect 284033 334237 284067 334271
rect 284033 334101 284067 334135
rect 282745 333965 282779 333999
rect 284493 333965 284527 333999
rect 282193 332129 282227 332163
rect 287805 332197 287839 332231
rect 283113 332061 283147 332095
rect 283113 331449 283147 331483
rect 286609 332061 286643 332095
rect 286701 332061 286735 332095
rect 286701 331857 286735 331891
rect 286609 331381 286643 331415
rect 287805 331245 287839 331279
rect 281733 329205 281767 329239
rect 291761 329545 291795 329579
rect 280445 328661 280479 328695
rect 291853 329477 291887 329511
rect 291853 328729 291887 328763
rect 291761 328661 291795 328695
rect 272717 326417 272751 326451
rect 474749 322881 474783 322915
rect 474749 322609 474783 322643
rect 272717 322473 272751 322507
rect 435925 239989 435959 240023
rect 445585 239853 445619 239887
rect 445861 239853 445895 239887
rect 445677 239785 445711 239819
rect 445953 239785 445987 239819
rect 435925 239649 435959 239683
rect 456165 239649 456199 239683
rect 455981 239513 456015 239547
rect 464721 239513 464755 239547
rect 464813 239513 464847 239547
rect 464997 239445 465031 239479
rect 464813 239377 464847 239411
rect 272441 5457 272475 5491
rect 272533 5457 272567 5491
rect 272533 5185 272567 5219
rect 272441 4845 272475 4879
rect 276121 4845 276155 4879
rect 583401 4777 583435 4811
rect 276121 4641 276155 4675
rect 276213 4641 276247 4675
rect 276213 4165 276247 4199
rect 233893 4097 233927 4131
rect 173081 3893 173115 3927
rect 169769 3077 169803 3111
rect 173081 3009 173115 3043
rect 208409 3893 208443 3927
rect 227729 3825 227763 3859
rect 233893 3757 233927 3791
rect 478245 4029 478279 4063
rect 208409 3009 208443 3043
rect 212825 3621 212859 3655
rect 227729 3621 227763 3655
rect 169585 2941 169619 2975
rect 212825 2941 212859 2975
rect 229569 3349 229603 3383
rect 465733 3349 465767 3383
rect 478245 3349 478279 3383
rect 465733 3213 465767 3247
rect 229569 2941 229603 2975
rect 344845 2941 344879 2975
rect 365637 2941 365671 2975
rect 344201 2873 344235 2907
rect 365637 2737 365671 2771
rect 367109 2941 367143 2975
rect 398389 2941 398423 2975
rect 405565 2941 405599 2975
rect 398205 2805 398239 2839
rect 405565 2805 405599 2839
rect 418721 2941 418755 2975
rect 367109 2737 367143 2771
rect 420285 2941 420319 2975
rect 420193 2805 420227 2839
rect 583401 2805 583435 2839
rect 418721 2737 418755 2771
<< metal1 >>
rect 254946 700952 254952 701004
rect 255004 700992 255010 701004
rect 397454 700992 397460 701004
rect 255004 700964 397460 700992
rect 255004 700952 255010 700964
rect 397454 700952 397460 700964
rect 397512 700952 397518 701004
rect 255038 700884 255044 700936
rect 255096 700924 255102 700936
rect 413646 700924 413652 700936
rect 255096 700896 413652 700924
rect 255096 700884 255102 700896
rect 413646 700884 413652 700896
rect 413704 700884 413710 700936
rect 89162 700816 89168 700868
rect 89220 700856 89226 700868
rect 259638 700856 259644 700868
rect 89220 700828 259644 700856
rect 89220 700816 89226 700828
rect 259638 700816 259644 700828
rect 259696 700816 259702 700868
rect 273898 700816 273904 700868
rect 273956 700856 273962 700868
rect 300118 700856 300124 700868
rect 273956 700828 300124 700856
rect 273956 700816 273962 700828
rect 300118 700816 300124 700828
rect 300176 700816 300182 700868
rect 72970 700748 72976 700800
rect 73028 700788 73034 700800
rect 259730 700788 259736 700800
rect 73028 700760 259736 700788
rect 73028 700748 73034 700760
rect 259730 700748 259736 700760
rect 259788 700748 259794 700800
rect 271138 700748 271144 700800
rect 271196 700788 271202 700800
rect 364978 700788 364984 700800
rect 271196 700760 364984 700788
rect 271196 700748 271202 700760
rect 364978 700748 364984 700760
rect 365036 700748 365042 700800
rect 253658 700680 253664 700732
rect 253716 700720 253722 700732
rect 462314 700720 462320 700732
rect 253716 700692 462320 700720
rect 253716 700680 253722 700692
rect 462314 700680 462320 700692
rect 462372 700680 462378 700732
rect 40494 700612 40500 700664
rect 40552 700652 40558 700664
rect 260834 700652 260840 700664
rect 40552 700624 260840 700652
rect 40552 700612 40558 700624
rect 260834 700612 260840 700624
rect 260892 700612 260898 700664
rect 269758 700612 269764 700664
rect 269816 700652 269822 700664
rect 429838 700652 429844 700664
rect 269816 700624 429844 700652
rect 269816 700612 269822 700624
rect 429838 700612 429844 700624
rect 429896 700612 429902 700664
rect 255130 700544 255136 700596
rect 255188 700584 255194 700596
rect 478506 700584 478512 700596
rect 255188 700556 478512 700584
rect 255188 700544 255194 700556
rect 478506 700544 478512 700556
rect 478564 700544 478570 700596
rect 24302 700476 24308 700528
rect 24360 700516 24366 700528
rect 261018 700516 261024 700528
rect 24360 700488 261024 700516
rect 24360 700476 24366 700488
rect 261018 700476 261024 700488
rect 261076 700476 261082 700528
rect 282178 700476 282184 700528
rect 282236 700516 282242 700528
rect 494790 700516 494796 700528
rect 282236 700488 494796 700516
rect 282236 700476 282242 700488
rect 494790 700476 494796 700488
rect 494848 700476 494854 700528
rect 170306 700408 170312 700460
rect 170364 700448 170370 700460
rect 240778 700448 240784 700460
rect 170364 700420 240784 700448
rect 170364 700408 170370 700420
rect 240778 700408 240784 700420
rect 240836 700408 240842 700460
rect 252186 700408 252192 700460
rect 252244 700448 252250 700460
rect 527174 700448 527180 700460
rect 252244 700420 527180 700448
rect 252244 700408 252250 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 8110 700340 8116 700392
rect 8168 700380 8174 700392
rect 260926 700380 260932 700392
rect 8168 700352 260932 700380
rect 8168 700340 8174 700352
rect 260926 700340 260932 700352
rect 260984 700340 260990 700392
rect 280798 700340 280804 700392
rect 280856 700380 280862 700392
rect 559650 700380 559656 700392
rect 280856 700352 559656 700380
rect 280856 700340 280862 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 105446 700272 105452 700324
rect 105504 700312 105510 700324
rect 242158 700312 242164 700324
rect 105504 700284 242164 700312
rect 105504 700272 105510 700284
rect 242158 700272 242164 700284
rect 242216 700272 242222 700324
rect 253750 700272 253756 700324
rect 253808 700312 253814 700324
rect 543458 700312 543464 700324
rect 253808 700284 543464 700312
rect 253808 700272 253814 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 137830 700204 137836 700256
rect 137888 700244 137894 700256
rect 258166 700244 258172 700256
rect 137888 700216 258172 700244
rect 137888 700204 137894 700216
rect 258166 700204 258172 700216
rect 258224 700204 258230 700256
rect 154114 700136 154120 700188
rect 154172 700176 154178 700188
rect 259546 700176 259552 700188
rect 154172 700148 259552 700176
rect 154172 700136 154178 700148
rect 259546 700136 259552 700148
rect 259604 700136 259610 700188
rect 256418 700068 256424 700120
rect 256476 700108 256482 700120
rect 348786 700108 348792 700120
rect 256476 700080 348792 700108
rect 256476 700068 256482 700080
rect 348786 700068 348792 700080
rect 348844 700068 348850 700120
rect 256510 700000 256516 700052
rect 256568 700040 256574 700052
rect 332502 700040 332508 700052
rect 256568 700012 332508 700040
rect 256568 700000 256574 700012
rect 332502 700000 332508 700012
rect 332560 700000 332566 700052
rect 202782 699932 202788 699984
rect 202840 699972 202846 699984
rect 258258 699972 258264 699984
rect 202840 699944 258264 699972
rect 202840 699932 202846 699944
rect 258258 699932 258264 699944
rect 258316 699932 258322 699984
rect 218974 699864 218980 699916
rect 219032 699904 219038 699916
rect 258350 699904 258356 699916
rect 219032 699876 258356 699904
rect 219032 699864 219038 699876
rect 258350 699864 258356 699876
rect 258408 699864 258414 699916
rect 257890 699796 257896 699848
rect 257948 699836 257954 699848
rect 283834 699836 283840 699848
rect 257948 699808 283840 699836
rect 257948 699796 257954 699808
rect 283834 699796 283840 699808
rect 283892 699796 283898 699848
rect 257982 699728 257988 699780
rect 258040 699768 258046 699780
rect 267642 699768 267648 699780
rect 258040 699740 267648 699768
rect 258040 699728 258046 699740
rect 267642 699728 267648 699740
rect 267700 699728 267706 699780
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 238018 699700 238024 699712
rect 235224 699672 238024 699700
rect 235224 699660 235230 699672
rect 238018 699660 238024 699672
rect 238076 699660 238082 699712
rect 252370 696940 252376 696992
rect 252428 696980 252434 696992
rect 580166 696980 580172 696992
rect 252428 696952 580172 696980
rect 252428 696940 252434 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 261110 683244 261116 683256
rect 3476 683216 261116 683244
rect 3476 683204 3482 683216
rect 261110 683204 261116 683216
rect 261168 683204 261174 683256
rect 252278 683136 252284 683188
rect 252336 683176 252342 683188
rect 580166 683176 580172 683188
rect 252336 683148 580172 683176
rect 252336 683136 252342 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3418 670760 3424 670812
rect 3476 670800 3482 670812
rect 262214 670800 262220 670812
rect 3476 670772 262220 670800
rect 3476 670760 3482 670772
rect 262214 670760 262220 670772
rect 262272 670760 262278 670812
rect 251082 670692 251088 670744
rect 251140 670732 251146 670744
rect 580166 670732 580172 670744
rect 251140 670704 580172 670732
rect 251140 670692 251146 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 262306 656928 262312 656940
rect 3476 656900 262312 656928
rect 3476 656888 3482 656900
rect 262306 656888 262312 656900
rect 262364 656888 262370 656940
rect 250990 643084 250996 643136
rect 251048 643124 251054 643136
rect 580166 643124 580172 643136
rect 251048 643096 580172 643124
rect 251048 643084 251054 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 262398 632108 262404 632120
rect 3476 632080 262404 632108
rect 3476 632068 3482 632080
rect 262398 632068 262404 632080
rect 262456 632068 262462 632120
rect 250898 630640 250904 630692
rect 250956 630680 250962 630692
rect 580166 630680 580172 630692
rect 250956 630652 580172 630680
rect 250956 630640 250962 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 263594 618304 263600 618316
rect 3200 618276 263600 618304
rect 3200 618264 3206 618276
rect 263594 618264 263600 618276
rect 263652 618264 263658 618316
rect 250806 616836 250812 616888
rect 250864 616876 250870 616888
rect 580166 616876 580172 616888
rect 250864 616848 580172 616876
rect 250864 616836 250870 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 263686 605860 263692 605872
rect 3292 605832 263692 605860
rect 3292 605820 3298 605832
rect 263686 605820 263692 605832
rect 263744 605820 263750 605872
rect 249702 590656 249708 590708
rect 249760 590696 249766 590708
rect 579798 590696 579804 590708
rect 249760 590668 579804 590696
rect 249760 590656 249766 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 263778 579680 263784 579692
rect 3384 579652 263784 579680
rect 3384 579640 3390 579652
rect 263778 579640 263784 579652
rect 263836 579640 263842 579692
rect 249610 576852 249616 576904
rect 249668 576892 249674 576904
rect 580166 576892 580172 576904
rect 249668 576864 580172 576892
rect 249668 576852 249674 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 264974 565876 264980 565888
rect 3476 565848 264980 565876
rect 3476 565836 3482 565848
rect 264974 565836 264980 565848
rect 265032 565836 265038 565888
rect 249518 563048 249524 563100
rect 249576 563088 249582 563100
rect 579798 563088 579804 563100
rect 249576 563060 579804 563088
rect 249576 563048 249582 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 263870 553432 263876 553444
rect 3476 553404 263876 553432
rect 3476 553392 3482 553404
rect 263870 553392 263876 553404
rect 263928 553392 263934 553444
rect 248322 536800 248328 536852
rect 248380 536840 248386 536852
rect 580166 536840 580172 536852
rect 248380 536812 580172 536840
rect 248380 536800 248386 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 265066 527184 265072 527196
rect 3476 527156 265072 527184
rect 3476 527144 3482 527156
rect 265066 527144 265072 527156
rect 265124 527144 265130 527196
rect 248230 524424 248236 524476
rect 248288 524464 248294 524476
rect 580166 524464 580172 524476
rect 248288 524436 580172 524464
rect 248288 524424 248294 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 265158 514808 265164 514820
rect 3476 514780 265164 514808
rect 3476 514768 3482 514780
rect 265158 514768 265164 514780
rect 265216 514768 265222 514820
rect 248138 510620 248144 510672
rect 248196 510660 248202 510672
rect 580166 510660 580172 510672
rect 248196 510632 580172 510660
rect 248196 510620 248202 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 265250 501004 265256 501016
rect 3108 500976 265256 501004
rect 3108 500964 3114 500976
rect 265250 500964 265256 500976
rect 265308 500964 265314 501016
rect 246942 484372 246948 484424
rect 247000 484412 247006 484424
rect 580166 484412 580172 484424
rect 247000 484384 580172 484412
rect 247000 484372 247006 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 266354 474756 266360 474768
rect 3476 474728 266360 474756
rect 3476 474716 3482 474728
rect 266354 474716 266360 474728
rect 266412 474716 266418 474768
rect 248046 470568 248052 470620
rect 248104 470608 248110 470620
rect 579982 470608 579988 470620
rect 248104 470580 579988 470608
rect 248104 470568 248110 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 266446 462380 266452 462392
rect 3292 462352 266452 462380
rect 3292 462340 3298 462352
rect 266446 462340 266452 462352
rect 266504 462340 266510 462392
rect 246850 456764 246856 456816
rect 246908 456804 246914 456816
rect 580166 456804 580172 456816
rect 246908 456776 580172 456804
rect 246908 456764 246914 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 266538 448576 266544 448588
rect 3200 448548 266544 448576
rect 3200 448536 3206 448548
rect 266538 448536 266544 448548
rect 266596 448536 266602 448588
rect 246758 430584 246764 430636
rect 246816 430624 246822 430636
rect 580166 430624 580172 430636
rect 246816 430596 580172 430624
rect 246816 430584 246822 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 267734 422328 267740 422340
rect 3476 422300 267740 422328
rect 3476 422288 3482 422300
rect 267734 422288 267740 422300
rect 267792 422288 267798 422340
rect 246666 418140 246672 418192
rect 246724 418180 246730 418192
rect 580166 418180 580172 418192
rect 246724 418152 580172 418180
rect 246724 418140 246730 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 267826 409884 267832 409896
rect 3200 409856 267832 409884
rect 3200 409844 3206 409856
rect 267826 409844 267832 409856
rect 267884 409844 267890 409896
rect 245562 404336 245568 404388
rect 245620 404376 245626 404388
rect 580166 404376 580172 404388
rect 245620 404348 580172 404376
rect 245620 404336 245626 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 268010 397508 268016 397520
rect 3476 397480 268016 397508
rect 3476 397468 3482 397480
rect 268010 397468 268016 397480
rect 268068 397468 268074 397520
rect 242158 391756 242164 391808
rect 242216 391796 242222 391808
rect 259730 391796 259736 391808
rect 242216 391768 259736 391796
rect 242216 391756 242222 391768
rect 259730 391756 259736 391768
rect 259788 391756 259794 391808
rect 262585 391799 262643 391805
rect 262585 391765 262597 391799
rect 262631 391796 262643 391799
rect 269758 391796 269764 391808
rect 262631 391768 269764 391796
rect 262631 391765 262643 391768
rect 262585 391759 262643 391765
rect 269758 391756 269764 391768
rect 269816 391756 269822 391808
rect 255682 391688 255688 391740
rect 255740 391728 255746 391740
rect 271138 391728 271144 391740
rect 255740 391700 271144 391728
rect 255740 391688 255746 391700
rect 271138 391688 271144 391700
rect 271196 391688 271202 391740
rect 256602 391552 256608 391604
rect 256660 391592 256666 391604
rect 273898 391592 273904 391604
rect 256660 391564 273904 391592
rect 256660 391552 256666 391564
rect 273898 391552 273904 391564
rect 273956 391552 273962 391604
rect 254578 391484 254584 391536
rect 254636 391524 254642 391536
rect 262585 391527 262643 391533
rect 262585 391524 262597 391527
rect 254636 391496 262597 391524
rect 254636 391484 254642 391496
rect 262585 391493 262597 391496
rect 262631 391493 262643 391527
rect 262585 391487 262643 391493
rect 240778 391416 240784 391468
rect 240836 391456 240842 391468
rect 258626 391456 258632 391468
rect 240836 391428 258632 391456
rect 240836 391416 240842 391428
rect 258626 391416 258632 391428
rect 258684 391416 258690 391468
rect 238018 391348 238024 391400
rect 238076 391388 238082 391400
rect 257614 391388 257620 391400
rect 238076 391360 257620 391388
rect 238076 391348 238082 391360
rect 257614 391348 257620 391360
rect 257672 391348 257678 391400
rect 252002 391280 252008 391332
rect 252060 391320 252066 391332
rect 280798 391320 280804 391332
rect 252060 391292 280804 391320
rect 252060 391280 252066 391292
rect 280798 391280 280804 391292
rect 280856 391280 280862 391332
rect 253474 391212 253480 391264
rect 253532 391252 253538 391264
rect 282178 391252 282184 391264
rect 253532 391224 282184 391252
rect 253532 391212 253538 391224
rect 282178 391212 282184 391224
rect 282236 391212 282242 391264
rect 242802 390464 242808 390516
rect 242860 390504 242866 390516
rect 242860 390476 253934 390504
rect 242860 390464 242866 390476
rect 245930 390396 245936 390448
rect 245988 390436 245994 390448
rect 246758 390436 246764 390448
rect 245988 390408 246764 390436
rect 245988 390396 245994 390408
rect 246758 390396 246764 390408
rect 246816 390396 246822 390448
rect 247402 390396 247408 390448
rect 247460 390436 247466 390448
rect 248046 390436 248052 390448
rect 247460 390408 248052 390436
rect 247460 390396 247466 390408
rect 248046 390396 248052 390408
rect 248104 390396 248110 390448
rect 248966 390396 248972 390448
rect 249024 390436 249030 390448
rect 249518 390436 249524 390448
rect 249024 390408 249524 390436
rect 249024 390396 249030 390408
rect 249518 390396 249524 390408
rect 249576 390396 249582 390448
rect 250070 390396 250076 390448
rect 250128 390436 250134 390448
rect 250714 390436 250720 390448
rect 250128 390408 250720 390436
rect 250128 390396 250134 390408
rect 250714 390396 250720 390408
rect 250772 390396 250778 390448
rect 251910 390396 251916 390448
rect 251968 390436 251974 390448
rect 252278 390436 252284 390448
rect 251968 390408 252284 390436
rect 251968 390396 251974 390408
rect 252278 390396 252284 390408
rect 252336 390396 252342 390448
rect 253014 390396 253020 390448
rect 253072 390436 253078 390448
rect 253750 390436 253756 390448
rect 253072 390408 253756 390436
rect 253072 390396 253078 390408
rect 253750 390396 253756 390408
rect 253808 390396 253814 390448
rect 243998 390328 244004 390380
rect 244056 390368 244062 390380
rect 244056 390340 244274 390368
rect 244056 390328 244062 390340
rect 244246 390300 244274 390340
rect 249334 390328 249340 390380
rect 249392 390368 249398 390380
rect 249702 390368 249708 390380
rect 249392 390340 249708 390368
rect 249392 390328 249398 390340
rect 249702 390328 249708 390340
rect 249760 390328 249766 390380
rect 250438 390328 250444 390380
rect 250496 390368 250502 390380
rect 250990 390368 250996 390380
rect 250496 390340 250996 390368
rect 250496 390328 250502 390340
rect 250990 390328 250996 390340
rect 251048 390328 251054 390380
rect 251542 390328 251548 390380
rect 251600 390368 251606 390380
rect 252370 390368 252376 390380
rect 251600 390340 252376 390368
rect 251600 390328 251606 390340
rect 252370 390328 252376 390340
rect 252428 390328 252434 390380
rect 253906 390368 253934 390476
rect 257154 390464 257160 390516
rect 257212 390504 257218 390516
rect 257982 390504 257988 390516
rect 257212 390476 257988 390504
rect 257212 390464 257218 390476
rect 257982 390464 257988 390476
rect 258040 390464 258046 390516
rect 258166 390464 258172 390516
rect 258224 390504 258230 390516
rect 258994 390504 259000 390516
rect 258224 390476 259000 390504
rect 258224 390464 258230 390476
rect 258994 390464 259000 390476
rect 259052 390464 259058 390516
rect 259638 390464 259644 390516
rect 259696 390504 259702 390516
rect 260466 390504 260472 390516
rect 259696 390476 260472 390504
rect 259696 390464 259702 390476
rect 260466 390464 260472 390476
rect 260524 390464 260530 390516
rect 262214 390464 262220 390516
rect 262272 390504 262278 390516
rect 262766 390504 262772 390516
rect 262272 390476 262772 390504
rect 262272 390464 262278 390476
rect 262766 390464 262772 390476
rect 262824 390464 262830 390516
rect 265158 390464 265164 390516
rect 265216 390504 265222 390516
rect 266078 390504 266084 390516
rect 265216 390476 266084 390504
rect 265216 390464 265222 390476
rect 266078 390464 266084 390476
rect 266136 390464 266142 390516
rect 266446 390464 266452 390516
rect 266504 390504 266510 390516
rect 267274 390504 267280 390516
rect 266504 390476 267280 390504
rect 266504 390464 266510 390476
rect 267274 390464 267280 390476
rect 267332 390464 267338 390516
rect 267826 390464 267832 390516
rect 267884 390504 267890 390516
rect 268378 390504 268384 390516
rect 267884 390476 268384 390504
rect 267884 390464 267890 390476
rect 268378 390464 268384 390476
rect 268436 390464 268442 390516
rect 280890 390464 280896 390516
rect 280948 390504 280954 390516
rect 291930 390504 291936 390516
rect 280948 390476 291936 390504
rect 280948 390464 280954 390476
rect 291930 390464 291936 390476
rect 291988 390464 291994 390516
rect 254210 390396 254216 390448
rect 254268 390436 254274 390448
rect 255130 390436 255136 390448
rect 254268 390408 255136 390436
rect 254268 390396 254274 390408
rect 255130 390396 255136 390408
rect 255188 390396 255194 390448
rect 256050 390396 256056 390448
rect 256108 390436 256114 390448
rect 256510 390436 256516 390448
rect 256108 390408 256516 390436
rect 256108 390396 256114 390408
rect 256510 390396 256516 390408
rect 256568 390396 256574 390448
rect 256605 390439 256663 390445
rect 256605 390405 256617 390439
rect 256651 390436 256663 390439
rect 540422 390436 540428 390448
rect 256651 390408 540428 390436
rect 256651 390405 256663 390408
rect 256605 390399 256663 390405
rect 540422 390396 540428 390408
rect 540480 390396 540486 390448
rect 544470 390368 544476 390380
rect 253906 390340 544476 390368
rect 544470 390328 544476 390340
rect 544528 390328 544534 390380
rect 547230 390300 547236 390312
rect 244246 390272 547236 390300
rect 547230 390260 547236 390272
rect 547288 390260 547294 390312
rect 245194 390192 245200 390244
rect 245252 390232 245258 390244
rect 245252 390204 287054 390232
rect 245252 390192 245258 390204
rect 241790 390124 241796 390176
rect 241848 390164 241854 390176
rect 281077 390167 281135 390173
rect 281077 390164 281089 390167
rect 241848 390136 281089 390164
rect 241848 390124 241854 390136
rect 281077 390133 281089 390136
rect 281123 390133 281135 390167
rect 285122 390164 285128 390176
rect 281077 390127 281135 390133
rect 281184 390136 285128 390164
rect 241422 390056 241428 390108
rect 241480 390096 241486 390108
rect 281184 390096 281212 390136
rect 285122 390124 285128 390136
rect 285180 390124 285186 390176
rect 285217 390167 285275 390173
rect 285217 390133 285229 390167
rect 285263 390164 285275 390167
rect 286502 390164 286508 390176
rect 285263 390136 286508 390164
rect 285263 390133 285275 390136
rect 285217 390127 285275 390133
rect 286502 390124 286508 390136
rect 286560 390124 286566 390176
rect 287026 390164 287054 390204
rect 289078 390164 289084 390176
rect 287026 390136 289084 390164
rect 289078 390124 289084 390136
rect 289136 390124 289142 390176
rect 284941 390099 284999 390105
rect 284941 390096 284953 390099
rect 241480 390068 281212 390096
rect 281276 390068 284953 390096
rect 241480 390056 241486 390068
rect 152458 389988 152464 390040
rect 152516 390028 152522 390040
rect 277486 390028 277492 390040
rect 152516 390000 277492 390028
rect 152516 389988 152522 390000
rect 277486 389988 277492 390000
rect 277544 389988 277550 390040
rect 281077 390031 281135 390037
rect 281077 389997 281089 390031
rect 281123 390028 281135 390031
rect 281276 390028 281304 390068
rect 284941 390065 284953 390068
rect 284987 390065 284999 390099
rect 284941 390059 284999 390065
rect 285030 390056 285036 390108
rect 285088 390096 285094 390108
rect 292206 390096 292212 390108
rect 285088 390068 292212 390096
rect 285088 390056 285094 390068
rect 292206 390056 292212 390068
rect 292264 390056 292270 390108
rect 281123 390000 281304 390028
rect 281123 389997 281135 390000
rect 281077 389991 281135 389997
rect 282362 389988 282368 390040
rect 282420 390028 282426 390040
rect 292022 390028 292028 390040
rect 282420 390000 292028 390028
rect 282420 389988 282426 390000
rect 292022 389988 292028 390000
rect 292080 389988 292086 390040
rect 248138 389920 248144 389972
rect 248196 389960 248202 389972
rect 248322 389960 248328 389972
rect 248196 389932 248328 389960
rect 248196 389920 248202 389932
rect 248322 389920 248328 389932
rect 248380 389920 248386 389972
rect 249061 389963 249119 389969
rect 249061 389929 249073 389963
rect 249107 389960 249119 389963
rect 395338 389960 395344 389972
rect 249107 389932 395344 389960
rect 249107 389929 249119 389932
rect 249061 389923 249119 389929
rect 395338 389920 395344 389932
rect 395396 389920 395402 389972
rect 40770 389852 40776 389904
rect 40828 389892 40834 389904
rect 273990 389892 273996 389904
rect 40828 389864 273996 389892
rect 40828 389852 40834 389864
rect 273990 389852 273996 389864
rect 274048 389852 274054 389904
rect 281350 389852 281356 389904
rect 281408 389892 281414 389904
rect 291838 389892 291844 389904
rect 281408 389864 291844 389892
rect 281408 389852 281414 389864
rect 291838 389852 291844 389864
rect 291896 389852 291902 389904
rect 39390 389784 39396 389836
rect 39448 389824 39454 389836
rect 272886 389824 272892 389836
rect 39448 389796 272892 389824
rect 39448 389784 39454 389796
rect 272886 389784 272892 389796
rect 272944 389784 272950 389836
rect 281258 389784 281264 389836
rect 281316 389824 281322 389836
rect 296070 389824 296076 389836
rect 281316 389796 296076 389824
rect 281316 389784 281322 389796
rect 296070 389784 296076 389796
rect 296128 389784 296134 389836
rect 36630 389716 36636 389768
rect 36688 389756 36694 389768
rect 271874 389756 271880 389768
rect 36688 389728 271880 389756
rect 36688 389716 36694 389728
rect 271874 389716 271880 389728
rect 271932 389716 271938 389768
rect 279694 389716 279700 389768
rect 279752 389756 279758 389768
rect 288066 389756 288072 389768
rect 279752 389728 288072 389756
rect 279752 389716 279758 389728
rect 288066 389716 288072 389728
rect 288124 389716 288130 389768
rect 35250 389648 35256 389700
rect 35308 389688 35314 389700
rect 270586 389688 270592 389700
rect 35308 389660 270592 389688
rect 35308 389648 35314 389660
rect 270586 389648 270592 389660
rect 270644 389648 270650 389700
rect 282730 389648 282736 389700
rect 282788 389688 282794 389700
rect 292114 389688 292120 389700
rect 282788 389660 292120 389688
rect 282788 389648 282794 389660
rect 292114 389648 292120 389660
rect 292172 389648 292178 389700
rect 33778 389580 33784 389632
rect 33836 389620 33842 389632
rect 275094 389620 275100 389632
rect 33836 389592 275100 389620
rect 33836 389580 33842 389592
rect 275094 389580 275100 389592
rect 275152 389580 275158 389632
rect 278682 389580 278688 389632
rect 278740 389620 278746 389632
rect 294690 389620 294696 389632
rect 278740 389592 294696 389620
rect 278740 389580 278746 389592
rect 294690 389580 294696 389592
rect 294748 389580 294754 389632
rect 35158 389512 35164 389564
rect 35216 389552 35222 389564
rect 276290 389552 276296 389564
rect 35216 389524 276296 389552
rect 35216 389512 35222 389524
rect 276290 389512 276296 389524
rect 276348 389512 276354 389564
rect 280062 389512 280068 389564
rect 280120 389552 280126 389564
rect 418890 389552 418896 389564
rect 280120 389524 418896 389552
rect 280120 389512 280126 389524
rect 418890 389512 418896 389524
rect 418948 389512 418954 389564
rect 15838 389444 15844 389496
rect 15896 389484 15902 389496
rect 269482 389484 269488 389496
rect 15896 389456 269488 389484
rect 15896 389444 15902 389456
rect 269482 389444 269488 389456
rect 269540 389444 269546 389496
rect 284570 389444 284576 389496
rect 284628 389484 284634 389496
rect 439682 389484 439688 389496
rect 284628 389456 439688 389484
rect 284628 389444 284634 389456
rect 439682 389444 439688 389456
rect 439740 389444 439746 389496
rect 21358 389376 21364 389428
rect 21416 389416 21422 389428
rect 277026 389416 277032 389428
rect 21416 389388 277032 389416
rect 21416 389376 21422 389388
rect 277026 389376 277032 389388
rect 277084 389376 277090 389428
rect 282822 389376 282828 389428
rect 282880 389416 282886 389428
rect 438302 389416 438308 389428
rect 282880 389388 438308 389416
rect 282880 389376 282886 389388
rect 438302 389376 438308 389388
rect 438360 389376 438366 389428
rect 242526 389308 242532 389360
rect 242584 389348 242590 389360
rect 256605 389351 256663 389357
rect 256605 389348 256617 389351
rect 242584 389320 256617 389348
rect 242584 389308 242590 389320
rect 256605 389317 256617 389320
rect 256651 389317 256663 389351
rect 256605 389311 256663 389317
rect 279326 389308 279332 389360
rect 279384 389348 279390 389360
rect 288158 389348 288164 389360
rect 279384 389320 288164 389348
rect 279384 389308 279390 389320
rect 288158 389308 288164 389320
rect 288216 389308 288222 389360
rect 240042 389240 240048 389292
rect 240100 389280 240106 389292
rect 249061 389283 249119 389289
rect 249061 389280 249073 389283
rect 240100 389252 249073 389280
rect 240100 389240 240106 389252
rect 249061 389249 249073 389252
rect 249107 389249 249119 389283
rect 249061 389243 249119 389249
rect 284202 389240 284208 389292
rect 284260 389280 284266 389292
rect 297358 389280 297364 389292
rect 284260 389252 297364 389280
rect 284260 389240 284266 389252
rect 297358 389240 297364 389252
rect 297416 389240 297422 389292
rect 283466 389172 283472 389224
rect 283524 389212 283530 389224
rect 293218 389212 293224 389224
rect 283524 389184 293224 389212
rect 283524 389172 283530 389184
rect 293218 389172 293224 389184
rect 293276 389172 293282 389224
rect 32490 389104 32496 389156
rect 32548 389144 32554 389156
rect 272150 389144 272156 389156
rect 32548 389116 272156 389144
rect 32548 389104 32554 389116
rect 272150 389104 272156 389116
rect 272208 389104 272214 389156
rect 236546 389036 236552 389088
rect 236604 389076 236610 389088
rect 295978 389076 295984 389088
rect 236604 389048 295984 389076
rect 236604 389036 236610 389048
rect 295978 389036 295984 389048
rect 296036 389036 296042 389088
rect 235810 388968 235816 389020
rect 235868 389008 235874 389020
rect 300118 389008 300124 389020
rect 235868 388980 300124 389008
rect 235868 388968 235874 388980
rect 300118 388968 300124 388980
rect 300176 388968 300182 389020
rect 236914 388900 236920 388952
rect 236972 388940 236978 388952
rect 302878 388940 302884 388952
rect 236972 388912 302884 388940
rect 236972 388900 236978 388912
rect 302878 388900 302884 388912
rect 302936 388900 302942 388952
rect 237650 388832 237656 388884
rect 237708 388872 237714 388884
rect 313918 388872 313924 388884
rect 237708 388844 313924 388872
rect 237708 388832 237714 388844
rect 313918 388832 313924 388844
rect 313976 388832 313982 388884
rect 235442 388764 235448 388816
rect 235500 388804 235506 388816
rect 318058 388804 318064 388816
rect 235500 388776 318064 388804
rect 235500 388764 235506 388776
rect 318058 388764 318064 388776
rect 318116 388764 318122 388816
rect 243630 388696 243636 388748
rect 243688 388736 243694 388748
rect 443638 388736 443644 388748
rect 243688 388708 443644 388736
rect 243688 388696 243694 388708
rect 443638 388696 443644 388708
rect 443696 388696 443702 388748
rect 33870 388628 33876 388680
rect 33928 388668 33934 388680
rect 270218 388668 270224 388680
rect 33928 388640 270224 388668
rect 33928 388628 33934 388640
rect 270218 388628 270224 388640
rect 270276 388628 270282 388680
rect 29638 388560 29644 388612
rect 29696 388600 29702 388612
rect 273622 388600 273628 388612
rect 29696 388572 273628 388600
rect 29696 388560 29702 388572
rect 273622 388560 273628 388572
rect 273680 388560 273686 388612
rect 21450 388492 21456 388544
rect 21508 388532 21514 388544
rect 272518 388532 272524 388544
rect 21508 388504 272524 388532
rect 21508 388492 21514 388504
rect 272518 388492 272524 388504
rect 272576 388492 272582 388544
rect 18690 388424 18696 388476
rect 18748 388464 18754 388476
rect 271322 388464 271328 388476
rect 18748 388436 271328 388464
rect 18748 388424 18754 388436
rect 271322 388424 271328 388436
rect 271380 388424 271386 388476
rect 17310 388356 17316 388408
rect 17368 388396 17374 388408
rect 270954 388396 270960 388408
rect 17368 388368 270960 388396
rect 17368 388356 17374 388368
rect 270954 388356 270960 388368
rect 271012 388356 271018 388408
rect 14642 388288 14648 388340
rect 14700 388328 14706 388340
rect 269850 388328 269856 388340
rect 14700 388300 269856 388328
rect 14700 388288 14706 388300
rect 269850 388288 269856 388300
rect 269908 388288 269914 388340
rect 18598 388220 18604 388272
rect 18656 388260 18662 388272
rect 276014 388260 276020 388272
rect 18656 388232 276020 388260
rect 18656 388220 18662 388232
rect 276014 388220 276020 388232
rect 276072 388220 276078 388272
rect 14550 388152 14556 388204
rect 14608 388192 14614 388204
rect 273484 388192 273490 388204
rect 14608 388164 273490 388192
rect 14608 388152 14614 388164
rect 273484 388152 273490 388164
rect 273542 388152 273548 388204
rect 7558 388084 7564 388136
rect 7616 388124 7622 388136
rect 268976 388124 268982 388136
rect 7616 388096 268982 388124
rect 7616 388084 7622 388096
rect 268976 388084 268982 388096
rect 269034 388084 269040 388136
rect 277992 388084 277998 388136
rect 278050 388124 278056 388136
rect 447778 388124 447784 388136
rect 278050 388096 447784 388124
rect 278050 388084 278056 388096
rect 447778 388084 447784 388096
rect 447836 388084 447842 388136
rect 11790 388016 11796 388068
rect 11848 388056 11854 388068
rect 274358 388056 274364 388068
rect 11848 388028 274364 388056
rect 11848 388016 11854 388028
rect 274358 388016 274364 388028
rect 274416 388016 274422 388068
rect 278590 388016 278596 388068
rect 278648 388056 278654 388068
rect 449158 388056 449164 388068
rect 278648 388028 449164 388056
rect 278648 388016 278654 388028
rect 449158 388016 449164 388028
rect 449216 388016 449222 388068
rect 4798 387948 4804 388000
rect 4856 387988 4862 388000
rect 275462 387988 275468 388000
rect 4856 387960 275468 387988
rect 4856 387948 4862 387960
rect 275462 387948 275468 387960
rect 275520 387948 275526 388000
rect 280522 387948 280528 388000
rect 280580 387988 280586 388000
rect 481634 387988 481640 388000
rect 280580 387960 481640 387988
rect 280580 387948 280586 387960
rect 481634 387948 481640 387960
rect 481692 387948 481698 388000
rect 3418 387880 3424 387932
rect 3476 387920 3482 387932
rect 276658 387920 276664 387932
rect 3476 387892 276664 387920
rect 3476 387880 3482 387892
rect 276658 387880 276664 387892
rect 276716 387880 276722 387932
rect 281994 387880 282000 387932
rect 282052 387920 282058 387932
rect 485774 387920 485780 387932
rect 282052 387892 485780 387920
rect 282052 387880 282058 387892
rect 485774 387880 485780 387892
rect 485832 387880 485838 387932
rect 243262 387812 243268 387864
rect 243320 387852 243326 387864
rect 537478 387852 537484 387864
rect 243320 387824 537484 387852
rect 243320 387812 243326 387824
rect 537478 387812 537484 387824
rect 537536 387812 537542 387864
rect 263594 387744 263600 387796
rect 263652 387784 263658 387796
rect 263870 387784 263876 387796
rect 263652 387756 263876 387784
rect 263652 387744 263658 387756
rect 263870 387744 263876 387756
rect 263928 387744 263934 387796
rect 237282 387308 237288 387320
rect 237243 387280 237288 387308
rect 237282 387268 237288 387280
rect 237340 387268 237346 387320
rect 238018 387308 238024 387320
rect 237979 387280 238024 387308
rect 238018 387268 238024 387280
rect 238076 387268 238082 387320
rect 238662 387268 238668 387320
rect 238720 387308 238726 387320
rect 239122 387308 239128 387320
rect 238720 387268 238754 387308
rect 239083 387280 239128 387308
rect 239122 387268 239128 387280
rect 239180 387268 239186 387320
rect 239950 387308 239956 387320
rect 239911 387280 239956 387308
rect 239950 387268 239956 387280
rect 240008 387268 240014 387320
rect 241054 387308 241060 387320
rect 241015 387280 241060 387308
rect 241054 387268 241060 387280
rect 241112 387268 241118 387320
rect 242158 387308 242164 387320
rect 242119 387280 242164 387308
rect 242158 387268 242164 387280
rect 242216 387268 242222 387320
rect 244274 387308 244280 387320
rect 244235 387280 244280 387308
rect 244274 387268 244280 387280
rect 244332 387268 244338 387320
rect 244826 387308 244832 387320
rect 244787 387280 244832 387308
rect 244826 387268 244832 387280
rect 244884 387268 244890 387320
rect 269114 387308 269120 387320
rect 269075 387280 269120 387308
rect 269114 387268 269120 387280
rect 269172 387268 269178 387320
rect 274726 387308 274732 387320
rect 274687 387280 274732 387308
rect 274726 387268 274732 387280
rect 274784 387268 274790 387320
rect 283834 387308 283840 387320
rect 283795 387280 283840 387308
rect 283834 387268 283840 387280
rect 283892 387268 283898 387320
rect 238726 387172 238754 387268
rect 580350 387172 580356 387184
rect 238726 387144 580356 387172
rect 580350 387132 580356 387144
rect 580408 387132 580414 387184
rect 17218 387064 17224 387116
rect 17276 387104 17282 387116
rect 274729 387107 274787 387113
rect 274729 387104 274741 387107
rect 17276 387076 274741 387104
rect 17276 387064 17282 387076
rect 274729 387073 274741 387076
rect 274775 387073 274787 387107
rect 274729 387067 274787 387073
rect 3510 386996 3516 387048
rect 3568 387036 3574 387048
rect 269117 387039 269175 387045
rect 269117 387036 269129 387039
rect 3568 387008 269129 387036
rect 3568 386996 3574 387008
rect 269117 387005 269129 387008
rect 269163 387005 269175 387039
rect 269117 386999 269175 387005
rect 288342 386996 288348 387048
rect 288400 387036 288406 387048
rect 471238 387036 471244 387048
rect 288400 387008 471244 387036
rect 288400 386996 288406 387008
rect 471238 386996 471244 387008
rect 471296 386996 471302 387048
rect 237285 386971 237343 386977
rect 237285 386937 237297 386971
rect 237331 386968 237343 386971
rect 555418 386968 555424 386980
rect 237331 386940 555424 386968
rect 237331 386937 237343 386940
rect 237285 386931 237343 386937
rect 555418 386928 555424 386940
rect 555476 386928 555482 386980
rect 244829 386903 244887 386909
rect 244829 386869 244841 386903
rect 244875 386900 244887 386903
rect 580902 386900 580908 386912
rect 244875 386872 580908 386900
rect 244875 386869 244887 386872
rect 244829 386863 244887 386869
rect 580902 386860 580908 386872
rect 580960 386860 580966 386912
rect 244277 386835 244335 386841
rect 244277 386801 244289 386835
rect 244323 386832 244335 386835
rect 580718 386832 580724 386844
rect 244323 386804 580724 386832
rect 244323 386801 244335 386804
rect 244277 386795 244335 386801
rect 580718 386792 580724 386804
rect 580776 386792 580782 386844
rect 242161 386767 242219 386773
rect 242161 386733 242173 386767
rect 242207 386764 242219 386767
rect 580810 386764 580816 386776
rect 242207 386736 580816 386764
rect 242207 386733 242219 386736
rect 242161 386727 242219 386733
rect 580810 386724 580816 386736
rect 580868 386724 580874 386776
rect 241057 386699 241115 386705
rect 241057 386665 241069 386699
rect 241103 386696 241115 386699
rect 580626 386696 580632 386708
rect 241103 386668 580632 386696
rect 241103 386665 241115 386668
rect 241057 386659 241115 386665
rect 580626 386656 580632 386668
rect 580684 386656 580690 386708
rect 239125 386631 239183 386637
rect 239125 386597 239137 386631
rect 239171 386628 239183 386631
rect 580442 386628 580448 386640
rect 239171 386600 580448 386628
rect 239171 386597 239183 386600
rect 239125 386591 239183 386597
rect 580442 386588 580448 386600
rect 580500 386588 580506 386640
rect 239953 386563 240011 386569
rect 239953 386529 239965 386563
rect 239999 386560 240011 386563
rect 580534 386560 580540 386572
rect 239999 386532 580540 386560
rect 239999 386529 240011 386532
rect 239953 386523 240011 386529
rect 580534 386520 580540 386532
rect 580592 386520 580598 386572
rect 238021 386495 238079 386501
rect 238021 386461 238033 386495
rect 238067 386492 238079 386495
rect 580258 386492 580264 386504
rect 238067 386464 580264 386492
rect 238067 386461 238079 386464
rect 238021 386455 238079 386461
rect 580258 386452 580264 386464
rect 580316 386452 580322 386504
rect 283837 386427 283895 386433
rect 283837 386393 283849 386427
rect 283883 386424 283895 386427
rect 293310 386424 293316 386436
rect 283883 386396 293316 386424
rect 283883 386393 283895 386396
rect 283837 386387 283895 386393
rect 293310 386384 293316 386396
rect 293368 386384 293374 386436
rect 288342 385024 288348 385076
rect 288400 385064 288406 385076
rect 298738 385064 298744 385076
rect 288400 385036 298744 385064
rect 288400 385024 288406 385036
rect 298738 385024 298744 385036
rect 298796 385024 298802 385076
rect 288342 383664 288348 383716
rect 288400 383704 288406 383716
rect 468478 383704 468484 383716
rect 288400 383676 468484 383704
rect 288400 383664 288406 383676
rect 468478 383664 468484 383676
rect 468536 383664 468542 383716
rect 287422 381692 287428 381744
rect 287480 381732 287486 381744
rect 294782 381732 294788 381744
rect 287480 381704 294788 381732
rect 287480 381692 287486 381704
rect 294782 381692 294788 381704
rect 294840 381692 294846 381744
rect 288342 379516 288348 379568
rect 288400 379556 288406 379568
rect 465718 379556 465724 379568
rect 288400 379528 465724 379556
rect 288400 379516 288406 379528
rect 465718 379516 465724 379528
rect 465776 379516 465782 379568
rect 288342 378156 288348 378208
rect 288400 378196 288406 378208
rect 297450 378196 297456 378208
rect 288400 378168 297456 378196
rect 288400 378156 288406 378168
rect 297450 378156 297456 378168
rect 297508 378156 297514 378208
rect 287422 376728 287428 376780
rect 287480 376768 287486 376780
rect 293402 376768 293408 376780
rect 287480 376740 293408 376768
rect 287480 376728 287486 376740
rect 293402 376728 293408 376740
rect 293460 376728 293466 376780
rect 287606 375368 287612 375420
rect 287664 375408 287670 375420
rect 293494 375408 293500 375420
rect 287664 375380 293500 375408
rect 287664 375368 287670 375380
rect 293494 375368 293500 375380
rect 293552 375368 293558 375420
rect 288342 374144 288348 374196
rect 288400 374184 288406 374196
rect 293586 374184 293592 374196
rect 288400 374156 293592 374184
rect 288400 374144 288406 374156
rect 293586 374144 293592 374156
rect 293644 374144 293650 374196
rect 287790 371628 287796 371680
rect 287848 371668 287854 371680
rect 292298 371668 292304 371680
rect 287848 371640 292304 371668
rect 287848 371628 287854 371640
rect 292298 371628 292304 371640
rect 292356 371628 292362 371680
rect 3326 371560 3332 371612
rect 3384 371600 3390 371612
rect 7558 371600 7564 371612
rect 3384 371572 7564 371600
rect 3384 371560 3390 371572
rect 7558 371560 7564 371572
rect 7616 371560 7622 371612
rect 287606 370540 287612 370592
rect 287664 370580 287670 370592
rect 290550 370580 290556 370592
rect 287664 370552 290556 370580
rect 287664 370540 287670 370552
rect 290550 370540 290556 370552
rect 290608 370540 290614 370592
rect 288342 368500 288348 368552
rect 288400 368540 288406 368552
rect 446398 368540 446404 368552
rect 288400 368512 446404 368540
rect 288400 368500 288406 368512
rect 446398 368500 446404 368512
rect 446456 368500 446462 368552
rect 287974 367072 287980 367124
rect 288032 367112 288038 367124
rect 297542 367112 297548 367124
rect 288032 367084 297548 367112
rect 288032 367072 288038 367084
rect 297542 367072 297548 367084
rect 297600 367072 297606 367124
rect 287606 365712 287612 365764
rect 287664 365752 287670 365764
rect 296162 365752 296168 365764
rect 287664 365724 296168 365752
rect 287664 365712 287670 365724
rect 296162 365712 296168 365724
rect 296220 365712 296226 365764
rect 289078 365644 289084 365696
rect 289136 365684 289142 365696
rect 580166 365684 580172 365696
rect 289136 365656 580172 365684
rect 289136 365644 289142 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 288342 364352 288348 364404
rect 288400 364392 288406 364404
rect 296254 364392 296260 364404
rect 288400 364364 296260 364392
rect 288400 364352 288406 364364
rect 296254 364352 296260 364364
rect 296312 364352 296318 364404
rect 287606 362312 287612 362364
rect 287664 362352 287670 362364
rect 296346 362352 296352 362364
rect 287664 362324 296352 362352
rect 287664 362312 287670 362324
rect 296346 362312 296352 362324
rect 296404 362312 296410 362364
rect 287606 360612 287612 360664
rect 287664 360652 287670 360664
rect 296438 360652 296444 360664
rect 287664 360624 296444 360652
rect 287664 360612 287670 360624
rect 296438 360612 296444 360624
rect 296496 360612 296502 360664
rect 287606 358980 287612 359032
rect 287664 359020 287670 359032
rect 289446 359020 289452 359032
rect 287664 358992 289452 359020
rect 287664 358980 287670 358992
rect 289446 358980 289452 358992
rect 289504 358980 289510 359032
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 15838 358748 15844 358760
rect 3384 358720 15844 358748
rect 3384 358708 3390 358720
rect 15838 358708 15844 358720
rect 15896 358708 15902 358760
rect 288342 357416 288348 357468
rect 288400 357456 288406 357468
rect 473998 357456 474004 357468
rect 288400 357428 474004 357456
rect 288400 357416 288406 357428
rect 473998 357416 474004 357428
rect 474056 357416 474062 357468
rect 287790 356056 287796 356108
rect 287848 356096 287854 356108
rect 298922 356096 298928 356108
rect 287848 356068 298928 356096
rect 287848 356056 287854 356068
rect 298922 356056 298928 356068
rect 298980 356056 298986 356108
rect 288342 354696 288348 354748
rect 288400 354736 288406 354748
rect 298830 354736 298836 354748
rect 288400 354708 298836 354736
rect 288400 354696 288406 354708
rect 298830 354696 298836 354708
rect 298888 354696 298894 354748
rect 287514 351908 287520 351960
rect 287572 351948 287578 351960
rect 472618 351948 472624 351960
rect 287572 351920 472624 351948
rect 287572 351908 287578 351920
rect 472618 351908 472624 351920
rect 472676 351908 472682 351960
rect 287238 351432 287244 351484
rect 287296 351472 287302 351484
rect 294874 351472 294880 351484
rect 287296 351444 294880 351472
rect 287296 351432 287302 351444
rect 294874 351432 294880 351444
rect 294932 351432 294938 351484
rect 232130 349800 232136 349852
rect 232188 349840 232194 349852
rect 232866 349840 232872 349852
rect 232188 349812 232872 349840
rect 232188 349800 232194 349812
rect 232866 349800 232872 349812
rect 232924 349800 232930 349852
rect 288342 349120 288348 349172
rect 288400 349160 288406 349172
rect 467098 349160 467104 349172
rect 288400 349132 467104 349160
rect 288400 349120 288406 349132
rect 467098 349120 467104 349132
rect 467156 349120 467162 349172
rect 287974 347760 287980 347812
rect 288032 347800 288038 347812
rect 299014 347800 299020 347812
rect 288032 347772 299020 347800
rect 288032 347760 288038 347772
rect 299014 347760 299020 347772
rect 299072 347760 299078 347812
rect 287974 346536 287980 346588
rect 288032 346576 288038 346588
rect 294966 346576 294972 346588
rect 288032 346548 294972 346576
rect 288032 346536 288038 346548
rect 294966 346536 294972 346548
rect 295024 346536 295030 346588
rect 288342 345040 288348 345092
rect 288400 345080 288406 345092
rect 295058 345080 295064 345092
rect 288400 345052 295064 345080
rect 288400 345040 288406 345052
rect 295058 345040 295064 345052
rect 295116 345040 295122 345092
rect 288342 342252 288348 342304
rect 288400 342292 288406 342304
rect 464338 342292 464344 342304
rect 288400 342264 464344 342292
rect 288400 342252 288406 342264
rect 464338 342252 464344 342264
rect 464396 342252 464402 342304
rect 288342 340892 288348 340944
rect 288400 340932 288406 340944
rect 297726 340932 297732 340944
rect 288400 340904 297732 340932
rect 288400 340892 288406 340904
rect 297726 340892 297732 340904
rect 297784 340892 297790 340944
rect 287790 339464 287796 339516
rect 287848 339504 287854 339516
rect 292390 339504 292396 339516
rect 287848 339476 292396 339504
rect 287848 339464 287854 339476
rect 292390 339464 292396 339476
rect 292448 339464 292454 339516
rect 446398 338716 446404 338768
rect 446456 338756 446462 338768
rect 488534 338756 488540 338768
rect 446456 338728 488540 338756
rect 446456 338716 446462 338728
rect 488534 338716 488540 338728
rect 488592 338716 488598 338768
rect 234522 338648 234528 338700
rect 234580 338688 234586 338700
rect 467834 338688 467840 338700
rect 234580 338660 467840 338688
rect 234580 338648 234586 338660
rect 467834 338648 467840 338660
rect 467892 338648 467898 338700
rect 232130 338580 232136 338632
rect 232188 338620 232194 338632
rect 297634 338620 297640 338632
rect 232188 338592 297640 338620
rect 232188 338580 232194 338592
rect 297634 338580 297640 338592
rect 297692 338580 297698 338632
rect 232866 338512 232872 338564
rect 232924 338552 232930 338564
rect 289538 338552 289544 338564
rect 232924 338524 289544 338552
rect 232924 338512 232930 338524
rect 289538 338512 289544 338524
rect 289596 338512 289602 338564
rect 278869 338283 278927 338289
rect 278869 338280 278881 338283
rect 275986 338252 278881 338280
rect 234614 338036 234620 338088
rect 234672 338076 234678 338088
rect 238665 338079 238723 338085
rect 234672 338048 237190 338076
rect 234672 338036 234678 338048
rect 233602 337968 233608 338020
rect 233660 338008 233666 338020
rect 235445 338011 235503 338017
rect 233660 337980 234614 338008
rect 233660 337968 233666 337980
rect 234586 337736 234614 337980
rect 235445 337977 235457 338011
rect 235491 338008 235503 338011
rect 235491 337980 235626 338008
rect 235491 337977 235503 337980
rect 235445 337971 235503 337977
rect 235598 337952 235626 337980
rect 237162 337952 237190 338048
rect 238665 338045 238677 338079
rect 238711 338045 238723 338079
rect 238665 338039 238723 338045
rect 238680 338008 238708 338039
rect 242161 338011 242219 338017
rect 238680 337980 239398 338008
rect 239370 337952 239398 337980
rect 242161 337977 242173 338011
rect 242207 338008 242219 338011
rect 242710 338008 242716 338020
rect 242207 337980 242716 338008
rect 242207 337977 242219 337980
rect 242161 337971 242219 337977
rect 242710 337968 242716 337980
rect 242768 337968 242774 338020
rect 242897 338011 242955 338017
rect 242897 337977 242909 338011
rect 242943 338008 242955 338011
rect 254489 338011 254547 338017
rect 242943 337980 249886 338008
rect 242943 337977 242955 337980
rect 242897 337971 242955 337977
rect 249858 337952 249886 337980
rect 254489 337977 254501 338011
rect 254535 338008 254547 338011
rect 254949 338011 255007 338017
rect 254949 338008 254961 338011
rect 254535 337980 254670 338008
rect 254535 337977 254547 337980
rect 254489 337971 254547 337977
rect 254642 337952 254670 337980
rect 254826 337980 254961 338008
rect 254826 337952 254854 337980
rect 254949 337977 254961 337980
rect 254995 337977 255007 338011
rect 269485 338011 269543 338017
rect 269485 338008 269497 338011
rect 254949 337971 255007 337977
rect 262278 337980 269497 338008
rect 262278 337952 262306 337980
rect 269485 337977 269497 337980
rect 269531 337977 269543 338011
rect 272613 338011 272671 338017
rect 272613 338008 272625 338011
rect 269485 337971 269543 337977
rect 272398 337980 272625 338008
rect 272398 337952 272426 337980
rect 272613 337977 272625 337980
rect 272659 337977 272671 338011
rect 272613 337971 272671 337977
rect 275986 337952 276014 338252
rect 278869 338249 278881 338252
rect 278915 338249 278927 338283
rect 278869 338243 278927 338249
rect 276201 338215 276259 338221
rect 276201 338181 276213 338215
rect 276247 338181 276259 338215
rect 276201 338175 276259 338181
rect 276216 338144 276244 338175
rect 282917 338147 282975 338153
rect 282917 338144 282929 338147
rect 276170 338116 276244 338144
rect 282518 338116 282929 338144
rect 276170 337952 276198 338116
rect 279237 338011 279295 338017
rect 279237 338008 279249 338011
rect 278930 337980 279249 338008
rect 234890 337900 234896 337952
rect 234948 337940 234954 337952
rect 235304 337940 235310 337952
rect 234948 337912 235310 337940
rect 234948 337900 234954 337912
rect 235304 337900 235310 337912
rect 235362 337900 235368 337952
rect 235580 337900 235586 337952
rect 235638 337900 235644 337952
rect 236181 337943 236239 337949
rect 236181 337909 236193 337943
rect 236227 337940 236239 337943
rect 236316 337940 236322 337952
rect 236227 337912 236322 337940
rect 236227 337909 236239 337912
rect 236181 337903 236239 337909
rect 236316 337900 236322 337912
rect 236374 337900 236380 337952
rect 237144 337900 237150 337952
rect 237202 337900 237208 337952
rect 237696 337900 237702 337952
rect 237754 337949 237760 337952
rect 237880 337949 237886 337952
rect 237754 337943 237803 337949
rect 237754 337909 237757 337943
rect 237791 337909 237803 337943
rect 237754 337903 237803 337909
rect 237837 337943 237886 337949
rect 237837 337909 237849 337943
rect 237883 337909 237886 337943
rect 237837 337903 237886 337909
rect 237754 337900 237760 337903
rect 237880 337900 237886 337903
rect 237938 337900 237944 337952
rect 238616 337949 238622 337952
rect 238573 337943 238622 337949
rect 238573 337909 238585 337943
rect 238619 337909 238622 337943
rect 238573 337903 238622 337909
rect 238616 337900 238622 337903
rect 238674 337900 238680 337952
rect 238708 337900 238714 337952
rect 238766 337949 238772 337952
rect 238892 337949 238898 337952
rect 238766 337943 238815 337949
rect 238766 337909 238769 337943
rect 238803 337909 238815 337943
rect 238766 337903 238815 337909
rect 238849 337943 238898 337949
rect 238849 337909 238861 337943
rect 238895 337909 238898 337943
rect 238849 337903 238898 337909
rect 238766 337900 238772 337903
rect 238892 337900 238898 337903
rect 238950 337900 238956 337952
rect 239260 337949 239266 337952
rect 239217 337943 239266 337949
rect 239217 337909 239229 337943
rect 239263 337909 239266 337943
rect 239217 337903 239266 337909
rect 239260 337900 239266 337903
rect 239318 337900 239324 337952
rect 239352 337900 239358 337952
rect 239410 337900 239416 337952
rect 239536 337949 239542 337952
rect 239493 337943 239542 337949
rect 239493 337909 239505 337943
rect 239539 337909 239542 337943
rect 239493 337903 239542 337909
rect 239536 337900 239542 337903
rect 239594 337900 239600 337952
rect 239720 337900 239726 337952
rect 239778 337900 239784 337952
rect 241100 337949 241106 337952
rect 241057 337943 241106 337949
rect 241057 337909 241069 337943
rect 241103 337909 241106 337943
rect 241057 337903 241106 337909
rect 241100 337900 241106 337903
rect 241158 337900 241164 337952
rect 241241 337943 241299 337949
rect 241241 337909 241253 337943
rect 241287 337940 241299 337943
rect 241376 337940 241382 337952
rect 241287 337912 241382 337940
rect 241287 337909 241299 337912
rect 241241 337903 241299 337909
rect 241376 337900 241382 337912
rect 241434 337900 241440 337952
rect 242388 337900 242394 337952
rect 242446 337940 242452 337952
rect 242805 337943 242863 337949
rect 242446 337900 242480 337940
rect 242805 337909 242817 337943
rect 242851 337940 242863 337943
rect 243124 337940 243130 337952
rect 242851 337912 243130 337940
rect 242851 337909 242863 337912
rect 242805 337903 242863 337909
rect 243124 337900 243130 337912
rect 243182 337900 243188 337952
rect 245197 337943 245255 337949
rect 245197 337909 245209 337943
rect 245243 337940 245255 337943
rect 245332 337940 245338 337952
rect 245243 337912 245338 337940
rect 245243 337909 245255 337912
rect 245197 337903 245255 337909
rect 245332 337900 245338 337912
rect 245390 337900 245396 337952
rect 245516 337949 245522 337952
rect 245473 337943 245522 337949
rect 245473 337909 245485 337943
rect 245519 337909 245522 337943
rect 245473 337903 245522 337909
rect 245516 337900 245522 337903
rect 245574 337900 245580 337952
rect 248276 337900 248282 337952
rect 248334 337949 248340 337952
rect 248334 337943 248383 337949
rect 248334 337909 248337 337943
rect 248371 337909 248383 337943
rect 248506 337940 248512 337952
rect 248467 337912 248512 337940
rect 248334 337903 248383 337909
rect 248334 337900 248340 337903
rect 248506 337900 248512 337912
rect 248564 337900 248570 337952
rect 249472 337940 249478 337952
rect 248616 337912 249478 337940
rect 234709 337875 234767 337881
rect 234709 337841 234721 337875
rect 234755 337872 234767 337875
rect 235488 337872 235494 337884
rect 234755 337844 235494 337872
rect 234755 337841 234767 337844
rect 234709 337835 234767 337841
rect 235488 337832 235494 337844
rect 235546 337832 235552 337884
rect 235856 337832 235862 337884
rect 235914 337881 235920 337884
rect 235914 337875 235963 337881
rect 235914 337841 235917 337875
rect 235951 337841 235963 337875
rect 235914 337835 235963 337841
rect 236917 337875 236975 337881
rect 236917 337841 236929 337875
rect 236963 337872 236975 337875
rect 237328 337872 237334 337884
rect 236963 337844 237334 337872
rect 236963 337841 236975 337844
rect 236917 337835 236975 337841
rect 235914 337832 235920 337835
rect 237328 337832 237334 337844
rect 237386 337832 237392 337884
rect 238064 337881 238070 337884
rect 238021 337875 238070 337881
rect 238021 337841 238033 337875
rect 238067 337841 238070 337875
rect 238021 337835 238070 337841
rect 238064 337832 238070 337835
rect 238122 337832 238128 337884
rect 238340 337832 238346 337884
rect 238398 337832 238404 337884
rect 238432 337832 238438 337884
rect 238490 337881 238496 337884
rect 238490 337875 238539 337881
rect 238490 337841 238493 337875
rect 238527 337841 238539 337875
rect 238490 337835 238539 337841
rect 238490 337832 238496 337835
rect 235672 337813 235678 337816
rect 235629 337807 235678 337813
rect 235629 337773 235641 337807
rect 235675 337773 235678 337807
rect 235629 337767 235678 337773
rect 235672 337764 235678 337767
rect 235730 337764 235736 337816
rect 236500 337813 236506 337816
rect 236457 337807 236506 337813
rect 236457 337773 236469 337807
rect 236503 337773 236506 337807
rect 236457 337767 236506 337773
rect 236500 337764 236506 337767
rect 236558 337764 236564 337816
rect 236592 337764 236598 337816
rect 236650 337813 236656 337816
rect 237512 337813 237518 337816
rect 236650 337807 236699 337813
rect 236650 337773 236653 337807
rect 236687 337773 236699 337807
rect 236650 337767 236699 337773
rect 237469 337807 237518 337813
rect 237469 337773 237481 337807
rect 237515 337773 237518 337807
rect 237469 337767 237518 337773
rect 236650 337764 236656 337767
rect 237512 337764 237518 337767
rect 237570 337764 237576 337816
rect 238358 337804 238386 337832
rect 239738 337816 239766 337900
rect 239904 337881 239910 337884
rect 239861 337875 239910 337881
rect 239861 337841 239873 337875
rect 239907 337841 239910 337875
rect 239861 337835 239910 337841
rect 239904 337832 239910 337835
rect 239962 337832 239968 337884
rect 240272 337832 240278 337884
rect 240330 337872 240336 337884
rect 240413 337875 240471 337881
rect 240413 337872 240425 337875
rect 240330 337844 240425 337872
rect 240330 337832 240336 337844
rect 240413 337841 240425 337844
rect 240459 337841 240471 337875
rect 240413 337835 240471 337841
rect 240548 337832 240554 337884
rect 240606 337872 240612 337884
rect 240689 337875 240747 337881
rect 240689 337872 240701 337875
rect 240606 337844 240701 337872
rect 240606 337832 240612 337844
rect 240689 337841 240701 337844
rect 240735 337841 240747 337875
rect 240689 337835 240747 337841
rect 241652 337832 241658 337884
rect 241710 337881 241716 337884
rect 241710 337875 241759 337881
rect 241710 337841 241713 337875
rect 241747 337841 241759 337875
rect 241710 337835 241759 337841
rect 241793 337875 241851 337881
rect 241793 337841 241805 337875
rect 241839 337872 241851 337875
rect 242296 337872 242302 337884
rect 241839 337844 242302 337872
rect 241839 337841 241851 337844
rect 241793 337835 241851 337841
rect 241710 337832 241716 337835
rect 242296 337832 242302 337844
rect 242354 337832 242360 337884
rect 242452 337816 242480 337900
rect 243032 337881 243038 337884
rect 242989 337875 243038 337881
rect 242989 337841 243001 337875
rect 243035 337841 243038 337875
rect 242989 337835 243038 337841
rect 243032 337832 243038 337835
rect 243090 337832 243096 337884
rect 243216 337832 243222 337884
rect 243274 337881 243280 337884
rect 243274 337875 243323 337881
rect 243274 337841 243277 337875
rect 243311 337841 243323 337875
rect 243274 337835 243323 337841
rect 243357 337875 243415 337881
rect 243357 337841 243369 337875
rect 243403 337872 243415 337875
rect 243584 337872 243590 337884
rect 243403 337844 243590 337872
rect 243403 337841 243415 337844
rect 243357 337835 243415 337841
rect 243274 337832 243280 337835
rect 243584 337832 243590 337844
rect 243642 337832 243648 337884
rect 243768 337832 243774 337884
rect 243826 337832 243832 337884
rect 244001 337875 244059 337881
rect 244001 337841 244013 337875
rect 244047 337872 244059 337875
rect 244228 337872 244234 337884
rect 244047 337844 244234 337872
rect 244047 337841 244059 337844
rect 244001 337835 244059 337841
rect 244228 337832 244234 337844
rect 244286 337832 244292 337884
rect 244369 337875 244427 337881
rect 244369 337841 244381 337875
rect 244415 337872 244427 337875
rect 244550 337872 244556 337884
rect 244415 337844 244556 337872
rect 244415 337841 244427 337844
rect 244369 337835 244427 337841
rect 244550 337832 244556 337844
rect 244608 337832 244614 337884
rect 245056 337832 245062 337884
rect 245114 337881 245120 337884
rect 245114 337875 245163 337881
rect 245114 337841 245117 337875
rect 245151 337841 245163 337875
rect 245114 337835 245163 337841
rect 245114 337832 245120 337835
rect 245884 337832 245890 337884
rect 245942 337832 245948 337884
rect 246117 337875 246175 337881
rect 246117 337841 246129 337875
rect 246163 337872 246175 337875
rect 246712 337872 246718 337884
rect 246163 337844 246718 337872
rect 246163 337841 246175 337844
rect 246117 337835 246175 337841
rect 246712 337832 246718 337844
rect 246770 337832 246776 337884
rect 246896 337881 246902 337884
rect 246853 337875 246902 337881
rect 246853 337841 246865 337875
rect 246899 337841 246902 337875
rect 246853 337835 246902 337841
rect 246896 337832 246902 337835
rect 246954 337832 246960 337884
rect 247037 337875 247095 337881
rect 247037 337841 247049 337875
rect 247083 337872 247095 337875
rect 247172 337872 247178 337884
rect 247083 337844 247178 337872
rect 247083 337841 247095 337844
rect 247037 337835 247095 337841
rect 247172 337832 247178 337844
rect 247230 337832 247236 337884
rect 247313 337875 247371 337881
rect 247313 337841 247325 337875
rect 247359 337872 247371 337875
rect 248092 337872 248098 337884
rect 247359 337844 248098 337872
rect 247359 337841 247371 337844
rect 247313 337835 247371 337841
rect 248092 337832 248098 337844
rect 248150 337832 248156 337884
rect 248417 337875 248475 337881
rect 248417 337841 248429 337875
rect 248463 337872 248475 337875
rect 248616 337872 248644 337912
rect 249472 337900 249478 337912
rect 249530 337900 249536 337952
rect 249840 337900 249846 337952
rect 249898 337900 249904 337952
rect 250533 337943 250591 337949
rect 250533 337909 250545 337943
rect 250579 337940 250591 337943
rect 250760 337940 250766 337952
rect 250579 337912 250766 337940
rect 250579 337909 250591 337912
rect 250533 337903 250591 337909
rect 250760 337900 250766 337912
rect 250818 337900 250824 337952
rect 250993 337943 251051 337949
rect 250993 337909 251005 337943
rect 251039 337940 251051 337943
rect 251128 337940 251134 337952
rect 251039 337912 251134 337940
rect 251039 337909 251051 337912
rect 250993 337903 251051 337909
rect 251128 337900 251134 337912
rect 251186 337900 251192 337952
rect 251220 337900 251226 337952
rect 251278 337900 251284 337952
rect 251404 337949 251410 337952
rect 251361 337943 251410 337949
rect 251361 337909 251373 337943
rect 251407 337909 251410 337943
rect 251361 337903 251410 337909
rect 251404 337900 251410 337903
rect 251462 337900 251468 337952
rect 251496 337900 251502 337952
rect 251554 337949 251560 337952
rect 251680 337949 251686 337952
rect 251554 337943 251603 337949
rect 251554 337909 251557 337943
rect 251591 337909 251603 337943
rect 251554 337903 251603 337909
rect 251637 337943 251686 337949
rect 251637 337909 251649 337943
rect 251683 337909 251686 337943
rect 251637 337903 251686 337909
rect 251554 337900 251560 337903
rect 251680 337900 251686 337903
rect 251738 337900 251744 337952
rect 252508 337949 252514 337952
rect 252465 337943 252514 337949
rect 252465 337909 252477 337943
rect 252511 337909 252514 337943
rect 252465 337903 252514 337909
rect 252508 337900 252514 337903
rect 252566 337900 252572 337952
rect 252649 337943 252707 337949
rect 252649 337909 252661 337943
rect 252695 337940 252707 337943
rect 253244 337940 253250 337952
rect 252695 337912 253250 337940
rect 252695 337909 252707 337912
rect 252649 337903 252707 337909
rect 253244 337900 253250 337912
rect 253302 337900 253308 337952
rect 253385 337943 253443 337949
rect 253385 337909 253397 337943
rect 253431 337940 253443 337943
rect 253520 337940 253526 337952
rect 253431 337912 253526 337940
rect 253431 337909 253443 337912
rect 253385 337903 253443 337909
rect 253520 337900 253526 337912
rect 253578 337900 253584 337952
rect 253796 337949 253802 337952
rect 253753 337943 253802 337949
rect 253753 337909 253765 337943
rect 253799 337909 253802 337943
rect 253753 337903 253802 337909
rect 253796 337900 253802 337903
rect 253854 337900 253860 337952
rect 254624 337900 254630 337952
rect 254682 337900 254688 337952
rect 254808 337900 254814 337952
rect 254866 337900 254872 337952
rect 255084 337940 255090 337952
rect 254918 337912 255090 337940
rect 248828 337881 248834 337884
rect 248463 337844 248644 337872
rect 248785 337875 248834 337881
rect 248463 337841 248475 337844
rect 248417 337835 248475 337841
rect 248785 337841 248797 337875
rect 248831 337841 248834 337875
rect 248785 337835 248834 337841
rect 248828 337832 248834 337835
rect 248886 337832 248892 337884
rect 248920 337832 248926 337884
rect 248978 337881 248984 337884
rect 248978 337875 249027 337881
rect 248978 337841 248981 337875
rect 249015 337841 249027 337875
rect 248978 337835 249027 337841
rect 249061 337875 249119 337881
rect 249061 337841 249073 337875
rect 249107 337872 249119 337875
rect 249288 337872 249294 337884
rect 249107 337844 249294 337872
rect 249107 337841 249119 337844
rect 249061 337835 249119 337841
rect 248978 337832 248984 337835
rect 249288 337832 249294 337844
rect 249346 337832 249352 337884
rect 249656 337881 249662 337884
rect 249613 337875 249662 337881
rect 249613 337841 249625 337875
rect 249659 337841 249662 337875
rect 249613 337835 249662 337841
rect 249656 337832 249662 337835
rect 249714 337832 249720 337884
rect 250116 337881 250122 337884
rect 250073 337875 250122 337881
rect 250073 337841 250085 337875
rect 250119 337841 250122 337875
rect 250073 337835 250122 337841
rect 250116 337832 250122 337835
rect 250174 337832 250180 337884
rect 238662 337804 238668 337816
rect 238358 337776 238668 337804
rect 238662 337764 238668 337776
rect 238720 337764 238726 337816
rect 238754 337764 238760 337816
rect 238812 337804 238818 337816
rect 239076 337804 239082 337816
rect 238812 337776 239082 337804
rect 238812 337764 238818 337776
rect 239076 337764 239082 337776
rect 239134 337764 239140 337816
rect 239738 337776 239772 337816
rect 239766 337764 239772 337776
rect 239824 337764 239830 337816
rect 242434 337764 242440 337816
rect 242492 337764 242498 337816
rect 242529 337807 242587 337813
rect 242529 337773 242541 337807
rect 242575 337804 242587 337807
rect 243786 337804 243814 337832
rect 244964 337813 244970 337816
rect 242575 337776 243814 337804
rect 244921 337807 244970 337813
rect 242575 337773 242587 337776
rect 242529 337767 242587 337773
rect 244921 337773 244933 337807
rect 244967 337773 244970 337807
rect 244921 337767 244970 337773
rect 244964 337764 244970 337767
rect 245022 337764 245028 337816
rect 245289 337807 245347 337813
rect 245289 337773 245301 337807
rect 245335 337804 245347 337807
rect 245424 337804 245430 337816
rect 245335 337776 245430 337804
rect 245335 337773 245347 337776
rect 245289 337767 245347 337773
rect 245424 337764 245430 337776
rect 245482 337764 245488 337816
rect 245749 337807 245807 337813
rect 245749 337773 245761 337807
rect 245795 337804 245807 337807
rect 245902 337804 245930 337832
rect 251238 337816 251266 337900
rect 252005 337875 252063 337881
rect 252005 337841 252017 337875
rect 252051 337872 252063 337875
rect 252784 337872 252790 337884
rect 252051 337844 252790 337872
rect 252051 337841 252063 337844
rect 252005 337835 252063 337841
rect 252784 337832 252790 337844
rect 252842 337832 252848 337884
rect 253109 337875 253167 337881
rect 253109 337841 253121 337875
rect 253155 337872 253167 337875
rect 253888 337872 253894 337884
rect 253155 337844 253894 337872
rect 253155 337841 253167 337844
rect 253109 337835 253167 337841
rect 253888 337832 253894 337844
rect 253946 337832 253952 337884
rect 254213 337875 254271 337881
rect 254213 337841 254225 337875
rect 254259 337872 254271 337875
rect 254440 337872 254446 337884
rect 254259 337844 254446 337872
rect 254259 337841 254271 337844
rect 254213 337835 254271 337841
rect 254440 337832 254446 337844
rect 254498 337832 254504 337884
rect 245795 337776 245930 337804
rect 249981 337807 250039 337813
rect 245795 337773 245807 337776
rect 245749 337767 245807 337773
rect 249981 337773 249993 337807
rect 250027 337804 250039 337807
rect 250668 337804 250674 337816
rect 250027 337776 250674 337804
rect 250027 337773 250039 337776
rect 249981 337767 250039 337773
rect 250668 337764 250674 337776
rect 250726 337764 250732 337816
rect 250809 337807 250867 337813
rect 250809 337773 250821 337807
rect 250855 337804 250867 337807
rect 250944 337804 250950 337816
rect 250855 337776 250950 337804
rect 250855 337773 250867 337776
rect 250809 337767 250867 337773
rect 250944 337764 250950 337776
rect 251002 337764 251008 337816
rect 251174 337764 251180 337816
rect 251232 337776 251266 337816
rect 251453 337807 251511 337813
rect 251232 337764 251238 337776
rect 251453 337773 251465 337807
rect 251499 337804 251511 337807
rect 251864 337804 251870 337816
rect 251499 337776 251870 337804
rect 251499 337773 251511 337776
rect 251453 337767 251511 337773
rect 251864 337764 251870 337776
rect 251922 337764 251928 337816
rect 253293 337807 253351 337813
rect 253293 337773 253305 337807
rect 253339 337804 253351 337807
rect 253428 337804 253434 337816
rect 253339 337776 253434 337804
rect 253339 337773 253351 337776
rect 253293 337767 253351 337773
rect 253428 337764 253434 337776
rect 253486 337764 253492 337816
rect 253569 337807 253627 337813
rect 253569 337773 253581 337807
rect 253615 337804 253627 337807
rect 253704 337804 253710 337816
rect 253615 337776 253710 337804
rect 253615 337773 253627 337776
rect 253569 337767 253627 337773
rect 253704 337764 253710 337776
rect 253762 337764 253768 337816
rect 254305 337807 254363 337813
rect 254305 337773 254317 337807
rect 254351 337804 254363 337807
rect 254918 337804 254946 337912
rect 255084 337900 255090 337912
rect 255142 337900 255148 337952
rect 255225 337943 255283 337949
rect 255225 337909 255237 337943
rect 255271 337940 255283 337943
rect 255360 337940 255366 337952
rect 255271 337912 255366 337940
rect 255271 337909 255283 337912
rect 255225 337903 255283 337909
rect 255360 337900 255366 337912
rect 255418 337900 255424 337952
rect 255636 337900 255642 337952
rect 255694 337940 255700 337952
rect 255777 337943 255835 337949
rect 255777 337940 255789 337943
rect 255694 337912 255789 337940
rect 255694 337900 255700 337912
rect 255777 337909 255789 337912
rect 255823 337909 255835 337943
rect 255777 337903 255835 337909
rect 255912 337900 255918 337952
rect 255970 337900 255976 337952
rect 256464 337900 256470 337952
rect 256522 337949 256528 337952
rect 256522 337943 256571 337949
rect 256522 337909 256525 337943
rect 256559 337909 256571 337943
rect 256522 337903 256571 337909
rect 256522 337900 256528 337903
rect 257108 337900 257114 337952
rect 257166 337949 257172 337952
rect 257166 337943 257215 337949
rect 257166 337909 257169 337943
rect 257203 337909 257215 337943
rect 257166 337903 257215 337909
rect 257166 337900 257172 337903
rect 257292 337900 257298 337952
rect 257350 337949 257356 337952
rect 257476 337949 257482 337952
rect 257350 337943 257399 337949
rect 257350 337909 257353 337943
rect 257387 337909 257399 337943
rect 257350 337903 257399 337909
rect 257433 337943 257482 337949
rect 257433 337909 257445 337943
rect 257479 337909 257482 337943
rect 257433 337903 257482 337909
rect 257350 337900 257356 337903
rect 257476 337900 257482 337903
rect 257534 337900 257540 337952
rect 257568 337900 257574 337952
rect 257626 337949 257632 337952
rect 257626 337943 257675 337949
rect 257626 337909 257629 337943
rect 257663 337909 257675 337943
rect 257626 337903 257675 337909
rect 257626 337900 257632 337903
rect 257844 337900 257850 337952
rect 257902 337940 257908 337952
rect 258672 337949 258678 337952
rect 257985 337943 258043 337949
rect 257985 337940 257997 337943
rect 257902 337912 257997 337940
rect 257902 337900 257908 337912
rect 257985 337909 257997 337912
rect 258031 337909 258043 337943
rect 257985 337903 258043 337909
rect 258629 337943 258678 337949
rect 258629 337909 258641 337943
rect 258675 337909 258678 337943
rect 258629 337903 258678 337909
rect 258672 337900 258678 337903
rect 258730 337900 258736 337952
rect 258856 337900 258862 337952
rect 258914 337949 258920 337952
rect 258914 337943 258963 337949
rect 258914 337909 258917 337943
rect 258951 337909 258963 337943
rect 258914 337903 258963 337909
rect 259089 337943 259147 337949
rect 259089 337909 259101 337943
rect 259135 337940 259147 337943
rect 259224 337940 259230 337952
rect 259135 337912 259230 337940
rect 259135 337909 259147 337912
rect 259089 337903 259147 337909
rect 258914 337900 258920 337903
rect 259224 337900 259230 337912
rect 259282 337900 259288 337952
rect 259408 337900 259414 337952
rect 259466 337949 259472 337952
rect 259466 337943 259515 337949
rect 259466 337909 259469 337943
rect 259503 337909 259515 337943
rect 259466 337903 259515 337909
rect 259466 337900 259472 337903
rect 259592 337900 259598 337952
rect 259650 337949 259656 337952
rect 259650 337943 259699 337949
rect 259650 337909 259653 337943
rect 259687 337909 259699 337943
rect 259650 337903 259699 337909
rect 259650 337900 259656 337903
rect 260052 337900 260058 337952
rect 260110 337940 260116 337952
rect 260193 337943 260251 337949
rect 260193 337940 260205 337943
rect 260110 337912 260205 337940
rect 260110 337900 260116 337912
rect 260193 337909 260205 337912
rect 260239 337909 260251 337943
rect 260193 337903 260251 337909
rect 260328 337900 260334 337952
rect 260386 337940 260392 337952
rect 260469 337943 260527 337949
rect 260469 337940 260481 337943
rect 260386 337912 260481 337940
rect 260386 337900 260392 337912
rect 260469 337909 260481 337912
rect 260515 337909 260527 337943
rect 260469 337903 260527 337909
rect 261248 337900 261254 337952
rect 261306 337940 261312 337952
rect 261757 337943 261815 337949
rect 261757 337940 261769 337943
rect 261306 337912 261769 337940
rect 261306 337900 261312 337912
rect 261757 337909 261769 337912
rect 261803 337909 261815 337943
rect 261757 337903 261815 337909
rect 262260 337900 262266 337952
rect 262318 337900 262324 337952
rect 262444 337949 262450 337952
rect 262401 337943 262450 337949
rect 262401 337909 262413 337943
rect 262447 337909 262450 337943
rect 262401 337903 262450 337909
rect 262444 337900 262450 337903
rect 262502 337900 262508 337952
rect 262536 337900 262542 337952
rect 262594 337940 262600 337952
rect 263229 337943 263287 337949
rect 263229 337940 263241 337943
rect 262594 337912 263241 337940
rect 262594 337900 262600 337912
rect 263229 337909 263241 337912
rect 263275 337909 263287 337943
rect 263229 337903 263287 337909
rect 264192 337900 264198 337952
rect 264250 337949 264256 337952
rect 264250 337943 264299 337949
rect 264250 337909 264253 337943
rect 264287 337909 264299 337943
rect 264250 337903 264299 337909
rect 264609 337943 264667 337949
rect 264609 337909 264621 337943
rect 264655 337940 264667 337943
rect 264744 337940 264750 337952
rect 264655 337912 264750 337940
rect 264655 337909 264667 337912
rect 264609 337903 264667 337909
rect 264250 337900 264256 337903
rect 264744 337900 264750 337912
rect 264802 337900 264808 337952
rect 264928 337900 264934 337952
rect 264986 337900 264992 337952
rect 265020 337900 265026 337952
rect 265078 337949 265084 337952
rect 265078 337943 265127 337949
rect 265078 337909 265081 337943
rect 265115 337909 265127 337943
rect 265078 337903 265127 337909
rect 265078 337900 265084 337903
rect 265204 337900 265210 337952
rect 265262 337949 265268 337952
rect 265262 337943 265311 337949
rect 265262 337909 265265 337943
rect 265299 337909 265311 337943
rect 265262 337903 265311 337909
rect 265262 337900 265268 337903
rect 265388 337900 265394 337952
rect 265446 337949 265452 337952
rect 265446 337943 265495 337949
rect 265446 337909 265449 337943
rect 265483 337909 265495 337943
rect 265446 337903 265495 337909
rect 265446 337900 265452 337903
rect 266492 337900 266498 337952
rect 266550 337949 266556 337952
rect 266676 337949 266682 337952
rect 266550 337943 266599 337949
rect 266550 337909 266553 337943
rect 266587 337909 266599 337943
rect 266550 337903 266599 337909
rect 266633 337943 266682 337949
rect 266633 337909 266645 337943
rect 266679 337909 266682 337943
rect 266633 337903 266682 337909
rect 266550 337900 266556 337903
rect 266676 337900 266682 337903
rect 266734 337900 266740 337952
rect 266768 337900 266774 337952
rect 266826 337949 266832 337952
rect 266826 337943 266875 337949
rect 266826 337909 266829 337943
rect 266863 337909 266875 337943
rect 266826 337903 266875 337909
rect 266826 337900 266832 337903
rect 267320 337900 267326 337952
rect 267378 337949 267384 337952
rect 267378 337943 267427 337949
rect 267378 337909 267381 337943
rect 267415 337909 267427 337943
rect 267378 337903 267427 337909
rect 267378 337900 267384 337903
rect 268332 337900 268338 337952
rect 268390 337949 268396 337952
rect 268390 337943 268439 337949
rect 268390 337909 268393 337943
rect 268427 337909 268439 337943
rect 268390 337903 268439 337909
rect 268390 337900 268396 337903
rect 268608 337900 268614 337952
rect 268666 337940 268672 337952
rect 268666 337900 268700 337940
rect 269068 337900 269074 337952
rect 269126 337940 269132 337952
rect 269209 337943 269267 337949
rect 269209 337940 269221 337943
rect 269126 337912 269221 337940
rect 269126 337900 269132 337912
rect 269209 337909 269221 337912
rect 269255 337909 269267 337943
rect 269209 337903 269267 337909
rect 269344 337900 269350 337952
rect 269402 337940 269408 337952
rect 270448 337949 270454 337952
rect 270037 337943 270095 337949
rect 270037 337940 270049 337943
rect 269402 337912 270049 337940
rect 269402 337900 269408 337912
rect 270037 337909 270049 337912
rect 270083 337909 270095 337943
rect 270037 337903 270095 337909
rect 270405 337943 270454 337949
rect 270405 337909 270417 337943
rect 270451 337909 270454 337943
rect 270405 337903 270454 337909
rect 270448 337900 270454 337903
rect 270506 337900 270512 337952
rect 270540 337900 270546 337952
rect 270598 337940 270604 337952
rect 271969 337943 272027 337949
rect 271969 337940 271981 337943
rect 270598 337912 271981 337940
rect 270598 337900 270604 337912
rect 271969 337909 271981 337912
rect 272015 337909 272027 337943
rect 271969 337903 272027 337909
rect 272061 337943 272119 337949
rect 272061 337909 272073 337943
rect 272107 337940 272119 337943
rect 272196 337940 272202 337952
rect 272107 337912 272202 337940
rect 272107 337909 272119 337912
rect 272061 337903 272119 337909
rect 272196 337900 272202 337912
rect 272254 337900 272260 337952
rect 272380 337900 272386 337952
rect 272438 337900 272444 337952
rect 272748 337900 272754 337952
rect 272806 337940 272812 337952
rect 272981 337943 273039 337949
rect 272981 337940 272993 337943
rect 272806 337912 272993 337940
rect 272806 337900 272812 337912
rect 272981 337909 272993 337912
rect 273027 337909 273039 337943
rect 272981 337903 273039 337909
rect 274220 337900 274226 337952
rect 274278 337940 274284 337952
rect 274453 337943 274511 337949
rect 274453 337940 274465 337943
rect 274278 337912 274465 337940
rect 274278 337900 274284 337912
rect 274453 337909 274465 337912
rect 274499 337909 274511 337943
rect 274453 337903 274511 337909
rect 274864 337900 274870 337952
rect 274922 337949 274928 337952
rect 274922 337943 274971 337949
rect 274922 337909 274925 337943
rect 274959 337909 274971 337943
rect 274922 337903 274971 337909
rect 274922 337900 274928 337903
rect 275140 337900 275146 337952
rect 275198 337940 275204 337952
rect 275465 337943 275523 337949
rect 275465 337940 275477 337943
rect 275198 337912 275477 337940
rect 275198 337900 275204 337912
rect 275465 337909 275477 337912
rect 275511 337909 275523 337943
rect 275465 337903 275523 337909
rect 275968 337900 275974 337952
rect 276026 337900 276032 337952
rect 276152 337900 276158 337952
rect 276210 337900 276216 337952
rect 276428 337900 276434 337952
rect 276486 337940 276492 337952
rect 276753 337943 276811 337949
rect 276753 337940 276765 337943
rect 276486 337912 276765 337940
rect 276486 337900 276492 337912
rect 276753 337909 276765 337912
rect 276799 337909 276811 337943
rect 276753 337903 276811 337909
rect 277072 337900 277078 337952
rect 277130 337940 277136 337952
rect 277581 337943 277639 337949
rect 277581 337940 277593 337943
rect 277130 337912 277593 337940
rect 277130 337900 277136 337912
rect 277581 337909 277593 337912
rect 277627 337909 277639 337943
rect 277581 337903 277639 337909
rect 278084 337900 278090 337952
rect 278142 337949 278148 337952
rect 278360 337949 278366 337952
rect 278142 337943 278191 337949
rect 278142 337909 278145 337943
rect 278179 337909 278191 337943
rect 278142 337903 278191 337909
rect 278317 337943 278366 337949
rect 278317 337909 278329 337943
rect 278363 337909 278366 337943
rect 278317 337903 278366 337909
rect 278142 337900 278148 337903
rect 278360 337900 278366 337903
rect 278418 337900 278424 337952
rect 278728 337900 278734 337952
rect 278786 337940 278792 337952
rect 278930 337940 278958 337980
rect 279237 337977 279249 337980
rect 279283 337977 279295 338011
rect 279237 337971 279295 337977
rect 282518 337952 282546 338116
rect 282917 338113 282929 338116
rect 282963 338113 282975 338147
rect 282917 338107 282975 338113
rect 287422 338104 287428 338156
rect 287480 338144 287486 338156
rect 296530 338144 296536 338156
rect 287480 338116 296536 338144
rect 287480 338104 287486 338116
rect 296530 338104 296536 338116
rect 296588 338104 296594 338156
rect 287701 338079 287759 338085
rect 287701 338076 287713 338079
rect 282610 338048 287713 338076
rect 278786 337912 278958 337940
rect 278786 337900 278792 337912
rect 279096 337900 279102 337952
rect 279154 337940 279160 337952
rect 281169 337943 281227 337949
rect 281169 337940 281181 337943
rect 279154 337912 281181 337940
rect 279154 337900 279160 337912
rect 281169 337909 281181 337912
rect 281215 337909 281227 337943
rect 281169 337903 281227 337909
rect 281304 337900 281310 337952
rect 281362 337949 281368 337952
rect 281362 337943 281411 337949
rect 281362 337909 281365 337943
rect 281399 337909 281411 337943
rect 281362 337903 281411 337909
rect 281362 337900 281368 337903
rect 281672 337900 281678 337952
rect 281730 337949 281736 337952
rect 281730 337943 281779 337949
rect 281730 337909 281733 337943
rect 281767 337909 281779 337943
rect 281730 337903 281779 337909
rect 281730 337900 281736 337903
rect 281856 337900 281862 337952
rect 281914 337940 281920 337952
rect 281997 337943 282055 337949
rect 281997 337940 282009 337943
rect 281914 337912 282009 337940
rect 281914 337900 281920 337912
rect 281997 337909 282009 337912
rect 282043 337909 282055 337943
rect 281997 337903 282055 337909
rect 282132 337900 282138 337952
rect 282190 337949 282196 337952
rect 282190 337943 282239 337949
rect 282190 337909 282193 337943
rect 282227 337909 282239 337943
rect 282190 337903 282239 337909
rect 282273 337943 282331 337949
rect 282273 337909 282285 337943
rect 282319 337940 282331 337943
rect 282408 337940 282414 337952
rect 282319 337912 282414 337940
rect 282319 337909 282331 337912
rect 282273 337903 282331 337909
rect 282190 337900 282196 337903
rect 282408 337900 282414 337912
rect 282466 337900 282472 337952
rect 282500 337900 282506 337952
rect 282558 337900 282564 337952
rect 254992 337832 254998 337884
rect 255050 337832 255056 337884
rect 255544 337872 255550 337884
rect 255424 337844 255550 337872
rect 254351 337776 254946 337804
rect 255010 337804 255038 337832
rect 255424 337816 255452 337844
rect 255544 337832 255550 337844
rect 255602 337832 255608 337884
rect 255930 337816 255958 337900
rect 256280 337832 256286 337884
rect 256338 337881 256344 337884
rect 256338 337875 256387 337881
rect 256338 337841 256341 337875
rect 256375 337841 256387 337875
rect 256338 337835 256387 337841
rect 256338 337832 256344 337835
rect 256648 337832 256654 337884
rect 256706 337872 256712 337884
rect 256881 337875 256939 337881
rect 256881 337872 256893 337875
rect 256706 337844 256893 337872
rect 256706 337832 256712 337844
rect 256881 337841 256893 337844
rect 256927 337841 256939 337875
rect 256881 337835 256939 337841
rect 257016 337832 257022 337884
rect 257074 337872 257080 337884
rect 258077 337875 258135 337881
rect 258077 337872 258089 337875
rect 257074 337844 258089 337872
rect 257074 337832 257080 337844
rect 258077 337841 258089 337844
rect 258123 337841 258135 337875
rect 258077 337835 258135 337841
rect 258488 337832 258494 337884
rect 258546 337881 258552 337884
rect 258546 337875 258595 337881
rect 258546 337841 258549 337875
rect 258583 337841 258595 337875
rect 258546 337835 258595 337841
rect 258546 337832 258552 337835
rect 258764 337832 258770 337884
rect 258822 337872 258828 337884
rect 260604 337881 260610 337884
rect 259825 337875 259883 337881
rect 259825 337872 259837 337875
rect 258822 337844 259837 337872
rect 258822 337832 258828 337844
rect 259825 337841 259837 337844
rect 259871 337841 259883 337875
rect 259825 337835 259883 337841
rect 260561 337875 260610 337881
rect 260561 337841 260573 337875
rect 260607 337841 260610 337875
rect 260561 337835 260610 337841
rect 260604 337832 260610 337835
rect 260662 337832 260668 337884
rect 261156 337881 261162 337884
rect 261113 337875 261162 337881
rect 261113 337841 261125 337875
rect 261159 337841 261162 337875
rect 261113 337835 261162 337841
rect 261156 337832 261162 337835
rect 261214 337832 261220 337884
rect 261432 337832 261438 337884
rect 261490 337872 261496 337884
rect 262168 337881 262174 337884
rect 262033 337875 262091 337881
rect 262033 337872 262045 337875
rect 261490 337844 262045 337872
rect 261490 337832 261496 337844
rect 262033 337841 262045 337844
rect 262079 337841 262091 337875
rect 262033 337835 262091 337841
rect 262125 337875 262174 337881
rect 262125 337841 262137 337875
rect 262171 337841 262174 337875
rect 262125 337835 262174 337841
rect 262168 337832 262174 337835
rect 262226 337832 262232 337884
rect 262628 337832 262634 337884
rect 262686 337881 262692 337884
rect 262686 337875 262735 337881
rect 262686 337841 262689 337875
rect 262723 337841 262735 337875
rect 262686 337835 262735 337841
rect 262686 337832 262692 337835
rect 262812 337832 262818 337884
rect 262870 337881 262876 337884
rect 262870 337875 262919 337881
rect 262870 337841 262873 337875
rect 262907 337841 262919 337875
rect 262870 337835 262919 337841
rect 262953 337875 263011 337881
rect 262953 337841 262965 337875
rect 262999 337872 263011 337875
rect 263088 337872 263094 337884
rect 262999 337844 263094 337872
rect 262999 337841 263011 337844
rect 262953 337835 263011 337841
rect 262870 337832 262876 337835
rect 263088 337832 263094 337844
rect 263146 337832 263152 337884
rect 263640 337832 263646 337884
rect 263698 337881 263704 337884
rect 263698 337875 263747 337881
rect 263698 337841 263701 337875
rect 263735 337841 263747 337875
rect 263698 337835 263747 337841
rect 263698 337832 263704 337835
rect 264376 337832 264382 337884
rect 264434 337872 264440 337884
rect 264517 337875 264575 337881
rect 264517 337872 264529 337875
rect 264434 337844 264529 337872
rect 264434 337832 264440 337844
rect 264517 337841 264529 337844
rect 264563 337841 264575 337875
rect 264946 337872 264974 337900
rect 266952 337881 266958 337884
rect 266357 337875 266415 337881
rect 266357 337872 266369 337875
rect 264946 337844 266369 337872
rect 264517 337835 264575 337841
rect 266357 337841 266369 337844
rect 266403 337841 266415 337875
rect 266357 337835 266415 337841
rect 266909 337875 266958 337881
rect 266909 337841 266921 337875
rect 266955 337841 266958 337875
rect 266909 337835 266958 337841
rect 266952 337832 266958 337835
rect 267010 337832 267016 337884
rect 267228 337832 267234 337884
rect 267286 337872 267292 337884
rect 267737 337875 267795 337881
rect 267737 337872 267749 337875
rect 267286 337844 267749 337872
rect 267286 337832 267292 337844
rect 267737 337841 267749 337844
rect 267783 337841 267795 337875
rect 267737 337835 267795 337841
rect 267872 337832 267878 337884
rect 267930 337872 267936 337884
rect 268148 337881 268154 337884
rect 268013 337875 268071 337881
rect 268013 337872 268025 337875
rect 267930 337844 268025 337872
rect 267930 337832 267936 337844
rect 268013 337841 268025 337844
rect 268059 337841 268071 337875
rect 268013 337835 268071 337841
rect 268105 337875 268154 337881
rect 268105 337841 268117 337875
rect 268151 337841 268154 337875
rect 268105 337835 268154 337841
rect 268148 337832 268154 337835
rect 268206 337832 268212 337884
rect 255133 337807 255191 337813
rect 255133 337804 255145 337807
rect 255010 337776 255145 337804
rect 254351 337773 254363 337776
rect 254305 337767 254363 337773
rect 255133 337773 255145 337776
rect 255179 337773 255191 337807
rect 255133 337767 255191 337773
rect 255406 337764 255412 337816
rect 255464 337764 255470 337816
rect 255930 337776 255964 337816
rect 255958 337764 255964 337776
rect 256016 337764 256022 337816
rect 257200 337764 257206 337816
rect 257258 337804 257264 337816
rect 257893 337807 257951 337813
rect 257893 337804 257905 337807
rect 257258 337776 257905 337804
rect 257258 337764 257264 337776
rect 257893 337773 257905 337776
rect 257939 337773 257951 337807
rect 257893 337767 257951 337773
rect 258304 337764 258310 337816
rect 258362 337813 258368 337816
rect 258362 337807 258411 337813
rect 258362 337773 258365 337807
rect 258399 337773 258411 337807
rect 258362 337767 258411 337773
rect 258362 337764 258368 337767
rect 260880 337764 260886 337816
rect 260938 337804 260944 337816
rect 265713 337807 265771 337813
rect 265713 337804 265725 337807
rect 260938 337776 265725 337804
rect 260938 337764 260944 337776
rect 265713 337773 265725 337776
rect 265759 337773 265771 337807
rect 265713 337767 265771 337773
rect 268424 337764 268430 337816
rect 268482 337813 268488 337816
rect 268482 337807 268531 337813
rect 268482 337773 268485 337807
rect 268519 337773 268531 337807
rect 268672 337804 268700 337900
rect 268792 337832 268798 337884
rect 268850 337881 268856 337884
rect 268976 337881 268982 337884
rect 268850 337875 268899 337881
rect 268850 337841 268853 337875
rect 268887 337841 268899 337875
rect 268850 337835 268899 337841
rect 268933 337875 268982 337881
rect 268933 337841 268945 337875
rect 268979 337841 268982 337875
rect 268933 337835 268982 337841
rect 268850 337832 268856 337835
rect 268976 337832 268982 337835
rect 269034 337832 269040 337884
rect 269761 337875 269819 337881
rect 269761 337841 269773 337875
rect 269807 337872 269819 337875
rect 269896 337872 269902 337884
rect 269807 337844 269902 337872
rect 269807 337841 269819 337844
rect 269761 337835 269819 337841
rect 269896 337832 269902 337844
rect 269954 337832 269960 337884
rect 270172 337832 270178 337884
rect 270230 337872 270236 337884
rect 270313 337875 270371 337881
rect 270313 337872 270325 337875
rect 270230 337844 270325 337872
rect 270230 337832 270236 337844
rect 270313 337841 270325 337844
rect 270359 337841 270371 337875
rect 270313 337835 270371 337841
rect 271000 337832 271006 337884
rect 271058 337881 271064 337884
rect 271368 337881 271374 337884
rect 271058 337875 271107 337881
rect 271058 337841 271061 337875
rect 271095 337841 271107 337875
rect 271058 337835 271107 337841
rect 271325 337875 271374 337881
rect 271325 337841 271337 337875
rect 271371 337841 271374 337875
rect 271325 337835 271374 337841
rect 271058 337832 271064 337835
rect 271368 337832 271374 337835
rect 271426 337832 271432 337884
rect 271506 337832 271512 337884
rect 271564 337872 271570 337884
rect 271564 337844 271609 337872
rect 271564 337832 271570 337844
rect 271644 337832 271650 337884
rect 271702 337872 271708 337884
rect 271785 337875 271843 337881
rect 271785 337872 271797 337875
rect 271702 337844 271797 337872
rect 271702 337832 271708 337844
rect 271785 337841 271797 337844
rect 271831 337841 271843 337875
rect 271785 337835 271843 337841
rect 271877 337875 271935 337881
rect 271877 337841 271889 337875
rect 271923 337872 271935 337875
rect 272840 337872 272846 337884
rect 271923 337844 272846 337872
rect 271923 337841 271935 337844
rect 271877 337835 271935 337841
rect 272840 337832 272846 337844
rect 272898 337832 272904 337884
rect 273760 337832 273766 337884
rect 273818 337881 273824 337884
rect 273944 337881 273950 337884
rect 273818 337875 273867 337881
rect 273818 337841 273821 337875
rect 273855 337841 273867 337875
rect 273818 337835 273867 337841
rect 273901 337875 273950 337881
rect 273901 337841 273913 337875
rect 273947 337841 273950 337875
rect 273901 337835 273950 337841
rect 273818 337832 273824 337835
rect 273944 337832 273950 337835
rect 274002 337832 274008 337884
rect 274128 337832 274134 337884
rect 274186 337872 274192 337884
rect 274361 337875 274419 337881
rect 274361 337872 274373 337875
rect 274186 337844 274373 337872
rect 274186 337832 274192 337844
rect 274361 337841 274373 337844
rect 274407 337841 274419 337875
rect 274361 337835 274419 337841
rect 275649 337875 275707 337881
rect 275649 337841 275661 337875
rect 275695 337872 275707 337875
rect 275784 337872 275790 337884
rect 275695 337844 275790 337872
rect 275695 337841 275707 337844
rect 275649 337835 275707 337841
rect 275784 337832 275790 337844
rect 275842 337832 275848 337884
rect 276336 337832 276342 337884
rect 276394 337872 276400 337884
rect 276569 337875 276627 337881
rect 276569 337872 276581 337875
rect 276394 337844 276581 337872
rect 276394 337832 276400 337844
rect 276569 337841 276581 337844
rect 276615 337841 276627 337875
rect 276569 337835 276627 337841
rect 277716 337832 277722 337884
rect 277774 337872 277780 337884
rect 277857 337875 277915 337881
rect 277857 337872 277869 337875
rect 277774 337844 277869 337872
rect 277774 337832 277780 337844
rect 277857 337841 277869 337844
rect 277903 337841 277915 337875
rect 277857 337835 277915 337841
rect 277992 337832 277998 337884
rect 278050 337872 278056 337884
rect 278225 337875 278283 337881
rect 278225 337872 278237 337875
rect 278050 337844 278237 337872
rect 278050 337832 278056 337844
rect 278225 337841 278237 337844
rect 278271 337841 278283 337875
rect 278225 337835 278283 337841
rect 279556 337832 279562 337884
rect 279614 337872 279620 337884
rect 279697 337875 279755 337881
rect 279697 337872 279709 337875
rect 279614 337844 279709 337872
rect 279614 337832 279620 337844
rect 279697 337841 279709 337844
rect 279743 337841 279755 337875
rect 279697 337835 279755 337841
rect 279789 337875 279847 337881
rect 279789 337841 279801 337875
rect 279835 337872 279847 337875
rect 280108 337872 280114 337884
rect 279835 337844 280114 337872
rect 279835 337841 279847 337844
rect 279789 337835 279847 337841
rect 280108 337832 280114 337844
rect 280166 337832 280172 337884
rect 280200 337832 280206 337884
rect 280258 337872 280264 337884
rect 280433 337875 280491 337881
rect 280433 337872 280445 337875
rect 280258 337844 280445 337872
rect 280258 337832 280264 337844
rect 280433 337841 280445 337844
rect 280479 337841 280491 337875
rect 280433 337835 280491 337841
rect 280568 337832 280574 337884
rect 280626 337872 280632 337884
rect 280709 337875 280767 337881
rect 280709 337872 280721 337875
rect 280626 337844 280721 337872
rect 280626 337832 280632 337844
rect 280709 337841 280721 337844
rect 280755 337841 280767 337875
rect 280709 337835 280767 337841
rect 280844 337832 280850 337884
rect 280902 337872 280908 337884
rect 282610 337872 282638 338048
rect 287701 338045 287713 338048
rect 287747 338045 287759 338079
rect 287701 338039 287759 338045
rect 285214 338008 285220 338020
rect 283898 337980 285220 338008
rect 283898 337952 283926 337980
rect 285214 337968 285220 337980
rect 285272 337968 285278 338020
rect 283880 337900 283886 337952
rect 283938 337900 283944 337952
rect 284064 337900 284070 337952
rect 284122 337940 284128 337952
rect 288250 337940 288256 337952
rect 284122 337912 288256 337940
rect 284122 337900 284128 337912
rect 288250 337900 288256 337912
rect 288308 337900 288314 337952
rect 280902 337844 282638 337872
rect 280902 337832 280908 337844
rect 284248 337832 284254 337884
rect 284306 337872 284312 337884
rect 284389 337875 284447 337881
rect 284389 337872 284401 337875
rect 284306 337844 284401 337872
rect 284306 337832 284312 337844
rect 284389 337841 284401 337844
rect 284435 337841 284447 337875
rect 284389 337835 284447 337841
rect 278777 337807 278835 337813
rect 278777 337804 278789 337807
rect 268672 337776 278789 337804
rect 268482 337767 268531 337773
rect 278777 337773 278789 337776
rect 278823 337773 278835 337807
rect 278777 337767 278835 337773
rect 268482 337764 268488 337767
rect 278912 337764 278918 337816
rect 278970 337804 278976 337816
rect 288069 337807 288127 337813
rect 288069 337804 288081 337807
rect 278970 337776 288081 337804
rect 278970 337764 278976 337776
rect 288069 337773 288081 337776
rect 288115 337773 288127 337807
rect 288069 337767 288127 337773
rect 436738 337736 436744 337748
rect 234586 337708 436744 337736
rect 436738 337696 436744 337708
rect 436796 337696 436802 337748
rect 479518 337668 479524 337680
rect 234586 337640 479524 337668
rect 232314 337492 232320 337544
rect 232372 337532 232378 337544
rect 234586 337532 234614 337640
rect 479518 337628 479524 337640
rect 479576 337628 479582 337680
rect 235442 337600 235448 337612
rect 235403 337572 235448 337600
rect 235442 337560 235448 337572
rect 235500 337560 235506 337612
rect 235626 337600 235632 337612
rect 235587 337572 235632 337600
rect 235626 337560 235632 337572
rect 235684 337560 235690 337612
rect 237745 337603 237803 337609
rect 237745 337569 237757 337603
rect 237791 337600 237803 337603
rect 237834 337600 237840 337612
rect 237791 337572 237840 337600
rect 237791 337569 237803 337572
rect 237745 337563 237803 337569
rect 237834 337560 237840 337572
rect 237892 337560 237898 337612
rect 238018 337600 238024 337612
rect 237979 337572 238024 337600
rect 238018 337560 238024 337572
rect 238076 337560 238082 337612
rect 238481 337603 238539 337609
rect 238481 337569 238493 337603
rect 238527 337600 238539 337603
rect 238570 337600 238576 337612
rect 238527 337572 238576 337600
rect 238527 337569 238539 337572
rect 238481 337563 238539 337569
rect 238570 337560 238576 337572
rect 238628 337560 238634 337612
rect 239217 337603 239275 337609
rect 239217 337569 239229 337603
rect 239263 337600 239275 337603
rect 239306 337600 239312 337612
rect 239263 337572 239312 337600
rect 239263 337569 239275 337572
rect 239217 337563 239275 337569
rect 239306 337560 239312 337572
rect 239364 337560 239370 337612
rect 239401 337603 239459 337609
rect 239401 337569 239413 337603
rect 239447 337600 239459 337603
rect 483014 337600 483020 337612
rect 239447 337572 483020 337600
rect 239447 337569 239459 337572
rect 239401 337563 239459 337569
rect 483014 337560 483020 337572
rect 483072 337560 483078 337612
rect 232372 337504 234614 337532
rect 232372 337492 232378 337504
rect 234982 337492 234988 337544
rect 235040 337532 235046 337544
rect 237469 337535 237527 337541
rect 237469 337532 237481 337535
rect 235040 337504 237481 337532
rect 235040 337492 235046 337504
rect 237469 337501 237481 337504
rect 237515 337501 237527 337535
rect 237469 337495 237527 337501
rect 240689 337535 240747 337541
rect 240689 337501 240701 337535
rect 240735 337532 240747 337535
rect 241146 337532 241152 337544
rect 240735 337504 241152 337532
rect 240735 337501 240747 337504
rect 240689 337495 240747 337501
rect 241146 337492 241152 337504
rect 241204 337492 241210 337544
rect 243354 337532 243360 337544
rect 243315 337504 243360 337532
rect 243354 337492 243360 337504
rect 243412 337492 243418 337544
rect 243998 337532 244004 337544
rect 243959 337504 244004 337532
rect 243998 337492 244004 337504
rect 244056 337492 244062 337544
rect 246114 337532 246120 337544
rect 246075 337504 246120 337532
rect 246114 337492 246120 337504
rect 246172 337492 246178 337544
rect 246850 337532 246856 337544
rect 246811 337504 246856 337532
rect 246850 337492 246856 337504
rect 246908 337492 246914 337544
rect 247034 337532 247040 337544
rect 246995 337504 247040 337532
rect 247034 337492 247040 337504
rect 247092 337492 247098 337544
rect 249058 337532 249064 337544
rect 249019 337504 249064 337532
rect 249058 337492 249064 337504
rect 249116 337492 249122 337544
rect 253106 337532 253112 337544
rect 253067 337504 253112 337532
rect 253106 337492 253112 337504
rect 253164 337492 253170 337544
rect 253290 337532 253296 337544
rect 253251 337504 253296 337532
rect 253290 337492 253296 337504
rect 253348 337492 253354 337544
rect 253750 337532 253756 337544
rect 253711 337504 253756 337532
rect 253750 337492 253756 337504
rect 253808 337492 253814 337544
rect 254029 337535 254087 337541
rect 254029 337501 254041 337535
rect 254075 337532 254087 337535
rect 254854 337532 254860 337544
rect 254075 337504 254860 337532
rect 254075 337501 254087 337504
rect 254029 337495 254087 337501
rect 254854 337492 254860 337504
rect 254912 337492 254918 337544
rect 256329 337535 256387 337541
rect 256329 337501 256341 337535
rect 256375 337532 256387 337535
rect 256418 337532 256424 337544
rect 256375 337504 256424 337532
rect 256375 337501 256387 337504
rect 256329 337495 256387 337501
rect 256418 337492 256424 337504
rect 256476 337492 256482 337544
rect 257157 337535 257215 337541
rect 257157 337501 257169 337535
rect 257203 337532 257215 337535
rect 257706 337532 257712 337544
rect 257203 337504 257712 337532
rect 257203 337501 257215 337504
rect 257157 337495 257215 337501
rect 257706 337492 257712 337504
rect 257764 337492 257770 337544
rect 258626 337492 258632 337544
rect 258684 337532 258690 337544
rect 259089 337535 259147 337541
rect 259089 337532 259101 337535
rect 258684 337504 259101 337532
rect 258684 337492 258690 337504
rect 259089 337501 259101 337504
rect 259135 337501 259147 337535
rect 259089 337495 259147 337501
rect 260193 337535 260251 337541
rect 260193 337501 260205 337535
rect 260239 337532 260251 337535
rect 260558 337532 260564 337544
rect 260239 337504 260564 337532
rect 260239 337501 260251 337504
rect 260193 337495 260251 337501
rect 260558 337492 260564 337504
rect 260616 337492 260622 337544
rect 262401 337535 262459 337541
rect 262401 337501 262413 337535
rect 262447 337532 262459 337535
rect 262766 337532 262772 337544
rect 262447 337504 262772 337532
rect 262447 337501 262459 337504
rect 262401 337495 262459 337501
rect 262766 337492 262772 337504
rect 262824 337492 262830 337544
rect 262950 337532 262956 337544
rect 262911 337504 262956 337532
rect 262950 337492 262956 337504
rect 263008 337492 263014 337544
rect 265434 337532 265440 337544
rect 265395 337504 265440 337532
rect 265434 337492 265440 337504
rect 265492 337492 265498 337544
rect 268010 337532 268016 337544
rect 267971 337504 268016 337532
rect 268010 337492 268016 337504
rect 268068 337492 268074 337544
rect 268841 337535 268899 337541
rect 268841 337501 268853 337535
rect 268887 337532 268899 337535
rect 269577 337535 269635 337541
rect 269577 337532 269589 337535
rect 268887 337504 269589 337532
rect 268887 337501 268899 337504
rect 268841 337495 268899 337501
rect 269577 337501 269589 337504
rect 269623 337501 269635 337535
rect 269758 337532 269764 337544
rect 269719 337504 269764 337532
rect 269577 337495 269635 337501
rect 269758 337492 269764 337504
rect 269816 337492 269822 337544
rect 270310 337532 270316 337544
rect 270271 337504 270316 337532
rect 270310 337492 270316 337504
rect 270368 337492 270374 337544
rect 271322 337532 271328 337544
rect 271283 337504 271328 337532
rect 271322 337492 271328 337504
rect 271380 337492 271386 337544
rect 271874 337532 271880 337544
rect 271835 337504 271880 337532
rect 271874 337492 271880 337504
rect 271932 337492 271938 337544
rect 272981 337535 273039 337541
rect 272981 337501 272993 337535
rect 273027 337532 273039 337535
rect 275278 337532 275284 337544
rect 273027 337504 275284 337532
rect 273027 337501 273039 337504
rect 272981 337495 273039 337501
rect 275278 337492 275284 337504
rect 275336 337492 275342 337544
rect 275649 337535 275707 337541
rect 275649 337501 275661 337535
rect 275695 337532 275707 337535
rect 275738 337532 275744 337544
rect 275695 337504 275744 337532
rect 275695 337501 275707 337504
rect 275649 337495 275707 337501
rect 275738 337492 275744 337504
rect 275796 337492 275802 337544
rect 276382 337492 276388 337544
rect 276440 337532 276446 337544
rect 276569 337535 276627 337541
rect 276569 337532 276581 337535
rect 276440 337504 276581 337532
rect 276440 337492 276446 337504
rect 276569 337501 276581 337504
rect 276615 337501 276627 337535
rect 276569 337495 276627 337501
rect 276937 337535 276995 337541
rect 276937 337501 276949 337535
rect 276983 337532 276995 337535
rect 277118 337532 277124 337544
rect 276983 337504 277124 337532
rect 276983 337501 276995 337504
rect 276937 337495 276995 337501
rect 277118 337492 277124 337504
rect 277176 337492 277182 337544
rect 278314 337532 278320 337544
rect 278275 337504 278320 337532
rect 278314 337492 278320 337504
rect 278372 337492 278378 337544
rect 282273 337535 282331 337541
rect 282273 337501 282285 337535
rect 282319 337532 282331 337535
rect 282362 337532 282368 337544
rect 282319 337504 282368 337532
rect 282319 337501 282331 337504
rect 282273 337495 282331 337501
rect 282362 337492 282368 337504
rect 282420 337492 282426 337544
rect 282549 337535 282607 337541
rect 282549 337501 282561 337535
rect 282595 337532 282607 337535
rect 282914 337532 282920 337544
rect 282595 337504 282920 337532
rect 282595 337501 282607 337504
rect 282549 337495 282607 337501
rect 282914 337492 282920 337504
rect 282972 337492 282978 337544
rect 283469 337535 283527 337541
rect 283469 337501 283481 337535
rect 283515 337532 283527 337535
rect 284110 337532 284116 337544
rect 283515 337504 284116 337532
rect 283515 337501 283527 337504
rect 283469 337495 283527 337501
rect 284110 337492 284116 337504
rect 284168 337492 284174 337544
rect 285030 337492 285036 337544
rect 285088 337532 285094 337544
rect 580902 337532 580908 337544
rect 285088 337504 580908 337532
rect 285088 337492 285094 337504
rect 580902 337492 580908 337504
rect 580960 337492 580966 337544
rect 234706 337424 234712 337476
rect 234764 337464 234770 337476
rect 530670 337464 530676 337476
rect 234764 337436 530676 337464
rect 234764 337424 234770 337436
rect 530670 337424 530676 337436
rect 530728 337424 530734 337476
rect 233510 337356 233516 337408
rect 233568 337396 233574 337408
rect 538306 337396 538312 337408
rect 233568 337368 538312 337396
rect 233568 337356 233574 337368
rect 538306 337356 538312 337368
rect 538364 337356 538370 337408
rect 232498 337288 232504 337340
rect 232556 337328 232562 337340
rect 239401 337331 239459 337337
rect 239401 337328 239413 337331
rect 232556 337300 239413 337328
rect 232556 337288 232562 337300
rect 239401 337297 239413 337300
rect 239447 337297 239459 337331
rect 239401 337291 239459 337297
rect 250809 337331 250867 337337
rect 250809 337297 250821 337331
rect 250855 337328 250867 337331
rect 250898 337328 250904 337340
rect 250855 337300 250904 337328
rect 250855 337297 250867 337300
rect 250809 337291 250867 337297
rect 250898 337288 250904 337300
rect 250956 337288 250962 337340
rect 250993 337331 251051 337337
rect 250993 337297 251005 337331
rect 251039 337328 251051 337331
rect 251082 337328 251088 337340
rect 251039 337300 251088 337328
rect 251039 337297 251051 337300
rect 250993 337291 251051 337297
rect 251082 337288 251088 337300
rect 251140 337288 251146 337340
rect 254213 337331 254271 337337
rect 254213 337297 254225 337331
rect 254259 337328 254271 337331
rect 254394 337328 254400 337340
rect 254259 337300 254400 337328
rect 254259 337297 254271 337300
rect 254213 337291 254271 337297
rect 254394 337288 254400 337300
rect 254452 337288 254458 337340
rect 254489 337331 254547 337337
rect 254489 337297 254501 337331
rect 254535 337328 254547 337331
rect 254854 337328 254860 337340
rect 254535 337300 254860 337328
rect 254535 337297 254547 337300
rect 254489 337291 254547 337297
rect 254854 337288 254860 337300
rect 254912 337288 254918 337340
rect 254946 337288 254952 337340
rect 255004 337328 255010 337340
rect 255133 337331 255191 337337
rect 255133 337328 255145 337331
rect 255004 337300 255145 337328
rect 255004 337288 255010 337300
rect 255133 337297 255145 337300
rect 255179 337297 255191 337331
rect 255133 337291 255191 337297
rect 255590 337288 255596 337340
rect 255648 337328 255654 337340
rect 255777 337331 255835 337337
rect 255777 337328 255789 337331
rect 255648 337300 255789 337328
rect 255648 337288 255654 337300
rect 255777 337297 255789 337300
rect 255823 337297 255835 337331
rect 255777 337291 255835 337297
rect 265253 337331 265311 337337
rect 265253 337297 265265 337331
rect 265299 337328 265311 337331
rect 268933 337331 268991 337337
rect 268933 337328 268945 337331
rect 265299 337300 268945 337328
rect 265299 337297 265311 337300
rect 265253 337291 265311 337297
rect 268933 337297 268945 337300
rect 268979 337297 268991 337331
rect 268933 337291 268991 337297
rect 275646 337288 275652 337340
rect 275704 337328 275710 337340
rect 275741 337331 275799 337337
rect 275741 337328 275753 337331
rect 275704 337300 275753 337328
rect 275704 337288 275710 337300
rect 275741 337297 275753 337300
rect 275787 337297 275799 337331
rect 278130 337328 278136 337340
rect 278091 337300 278136 337328
rect 275741 337291 275799 337297
rect 278130 337288 278136 337300
rect 278188 337288 278194 337340
rect 278958 337288 278964 337340
rect 279016 337328 279022 337340
rect 292761 337331 292819 337337
rect 292761 337328 292773 337331
rect 279016 337300 292773 337328
rect 279016 337288 279022 337300
rect 292761 337297 292773 337300
rect 292807 337297 292819 337331
rect 292761 337291 292819 337297
rect 293788 337300 299474 337328
rect 236178 337260 236184 337272
rect 236139 337232 236184 337260
rect 236178 337220 236184 337232
rect 236236 337220 236242 337272
rect 237558 337220 237564 337272
rect 237616 337260 237622 337272
rect 237837 337263 237895 337269
rect 237837 337260 237849 337263
rect 237616 337232 237849 337260
rect 237616 337220 237622 337232
rect 237837 337229 237849 337232
rect 237883 337229 237895 337263
rect 237837 337223 237895 337229
rect 265713 337263 265771 337269
rect 265713 337229 265725 337263
rect 265759 337260 265771 337263
rect 268841 337263 268899 337269
rect 268841 337260 268853 337263
rect 265759 337232 268853 337260
rect 265759 337229 265771 337232
rect 265713 337223 265771 337229
rect 268841 337229 268853 337232
rect 268887 337229 268899 337263
rect 268841 337223 268899 337229
rect 270037 337263 270095 337269
rect 270037 337229 270049 337263
rect 270083 337260 270095 337263
rect 293788 337260 293816 337300
rect 270083 337232 293816 337260
rect 299446 337260 299474 337300
rect 420914 337260 420920 337272
rect 299446 337232 420920 337260
rect 270083 337229 270095 337232
rect 270037 337223 270095 337229
rect 420914 337220 420920 337232
rect 420972 337220 420978 337272
rect 254762 337152 254768 337204
rect 254820 337192 254826 337204
rect 254949 337195 255007 337201
rect 254949 337192 254961 337195
rect 254820 337164 254961 337192
rect 254820 337152 254826 337164
rect 254949 337161 254961 337164
rect 254995 337161 255007 337195
rect 254949 337155 255007 337161
rect 266906 337152 266912 337204
rect 266964 337192 266970 337204
rect 268749 337195 268807 337201
rect 268749 337192 268761 337195
rect 266964 337164 268761 337192
rect 266964 337152 266970 337164
rect 268749 337161 268761 337164
rect 268795 337161 268807 337195
rect 268749 337155 268807 337161
rect 269209 337195 269267 337201
rect 269209 337161 269221 337195
rect 269255 337192 269267 337195
rect 269298 337192 269304 337204
rect 269255 337164 269304 337192
rect 269255 337161 269267 337164
rect 269209 337155 269267 337161
rect 269298 337152 269304 337164
rect 269356 337152 269362 337204
rect 273530 337152 273536 337204
rect 273588 337192 273594 337204
rect 292761 337195 292819 337201
rect 273588 337164 279096 337192
rect 273588 337152 273594 337164
rect 271969 337127 272027 337133
rect 271969 337093 271981 337127
rect 272015 337124 272027 337127
rect 277305 337127 277363 337133
rect 277305 337124 277317 337127
rect 272015 337096 277317 337124
rect 272015 337093 272027 337096
rect 271969 337087 272027 337093
rect 277305 337093 277317 337096
rect 277351 337093 277363 337127
rect 277305 337087 277363 337093
rect 277581 337127 277639 337133
rect 277581 337093 277593 337127
rect 277627 337124 277639 337127
rect 278590 337124 278596 337136
rect 277627 337096 278596 337124
rect 277627 337093 277639 337096
rect 277581 337087 277639 337093
rect 278590 337084 278596 337096
rect 278648 337084 278654 337136
rect 279068 337124 279096 337164
rect 292761 337161 292773 337195
rect 292807 337192 292819 337195
rect 536834 337192 536840 337204
rect 292807 337164 536840 337192
rect 292807 337161 292819 337164
rect 292761 337155 292819 337161
rect 536834 337152 536840 337164
rect 536892 337152 536898 337204
rect 279068 337096 279464 337124
rect 268013 337059 268071 337065
rect 268013 337025 268025 337059
rect 268059 337056 268071 337059
rect 273073 337059 273131 337065
rect 273073 337056 273085 337059
rect 268059 337028 273085 337056
rect 268059 337025 268071 337028
rect 268013 337019 268071 337025
rect 273073 337025 273085 337028
rect 273119 337025 273131 337059
rect 273073 337019 273131 337025
rect 279142 337016 279148 337068
rect 279200 337056 279206 337068
rect 279326 337056 279332 337068
rect 279200 337028 279332 337056
rect 279200 337016 279206 337028
rect 279326 337016 279332 337028
rect 279384 337016 279390 337068
rect 279436 337056 279464 337096
rect 279510 337084 279516 337136
rect 279568 337124 279574 337136
rect 287517 337127 287575 337133
rect 287517 337124 287529 337127
rect 279568 337096 287529 337124
rect 279568 337084 279574 337096
rect 287517 337093 287529 337096
rect 287563 337093 287575 337127
rect 287517 337087 287575 337093
rect 288069 337127 288127 337133
rect 288069 337093 288081 337127
rect 288115 337124 288127 337127
rect 538214 337124 538220 337136
rect 288115 337096 538220 337124
rect 288115 337093 288127 337096
rect 288069 337087 288127 337093
rect 538214 337084 538220 337096
rect 538272 337084 538278 337136
rect 279881 337059 279939 337065
rect 279881 337056 279893 337059
rect 279436 337028 279893 337056
rect 279881 337025 279893 337028
rect 279927 337025 279939 337059
rect 282914 337056 282920 337068
rect 282875 337028 282920 337056
rect 279881 337019 279939 337025
rect 282914 337016 282920 337028
rect 282972 337016 282978 337068
rect 283282 337016 283288 337068
rect 283340 337056 283346 337068
rect 283650 337056 283656 337068
rect 283340 337028 283656 337056
rect 283340 337016 283346 337028
rect 283650 337016 283656 337028
rect 283708 337016 283714 337068
rect 538858 337056 538864 337068
rect 283760 337028 538864 337056
rect 241701 336991 241759 336997
rect 241701 336957 241713 336991
rect 241747 336988 241759 336991
rect 242710 336988 242716 337000
rect 241747 336960 242716 336988
rect 241747 336957 241759 336960
rect 241701 336951 241759 336957
rect 242710 336948 242716 336960
rect 242768 336948 242774 337000
rect 265066 336948 265072 337000
rect 265124 336988 265130 337000
rect 268197 336991 268255 336997
rect 268197 336988 268209 336991
rect 265124 336960 268209 336988
rect 265124 336948 265130 336960
rect 268197 336957 268209 336960
rect 268243 336957 268255 336991
rect 268197 336951 268255 336957
rect 272797 336991 272855 336997
rect 272797 336957 272809 336991
rect 272843 336988 272855 336991
rect 274269 336991 274327 336997
rect 274269 336988 274281 336991
rect 272843 336960 274281 336988
rect 272843 336957 272855 336960
rect 272797 336951 272855 336957
rect 274269 336957 274281 336960
rect 274315 336957 274327 336991
rect 274269 336951 274327 336957
rect 276290 336948 276296 337000
rect 276348 336988 276354 337000
rect 276750 336988 276756 337000
rect 276348 336960 276756 336988
rect 276348 336948 276354 336960
rect 276750 336948 276756 336960
rect 276808 336948 276814 337000
rect 276845 336991 276903 336997
rect 276845 336957 276857 336991
rect 276891 336988 276903 336991
rect 276934 336988 276940 337000
rect 276891 336960 276940 336988
rect 276891 336957 276903 336960
rect 276845 336951 276903 336957
rect 276934 336948 276940 336960
rect 276992 336948 276998 337000
rect 281169 336991 281227 336997
rect 281169 336957 281181 336991
rect 281215 336988 281227 336991
rect 283760 336988 283788 337028
rect 538858 337016 538864 337028
rect 538916 337016 538922 337068
rect 281215 336960 283788 336988
rect 281215 336957 281227 336960
rect 281169 336951 281227 336957
rect 287606 336948 287612 337000
rect 287664 336988 287670 337000
rect 538950 336988 538956 337000
rect 287664 336960 538956 336988
rect 287664 336948 287670 336960
rect 538950 336948 538956 336960
rect 539008 336948 539014 337000
rect 237834 336920 237840 336932
rect 219406 336892 237840 336920
rect 33134 336744 33140 336796
rect 33192 336784 33198 336796
rect 219406 336784 219434 336892
rect 237834 336880 237840 336892
rect 237892 336880 237898 336932
rect 243725 336923 243783 336929
rect 243725 336889 243737 336923
rect 243771 336920 243783 336923
rect 243906 336920 243912 336932
rect 243771 336892 243912 336920
rect 243771 336889 243783 336892
rect 243725 336883 243783 336889
rect 243906 336880 243912 336892
rect 243964 336880 243970 336932
rect 264606 336880 264612 336932
rect 264664 336920 264670 336932
rect 272981 336923 273039 336929
rect 272981 336920 272993 336923
rect 264664 336892 272993 336920
rect 264664 336880 264670 336892
rect 272981 336889 272993 336892
rect 273027 336889 273039 336923
rect 272981 336883 273039 336889
rect 275370 336880 275376 336932
rect 275428 336920 275434 336932
rect 279973 336923 280031 336929
rect 279973 336920 279985 336923
rect 275428 336892 279985 336920
rect 275428 336880 275434 336892
rect 279973 336889 279985 336892
rect 280019 336889 280031 336923
rect 279973 336883 280031 336889
rect 283006 336880 283012 336932
rect 283064 336920 283070 336932
rect 285217 336923 285275 336929
rect 285217 336920 285229 336923
rect 283064 336892 285229 336920
rect 283064 336880 283070 336892
rect 285217 336889 285229 336892
rect 285263 336889 285275 336923
rect 285217 336883 285275 336889
rect 287517 336923 287575 336929
rect 287517 336889 287529 336923
rect 287563 336920 287575 336923
rect 543734 336920 543740 336932
rect 287563 336892 543740 336920
rect 287563 336889 287575 336892
rect 287517 336883 287575 336889
rect 543734 336880 543740 336892
rect 543792 336880 543798 336932
rect 237374 336812 237380 336864
rect 237432 336852 237438 336864
rect 242253 336855 242311 336861
rect 242253 336852 242265 336855
rect 237432 336824 242265 336852
rect 237432 336812 237438 336824
rect 242253 336821 242265 336824
rect 242299 336821 242311 336855
rect 242253 336815 242311 336821
rect 269206 336812 269212 336864
rect 269264 336852 269270 336864
rect 273257 336855 273315 336861
rect 273257 336852 273269 336855
rect 269264 336824 270494 336852
rect 269264 336812 269270 336824
rect 33192 336756 219434 336784
rect 33192 336744 33198 336756
rect 240410 336744 240416 336796
rect 240468 336784 240474 336796
rect 240686 336784 240692 336796
rect 240468 336756 240692 336784
rect 240468 336744 240474 336756
rect 240686 336744 240692 336756
rect 240744 336744 240750 336796
rect 241606 336784 241612 336796
rect 241567 336756 241612 336784
rect 241606 336744 241612 336756
rect 241664 336744 241670 336796
rect 263229 336787 263287 336793
rect 263229 336753 263241 336787
rect 263275 336784 263287 336787
rect 266998 336784 267004 336796
rect 263275 336756 267004 336784
rect 263275 336753 263287 336756
rect 263229 336747 263287 336753
rect 266998 336744 267004 336756
rect 267056 336744 267062 336796
rect 267384 336756 268976 336784
rect 103422 336676 103428 336728
rect 103480 336716 103486 336728
rect 238941 336719 238999 336725
rect 238941 336716 238953 336719
rect 103480 336688 238953 336716
rect 103480 336676 103486 336688
rect 238941 336685 238953 336688
rect 238987 336685 238999 336719
rect 238941 336679 238999 336685
rect 240134 336676 240140 336728
rect 240192 336716 240198 336728
rect 247770 336716 247776 336728
rect 240192 336688 247776 336716
rect 240192 336676 240198 336688
rect 247770 336676 247776 336688
rect 247828 336676 247834 336728
rect 259825 336719 259883 336725
rect 259825 336685 259837 336719
rect 259871 336716 259883 336719
rect 263318 336716 263324 336728
rect 259871 336688 263324 336716
rect 259871 336685 259883 336688
rect 259825 336679 259883 336685
rect 263318 336676 263324 336688
rect 263376 336676 263382 336728
rect 266262 336676 266268 336728
rect 266320 336716 266326 336728
rect 267384 336716 267412 336756
rect 266320 336688 267412 336716
rect 268948 336716 268976 336756
rect 269117 336719 269175 336725
rect 269117 336716 269129 336719
rect 268948 336688 269129 336716
rect 266320 336676 266326 336688
rect 269117 336685 269129 336688
rect 269163 336685 269175 336719
rect 270466 336716 270494 336824
rect 272904 336824 273269 336852
rect 272904 336716 272932 336824
rect 273257 336821 273269 336824
rect 273303 336821 273315 336855
rect 273257 336815 273315 336821
rect 275094 336812 275100 336864
rect 275152 336852 275158 336864
rect 277029 336855 277087 336861
rect 277029 336852 277041 336855
rect 275152 336824 277041 336852
rect 275152 336812 275158 336824
rect 277029 336821 277041 336824
rect 277075 336821 277087 336855
rect 277394 336852 277400 336864
rect 277355 336824 277400 336852
rect 277029 336815 277087 336821
rect 277394 336812 277400 336824
rect 277452 336812 277458 336864
rect 279602 336812 279608 336864
rect 279660 336852 279666 336864
rect 279697 336855 279755 336861
rect 279697 336852 279709 336855
rect 279660 336824 279709 336852
rect 279660 336812 279666 336824
rect 279697 336821 279709 336824
rect 279743 336821 279755 336855
rect 279697 336815 279755 336821
rect 280709 336855 280767 336861
rect 280709 336821 280721 336855
rect 280755 336852 280767 336855
rect 557534 336852 557540 336864
rect 280755 336824 557540 336852
rect 280755 336821 280767 336824
rect 280709 336815 280767 336821
rect 557534 336812 557540 336824
rect 557592 336812 557598 336864
rect 273165 336787 273223 336793
rect 273165 336753 273177 336787
rect 273211 336784 273223 336787
rect 273717 336787 273775 336793
rect 273717 336784 273729 336787
rect 273211 336756 273729 336784
rect 273211 336753 273223 336756
rect 273165 336747 273223 336753
rect 273717 336753 273729 336756
rect 273763 336753 273775 336787
rect 273717 336747 273775 336753
rect 273809 336787 273867 336793
rect 273809 336753 273821 336787
rect 273855 336784 273867 336787
rect 274266 336784 274272 336796
rect 273855 336756 274272 336784
rect 273855 336753 273867 336756
rect 273809 336747 273867 336753
rect 274266 336744 274272 336756
rect 274324 336744 274330 336796
rect 274726 336744 274732 336796
rect 274784 336784 274790 336796
rect 279510 336784 279516 336796
rect 274784 336756 279516 336784
rect 274784 336744 274790 336756
rect 279510 336744 279516 336756
rect 279568 336744 279574 336796
rect 287701 336787 287759 336793
rect 287701 336753 287713 336787
rect 287747 336784 287759 336787
rect 561674 336784 561680 336796
rect 287747 336756 561680 336784
rect 287747 336753 287759 336756
rect 287701 336747 287759 336753
rect 561674 336744 561680 336756
rect 561732 336744 561738 336796
rect 270466 336688 272932 336716
rect 273073 336719 273131 336725
rect 269117 336679 269175 336685
rect 273073 336685 273085 336719
rect 273119 336716 273131 336719
rect 341518 336716 341524 336728
rect 273119 336688 341524 336716
rect 273119 336685 273131 336688
rect 273073 336679 273131 336685
rect 341518 336676 341524 336688
rect 341576 336676 341582 336728
rect 96522 336608 96528 336660
rect 96580 336648 96586 336660
rect 242802 336648 242808 336660
rect 96580 336620 242808 336648
rect 96580 336608 96586 336620
rect 242802 336608 242808 336620
rect 242860 336608 242866 336660
rect 249058 336608 249064 336660
rect 249116 336648 249122 336660
rect 254118 336648 254124 336660
rect 249116 336620 254124 336648
rect 249116 336608 249122 336620
rect 254118 336608 254124 336620
rect 254176 336608 254182 336660
rect 259270 336608 259276 336660
rect 259328 336648 259334 336660
rect 261389 336651 261447 336657
rect 261389 336648 261401 336651
rect 259328 336620 261401 336648
rect 259328 336608 259334 336620
rect 261389 336617 261401 336620
rect 261435 336617 261447 336651
rect 261389 336611 261447 336617
rect 263962 336608 263968 336660
rect 264020 336648 264026 336660
rect 268013 336651 268071 336657
rect 268013 336648 268025 336651
rect 264020 336620 268025 336648
rect 264020 336608 264026 336620
rect 268013 336617 268025 336620
rect 268059 336617 268071 336651
rect 268013 336611 268071 336617
rect 268102 336608 268108 336660
rect 268160 336648 268166 336660
rect 272797 336651 272855 336657
rect 272797 336648 272809 336651
rect 268160 336620 268700 336648
rect 268160 336608 268166 336620
rect 95142 336540 95148 336592
rect 95200 336580 95206 336592
rect 242161 336583 242219 336589
rect 242161 336580 242173 336583
rect 95200 336552 242173 336580
rect 95200 336540 95206 336552
rect 242161 336549 242173 336552
rect 242207 336549 242219 336583
rect 242161 336543 242219 336549
rect 242253 336583 242311 336589
rect 242253 336549 242265 336583
rect 242299 336580 242311 336583
rect 243909 336583 243967 336589
rect 243909 336580 243921 336583
rect 242299 336552 243921 336580
rect 242299 336549 242311 336552
rect 242253 336543 242311 336549
rect 243909 336549 243921 336552
rect 243955 336549 243967 336583
rect 243909 336543 243967 336549
rect 259914 336540 259920 336592
rect 259972 336580 259978 336592
rect 263229 336583 263287 336589
rect 263229 336580 263241 336583
rect 259972 336552 263241 336580
rect 259972 336540 259978 336552
rect 263229 336549 263241 336552
rect 263275 336549 263287 336583
rect 268672 336580 268700 336620
rect 268948 336620 272809 336648
rect 268948 336580 268976 336620
rect 272797 336617 272809 336620
rect 272843 336617 272855 336651
rect 272797 336611 272855 336617
rect 272981 336651 273039 336657
rect 272981 336617 272993 336651
rect 273027 336648 273039 336651
rect 344278 336648 344284 336660
rect 273027 336620 344284 336648
rect 273027 336617 273039 336620
rect 272981 336611 273039 336617
rect 344278 336608 344284 336620
rect 344336 336608 344342 336660
rect 268672 336552 268976 336580
rect 269209 336583 269267 336589
rect 263229 336543 263287 336549
rect 269209 336549 269221 336583
rect 269255 336580 269267 336583
rect 273165 336583 273223 336589
rect 269255 336552 273116 336580
rect 269255 336549 269267 336552
rect 269209 336543 269267 336549
rect 46842 336472 46848 336524
rect 46900 336512 46906 336524
rect 238757 336515 238815 336521
rect 238757 336512 238769 336515
rect 46900 336484 238769 336512
rect 46900 336472 46906 336484
rect 238757 336481 238769 336484
rect 238803 336481 238815 336515
rect 241241 336515 241299 336521
rect 241241 336512 241253 336515
rect 238757 336475 238815 336481
rect 238864 336484 241253 336512
rect 78582 336404 78588 336456
rect 78640 336444 78646 336456
rect 238864 336444 238892 336484
rect 241241 336481 241253 336484
rect 241287 336481 241299 336515
rect 241241 336475 241299 336481
rect 241333 336515 241391 336521
rect 241333 336481 241345 336515
rect 241379 336512 241391 336515
rect 243446 336512 243452 336524
rect 241379 336484 243452 336512
rect 241379 336481 241391 336484
rect 241333 336475 241391 336481
rect 243446 336472 243452 336484
rect 243504 336472 243510 336524
rect 259641 336515 259699 336521
rect 259641 336481 259653 336515
rect 259687 336512 259699 336515
rect 263045 336515 263103 336521
rect 263045 336512 263057 336515
rect 259687 336484 263057 336512
rect 259687 336481 259699 336484
rect 259641 336475 259699 336481
rect 263045 336481 263057 336484
rect 263091 336481 263103 336515
rect 263045 336475 263103 336481
rect 267458 336472 267464 336524
rect 267516 336512 267522 336524
rect 272981 336515 273039 336521
rect 272981 336512 272993 336515
rect 267516 336484 272993 336512
rect 267516 336472 267522 336484
rect 272981 336481 272993 336484
rect 273027 336481 273039 336515
rect 273088 336512 273116 336552
rect 273165 336549 273177 336583
rect 273211 336580 273223 336583
rect 348418 336580 348424 336592
rect 273211 336552 348424 336580
rect 273211 336549 273223 336552
rect 273165 336543 273223 336549
rect 348418 336540 348424 336552
rect 348476 336540 348482 336592
rect 274177 336515 274235 336521
rect 273088 336484 273346 336512
rect 272981 336475 273039 336481
rect 78640 336416 238892 336444
rect 238941 336447 238999 336453
rect 78640 336404 78646 336416
rect 238941 336413 238953 336447
rect 238987 336444 238999 336447
rect 238987 336416 240364 336444
rect 238987 336413 238999 336416
rect 238941 336407 238999 336413
rect 45462 336336 45468 336388
rect 45520 336376 45526 336388
rect 238573 336379 238631 336385
rect 238573 336376 238585 336379
rect 45520 336348 238585 336376
rect 45520 336336 45526 336348
rect 238573 336345 238585 336348
rect 238619 336345 238631 336379
rect 238573 336339 238631 336345
rect 238846 336336 238852 336388
rect 238904 336376 238910 336388
rect 239493 336379 239551 336385
rect 239493 336376 239505 336379
rect 238904 336348 239505 336376
rect 238904 336336 238910 336348
rect 239493 336345 239505 336348
rect 239539 336345 239551 336379
rect 239493 336339 239551 336345
rect 240226 336336 240232 336388
rect 240284 336336 240290 336388
rect 240336 336376 240364 336416
rect 240686 336404 240692 336456
rect 240744 336444 240750 336456
rect 244182 336444 244188 336456
rect 240744 336416 244188 336444
rect 240744 336404 240750 336416
rect 244182 336404 244188 336416
rect 244240 336404 244246 336456
rect 263410 336404 263416 336456
rect 263468 336444 263474 336456
rect 272613 336447 272671 336453
rect 272613 336444 272625 336447
rect 263468 336416 272625 336444
rect 263468 336404 263474 336416
rect 272613 336413 272625 336416
rect 272659 336413 272671 336447
rect 273318 336444 273346 336484
rect 274177 336481 274189 336515
rect 274223 336512 274235 336515
rect 355318 336512 355324 336524
rect 274223 336484 355324 336512
rect 274223 336481 274235 336484
rect 274177 336475 274235 336481
rect 355318 336472 355324 336484
rect 355376 336472 355382 336524
rect 362218 336444 362224 336456
rect 273318 336416 362224 336444
rect 272613 336407 272671 336413
rect 362218 336404 362224 336416
rect 362276 336404 362282 336456
rect 241333 336379 241391 336385
rect 241333 336376 241345 336379
rect 240336 336348 241345 336376
rect 241333 336345 241345 336348
rect 241379 336345 241391 336379
rect 241333 336339 241391 336345
rect 243446 336336 243452 336388
rect 243504 336376 243510 336388
rect 245105 336379 245163 336385
rect 245105 336376 245117 336379
rect 243504 336348 245117 336376
rect 243504 336336 243510 336348
rect 245105 336345 245117 336348
rect 245151 336345 245163 336379
rect 245105 336339 245163 336345
rect 261110 336336 261116 336388
rect 261168 336376 261174 336388
rect 272797 336379 272855 336385
rect 272797 336376 272809 336379
rect 261168 336348 272809 336376
rect 261168 336336 261174 336348
rect 272797 336345 272809 336348
rect 272843 336345 272855 336379
rect 369118 336376 369124 336388
rect 272797 336339 272855 336345
rect 273180 336348 369124 336376
rect 89622 336268 89628 336320
rect 89680 336308 89686 336320
rect 237285 336311 237343 336317
rect 237285 336308 237297 336311
rect 89680 336280 237297 336308
rect 89680 336268 89686 336280
rect 237285 336277 237297 336280
rect 237331 336277 237343 336311
rect 240244 336308 240272 336336
rect 237285 336271 237343 336277
rect 237392 336280 240272 336308
rect 64782 336200 64788 336252
rect 64840 336240 64846 336252
rect 237392 336240 237420 336280
rect 261662 336268 261668 336320
rect 261720 336308 261726 336320
rect 264238 336308 264244 336320
rect 261720 336280 264244 336308
rect 261720 336268 261726 336280
rect 264238 336268 264244 336280
rect 264296 336268 264302 336320
rect 267734 336268 267740 336320
rect 267792 336308 267798 336320
rect 268378 336308 268384 336320
rect 267792 336280 268384 336308
rect 267792 336268 267798 336280
rect 268378 336268 268384 336280
rect 268436 336268 268442 336320
rect 268749 336311 268807 336317
rect 268749 336277 268761 336311
rect 268795 336308 268807 336311
rect 273180 336308 273208 336348
rect 369118 336336 369124 336348
rect 369176 336336 369182 336388
rect 268795 336280 273208 336308
rect 273717 336311 273775 336317
rect 268795 336277 268807 336280
rect 268749 336271 268807 336277
rect 273717 336277 273729 336311
rect 273763 336308 273775 336311
rect 376018 336308 376024 336320
rect 273763 336280 376024 336308
rect 273763 336277 273775 336280
rect 273717 336271 273775 336277
rect 376018 336268 376024 336280
rect 376076 336268 376082 336320
rect 64840 336212 237420 336240
rect 64840 336200 64846 336212
rect 237834 336200 237840 336252
rect 237892 336240 237898 336252
rect 239401 336243 239459 336249
rect 239401 336240 239413 336243
rect 237892 336212 239413 336240
rect 237892 336200 237898 336212
rect 239401 336209 239413 336212
rect 239447 336209 239459 336243
rect 239401 336203 239459 336209
rect 240226 336200 240232 336252
rect 240284 336240 240290 336252
rect 248690 336240 248696 336252
rect 240284 336212 248696 336240
rect 240284 336200 240290 336212
rect 248690 336200 248696 336212
rect 248748 336200 248754 336252
rect 257985 336243 258043 336249
rect 257985 336209 257997 336243
rect 258031 336240 258043 336243
rect 260834 336240 260840 336252
rect 258031 336212 260840 336240
rect 258031 336209 258043 336212
rect 257985 336203 258043 336209
rect 260834 336200 260840 336212
rect 260892 336200 260898 336252
rect 262214 336200 262220 336252
rect 262272 336240 262278 336252
rect 263502 336240 263508 336252
rect 262272 336212 263508 336240
rect 262272 336200 262278 336212
rect 263502 336200 263508 336212
rect 263560 336200 263566 336252
rect 265710 336200 265716 336252
rect 265768 336240 265774 336252
rect 265768 336212 268148 336240
rect 265768 336200 265774 336212
rect 39942 336132 39948 336184
rect 40000 336172 40006 336184
rect 238110 336172 238116 336184
rect 40000 336144 238116 336172
rect 40000 336132 40006 336144
rect 238110 336132 238116 336144
rect 238168 336132 238174 336184
rect 238202 336132 238208 336184
rect 238260 336172 238266 336184
rect 238849 336175 238907 336181
rect 238849 336172 238861 336175
rect 238260 336144 238861 336172
rect 238260 336132 238266 336144
rect 238849 336141 238861 336144
rect 238895 336141 238907 336175
rect 238849 336135 238907 336141
rect 239217 336175 239275 336181
rect 239217 336141 239229 336175
rect 239263 336172 239275 336175
rect 243722 336172 243728 336184
rect 239263 336144 243728 336172
rect 239263 336141 239275 336144
rect 239217 336135 239275 336141
rect 243722 336132 243728 336144
rect 243780 336132 243786 336184
rect 261938 336132 261944 336184
rect 261996 336172 262002 336184
rect 267274 336172 267280 336184
rect 261996 336144 267280 336172
rect 261996 336132 262002 336144
rect 267274 336132 267280 336144
rect 267332 336132 267338 336184
rect 24762 336064 24768 336116
rect 24820 336104 24826 336116
rect 236914 336104 236920 336116
rect 24820 336076 236920 336104
rect 24820 336064 24826 336076
rect 236914 336064 236920 336076
rect 236972 336064 236978 336116
rect 238754 336064 238760 336116
rect 238812 336104 238818 336116
rect 252005 336107 252063 336113
rect 252005 336104 252017 336107
rect 238812 336076 252017 336104
rect 238812 336064 238818 336076
rect 252005 336073 252017 336076
rect 252051 336073 252063 336107
rect 252005 336067 252063 336073
rect 260282 336064 260288 336116
rect 260340 336104 260346 336116
rect 260340 336076 262904 336104
rect 260340 336064 260346 336076
rect 233602 335996 233608 336048
rect 233660 336036 233666 336048
rect 237193 336039 237251 336045
rect 237193 336036 237205 336039
rect 233660 336008 237205 336036
rect 233660 335996 233666 336008
rect 237193 336005 237205 336008
rect 237239 336005 237251 336039
rect 237193 335999 237251 336005
rect 237285 336039 237343 336045
rect 237285 336005 237297 336039
rect 237331 336036 237343 336039
rect 242250 336036 242256 336048
rect 237331 336008 242256 336036
rect 237331 336005 237343 336008
rect 237285 335999 237343 336005
rect 242250 335996 242256 336008
rect 242308 335996 242314 336048
rect 242802 335996 242808 336048
rect 242860 336036 242866 336048
rect 243817 336039 243875 336045
rect 243817 336036 243829 336039
rect 242860 336008 243829 336036
rect 242860 335996 242866 336008
rect 243817 336005 243829 336008
rect 243863 336005 243875 336039
rect 243817 335999 243875 336005
rect 243909 336039 243967 336045
rect 243909 336005 243921 336039
rect 243955 336036 243967 336039
rect 256786 336036 256792 336048
rect 243955 336008 256792 336036
rect 243955 336005 243967 336008
rect 243909 335999 243967 336005
rect 256786 335996 256792 336008
rect 256844 335996 256850 336048
rect 257341 336039 257399 336045
rect 257341 336005 257353 336039
rect 257387 336036 257399 336039
rect 257387 336008 262812 336036
rect 257387 336005 257399 336008
rect 257341 335999 257399 336005
rect 117222 335928 117228 335980
rect 117280 335968 117286 335980
rect 244458 335968 244464 335980
rect 117280 335940 244464 335968
rect 117280 335928 117286 335940
rect 244458 335928 244464 335940
rect 244516 335928 244522 335980
rect 244553 335971 244611 335977
rect 244553 335937 244565 335971
rect 244599 335968 244611 335971
rect 250622 335968 250628 335980
rect 244599 335940 250628 335968
rect 244599 335937 244611 335940
rect 244553 335931 244611 335937
rect 250622 335928 250628 335940
rect 250680 335928 250686 335980
rect 262030 335968 262036 335980
rect 261991 335940 262036 335968
rect 262030 335928 262036 335940
rect 262088 335928 262094 335980
rect 119982 335860 119988 335912
rect 120040 335900 120046 335912
rect 239033 335903 239091 335909
rect 239033 335900 239045 335903
rect 120040 335872 239045 335900
rect 120040 335860 120046 335872
rect 239033 335869 239045 335872
rect 239079 335869 239091 335903
rect 239033 335863 239091 335869
rect 239122 335860 239128 335912
rect 239180 335900 239186 335912
rect 244369 335903 244427 335909
rect 244369 335900 244381 335903
rect 239180 335872 244381 335900
rect 239180 335860 239186 335872
rect 244369 335869 244381 335872
rect 244415 335869 244427 335903
rect 244369 335863 244427 335869
rect 244829 335903 244887 335909
rect 244829 335869 244841 335903
rect 244875 335900 244887 335903
rect 251542 335900 251548 335912
rect 244875 335872 251548 335900
rect 244875 335869 244887 335872
rect 244829 335863 244887 335869
rect 251542 335860 251548 335872
rect 251600 335860 251606 335912
rect 255958 335860 255964 335912
rect 256016 335900 256022 335912
rect 259454 335900 259460 335912
rect 256016 335872 259460 335900
rect 256016 335860 256022 335872
rect 259454 335860 259460 335872
rect 259512 335860 259518 335912
rect 262784 335900 262812 336008
rect 262876 335968 262904 336076
rect 262950 336064 262956 336116
rect 263008 336104 263014 336116
rect 268013 336107 268071 336113
rect 268013 336104 268025 336107
rect 263008 336076 268025 336104
rect 263008 336064 263014 336076
rect 268013 336073 268025 336076
rect 268059 336073 268071 336107
rect 268120 336104 268148 336212
rect 269390 336200 269396 336252
rect 269448 336240 269454 336252
rect 270310 336240 270316 336252
rect 269448 336212 270316 336240
rect 269448 336200 269454 336212
rect 270310 336200 270316 336212
rect 270368 336200 270374 336252
rect 274177 336243 274235 336249
rect 274177 336240 274189 336243
rect 272352 336212 274189 336240
rect 268381 336175 268439 336181
rect 268381 336141 268393 336175
rect 268427 336172 268439 336175
rect 272153 336175 272211 336181
rect 272153 336172 272165 336175
rect 268427 336144 272165 336172
rect 268427 336141 268439 336144
rect 268381 336135 268439 336141
rect 272153 336141 272165 336144
rect 272199 336141 272211 336175
rect 272153 336135 272211 336141
rect 272352 336104 272380 336212
rect 274177 336209 274189 336212
rect 274223 336209 274235 336243
rect 274177 336203 274235 336209
rect 274269 336243 274327 336249
rect 274269 336209 274281 336243
rect 274315 336240 274327 336243
rect 382918 336240 382924 336252
rect 274315 336212 382924 336240
rect 274315 336209 274327 336212
rect 274269 336203 274327 336209
rect 382918 336200 382924 336212
rect 382976 336200 382982 336252
rect 272429 336175 272487 336181
rect 272429 336141 272441 336175
rect 272475 336172 272487 336175
rect 391198 336172 391204 336184
rect 272475 336144 391204 336172
rect 272475 336141 272487 336144
rect 272429 336135 272487 336141
rect 391198 336132 391204 336144
rect 391256 336132 391262 336184
rect 268120 336076 272380 336104
rect 272613 336107 272671 336113
rect 268013 336067 268071 336073
rect 272613 336073 272625 336107
rect 272659 336104 272671 336107
rect 273257 336107 273315 336113
rect 272659 336076 273116 336104
rect 272659 336073 272671 336076
rect 272613 336067 272671 336073
rect 263045 336039 263103 336045
rect 263045 336005 263057 336039
rect 263091 336036 263103 336039
rect 267734 336036 267740 336048
rect 263091 336008 267740 336036
rect 263091 336005 263103 336008
rect 263045 335999 263103 336005
rect 267734 335996 267740 336008
rect 267792 335996 267798 336048
rect 269482 335996 269488 336048
rect 269540 336036 269546 336048
rect 273088 336036 273116 336076
rect 273257 336073 273269 336107
rect 273303 336104 273315 336107
rect 277949 336107 278007 336113
rect 277949 336104 277961 336107
rect 273303 336076 277961 336104
rect 273303 336073 273315 336076
rect 273257 336067 273315 336073
rect 277949 336073 277961 336076
rect 277995 336073 278007 336107
rect 277949 336067 278007 336073
rect 278225 336107 278283 336113
rect 278225 336073 278237 336107
rect 278271 336104 278283 336107
rect 279418 336104 279424 336116
rect 278271 336076 279424 336104
rect 278271 336073 278283 336076
rect 278225 336067 278283 336073
rect 279418 336064 279424 336076
rect 279476 336064 279482 336116
rect 279513 336107 279571 336113
rect 279513 336073 279525 336107
rect 279559 336104 279571 336107
rect 404998 336104 405004 336116
rect 279559 336076 405004 336104
rect 279559 336073 279571 336076
rect 279513 336067 279571 336073
rect 404998 336064 405004 336076
rect 405056 336064 405062 336116
rect 273809 336039 273867 336045
rect 269540 336008 273024 336036
rect 273088 336008 273254 336036
rect 269540 335996 269546 336008
rect 263413 335971 263471 335977
rect 263413 335968 263425 335971
rect 262876 335940 263425 335968
rect 263413 335937 263425 335940
rect 263459 335937 263471 335971
rect 263413 335931 263471 335937
rect 268197 335971 268255 335977
rect 268197 335937 268209 335971
rect 268243 335968 268255 335971
rect 268243 335940 271920 335968
rect 268243 335937 268255 335940
rect 268197 335931 268255 335937
rect 262784 335872 263364 335900
rect 171778 335792 171784 335844
rect 171836 335832 171842 335844
rect 238941 335835 238999 335841
rect 238941 335832 238953 335835
rect 171836 335804 238953 335832
rect 171836 335792 171842 335804
rect 238941 335801 238953 335804
rect 238987 335801 238999 335835
rect 238941 335795 238999 335801
rect 239401 335835 239459 335841
rect 239401 335801 239413 335835
rect 239447 335832 239459 335835
rect 242345 335835 242403 335841
rect 242345 335832 242357 335835
rect 239447 335804 242357 335832
rect 239447 335801 239459 335804
rect 239401 335795 239459 335801
rect 242345 335801 242357 335804
rect 242391 335801 242403 335835
rect 242345 335795 242403 335801
rect 244737 335835 244795 335841
rect 244737 335801 244749 335835
rect 244783 335832 244795 335835
rect 248138 335832 248144 335844
rect 244783 335804 248144 335832
rect 244783 335801 244795 335804
rect 244737 335795 244795 335801
rect 248138 335792 248144 335804
rect 248196 335792 248202 335844
rect 256142 335792 256148 335844
rect 256200 335832 256206 335844
rect 258718 335832 258724 335844
rect 256200 335804 258724 335832
rect 256200 335792 256206 335804
rect 258718 335792 258724 335804
rect 258776 335792 258782 335844
rect 262950 335792 262956 335844
rect 263008 335832 263014 335844
rect 263226 335832 263232 335844
rect 263008 335804 263232 335832
rect 263008 335792 263014 335804
rect 263226 335792 263232 335804
rect 263284 335792 263290 335844
rect 263336 335832 263364 335872
rect 264974 335860 264980 335912
rect 265032 335900 265038 335912
rect 268470 335900 268476 335912
rect 265032 335872 268476 335900
rect 265032 335860 265038 335872
rect 268470 335860 268476 335872
rect 268528 335860 268534 335912
rect 269666 335860 269672 335912
rect 269724 335900 269730 335912
rect 270310 335900 270316 335912
rect 269724 335872 270316 335900
rect 269724 335860 269730 335872
rect 270310 335860 270316 335872
rect 270368 335860 270374 335912
rect 271892 335900 271920 335940
rect 271966 335928 271972 335980
rect 272024 335968 272030 335980
rect 272518 335968 272524 335980
rect 272024 335940 272524 335968
rect 272024 335928 272030 335940
rect 272518 335928 272524 335940
rect 272576 335928 272582 335980
rect 272996 335968 273024 336008
rect 273073 335971 273131 335977
rect 273073 335968 273085 335971
rect 272996 335940 273085 335968
rect 273073 335937 273085 335940
rect 273119 335937 273131 335971
rect 273226 335968 273254 336008
rect 273809 336005 273821 336039
rect 273855 336036 273867 336039
rect 407758 336036 407764 336048
rect 273855 336008 407764 336036
rect 273855 336005 273867 336008
rect 273809 335999 273867 336005
rect 407758 335996 407764 336008
rect 407816 335996 407822 336048
rect 337378 335968 337384 335980
rect 273226 335940 337384 335968
rect 273073 335931 273131 335937
rect 337378 335928 337384 335940
rect 337436 335928 337442 335980
rect 273165 335903 273223 335909
rect 273165 335900 273177 335903
rect 271892 335872 273177 335900
rect 273165 335869 273177 335872
rect 273211 335869 273223 335903
rect 273165 335863 273223 335869
rect 274726 335860 274732 335912
rect 274784 335900 274790 335912
rect 275922 335900 275928 335912
rect 274784 335872 275928 335900
rect 274784 335860 274790 335872
rect 275922 335860 275928 335872
rect 275980 335860 275986 335912
rect 277394 335860 277400 335912
rect 277452 335900 277458 335912
rect 278498 335900 278504 335912
rect 277452 335872 278504 335900
rect 277452 335860 277458 335872
rect 278498 335860 278504 335872
rect 278556 335860 278562 335912
rect 278685 335903 278743 335909
rect 278685 335869 278697 335903
rect 278731 335900 278743 335903
rect 279513 335903 279571 335909
rect 279513 335900 279525 335903
rect 278731 335872 279525 335900
rect 278731 335869 278743 335872
rect 278685 335863 278743 335869
rect 279513 335869 279525 335872
rect 279559 335869 279571 335903
rect 279513 335863 279571 335869
rect 280338 335860 280344 335912
rect 280396 335900 280402 335912
rect 281813 335903 281871 335909
rect 281813 335900 281825 335903
rect 280396 335872 281825 335900
rect 280396 335860 280402 335872
rect 281813 335869 281825 335872
rect 281859 335869 281871 335903
rect 281813 335863 281871 335869
rect 283282 335860 283288 335912
rect 283340 335900 283346 335912
rect 284389 335903 284447 335909
rect 283340 335872 284340 335900
rect 283340 335860 283346 335872
rect 264514 335832 264520 335844
rect 263336 335804 264520 335832
rect 264514 335792 264520 335804
rect 264572 335792 264578 335844
rect 269850 335832 269856 335844
rect 266740 335804 269856 335832
rect 178678 335724 178684 335776
rect 178736 335764 178742 335776
rect 239030 335764 239036 335776
rect 178736 335736 239036 335764
rect 178736 335724 178742 335736
rect 239030 335724 239036 335736
rect 239088 335724 239094 335776
rect 239125 335767 239183 335773
rect 239125 335733 239137 335767
rect 239171 335764 239183 335767
rect 243725 335767 243783 335773
rect 243725 335764 243737 335767
rect 239171 335736 243737 335764
rect 239171 335733 239183 335736
rect 239125 335727 239183 335733
rect 243725 335733 243737 335736
rect 243771 335733 243783 335767
rect 243725 335727 243783 335733
rect 243817 335767 243875 335773
rect 243817 335733 243829 335767
rect 243863 335764 243875 335767
rect 245286 335764 245292 335776
rect 243863 335736 245292 335764
rect 243863 335733 243875 335736
rect 243817 335727 243875 335733
rect 245286 335724 245292 335736
rect 245344 335724 245350 335776
rect 257246 335724 257252 335776
rect 257304 335764 257310 335776
rect 257890 335764 257896 335776
rect 257304 335736 257896 335764
rect 257304 335724 257310 335736
rect 257890 335724 257896 335736
rect 257948 335724 257954 335776
rect 263505 335767 263563 335773
rect 263505 335733 263517 335767
rect 263551 335764 263563 335767
rect 266740 335764 266768 335804
rect 269850 335792 269856 335804
rect 269908 335792 269914 335844
rect 273898 335792 273904 335844
rect 273956 335832 273962 335844
rect 274174 335832 274180 335844
rect 273956 335804 274180 335832
rect 273956 335792 273962 335804
rect 274174 335792 274180 335804
rect 274232 335792 274238 335844
rect 274453 335835 274511 335841
rect 274453 335801 274465 335835
rect 274499 335832 274511 335835
rect 278777 335835 278835 335841
rect 274499 335804 278636 335832
rect 274499 335801 274511 335804
rect 274453 335795 274511 335801
rect 263551 335736 266768 335764
rect 268013 335767 268071 335773
rect 263551 335733 263563 335736
rect 263505 335727 263563 335733
rect 268013 335733 268025 335767
rect 268059 335764 268071 335767
rect 269485 335767 269543 335773
rect 268059 335736 268332 335764
rect 268059 335733 268071 335736
rect 268013 335727 268071 335733
rect 180058 335656 180064 335708
rect 180116 335696 180122 335708
rect 239217 335699 239275 335705
rect 239217 335696 239229 335699
rect 180116 335668 239229 335696
rect 180116 335656 180122 335668
rect 239217 335665 239229 335668
rect 239263 335665 239275 335699
rect 239217 335659 239275 335665
rect 239309 335699 239367 335705
rect 239309 335665 239321 335699
rect 239355 335696 239367 335699
rect 244918 335696 244924 335708
rect 239355 335668 244924 335696
rect 239355 335665 239367 335668
rect 239309 335659 239367 335665
rect 244918 335656 244924 335668
rect 244976 335656 244982 335708
rect 245565 335699 245623 335705
rect 245565 335665 245577 335699
rect 245611 335696 245623 335699
rect 251266 335696 251272 335708
rect 245611 335668 251272 335696
rect 245611 335665 245623 335668
rect 245565 335659 245623 335665
rect 251266 335656 251272 335668
rect 251324 335656 251330 335708
rect 259546 335656 259552 335708
rect 259604 335696 259610 335708
rect 261110 335696 261116 335708
rect 259604 335668 261116 335696
rect 259604 335656 259610 335668
rect 261110 335656 261116 335668
rect 261168 335656 261174 335708
rect 268304 335696 268332 335736
rect 269485 335733 269497 335767
rect 269531 335764 269543 335767
rect 278501 335767 278559 335773
rect 278501 335764 278513 335767
rect 269531 335736 278513 335764
rect 269531 335733 269543 335736
rect 269485 335727 269543 335733
rect 278501 335733 278513 335736
rect 278547 335733 278559 335767
rect 278608 335764 278636 335804
rect 278777 335801 278789 335835
rect 278823 335832 278835 335835
rect 282733 335835 282791 335841
rect 282733 335832 282745 335835
rect 278823 335804 282745 335832
rect 278823 335801 278835 335804
rect 278777 335795 278835 335801
rect 282733 335801 282745 335804
rect 282779 335801 282791 335835
rect 282733 335795 282791 335801
rect 283190 335792 283196 335844
rect 283248 335832 283254 335844
rect 283466 335832 283472 335844
rect 283248 335804 283472 335832
rect 283248 335792 283254 335804
rect 283466 335792 283472 335804
rect 283524 335792 283530 335844
rect 284312 335832 284340 335872
rect 284389 335869 284401 335903
rect 284435 335900 284447 335903
rect 344554 335900 344560 335912
rect 284435 335872 344560 335900
rect 284435 335869 284447 335872
rect 284389 335863 284447 335869
rect 344554 335860 344560 335872
rect 344612 335860 344618 335912
rect 344462 335832 344468 335844
rect 284312 335804 344468 335832
rect 344462 335792 344468 335804
rect 344520 335792 344526 335844
rect 280798 335764 280804 335776
rect 278608 335736 280804 335764
rect 278501 335727 278559 335733
rect 280798 335724 280804 335736
rect 280856 335724 280862 335776
rect 281994 335724 282000 335776
rect 282052 335764 282058 335776
rect 282822 335764 282828 335776
rect 282052 335736 282828 335764
rect 282052 335724 282058 335736
rect 282822 335724 282828 335736
rect 282880 335724 282886 335776
rect 285217 335767 285275 335773
rect 285217 335733 285229 335767
rect 285263 335764 285275 335767
rect 344370 335764 344376 335776
rect 285263 335736 344376 335764
rect 285263 335733 285275 335736
rect 285217 335727 285275 335733
rect 344370 335724 344376 335736
rect 344428 335724 344434 335776
rect 316678 335696 316684 335708
rect 268304 335668 316684 335696
rect 316678 335656 316684 335668
rect 316736 335656 316742 335708
rect 231118 335588 231124 335640
rect 231176 335628 231182 335640
rect 236822 335628 236828 335640
rect 231176 335600 236828 335628
rect 231176 335588 231182 335600
rect 236822 335588 236828 335600
rect 236880 335588 236886 335640
rect 237193 335631 237251 335637
rect 237193 335597 237205 335631
rect 237239 335628 237251 335631
rect 243814 335628 243820 335640
rect 237239 335600 243820 335628
rect 237239 335597 237251 335600
rect 237193 335591 237251 335597
rect 243814 335588 243820 335600
rect 243872 335588 243878 335640
rect 244461 335631 244519 335637
rect 244461 335628 244473 335631
rect 243924 335600 244473 335628
rect 234801 335563 234859 335569
rect 234801 335529 234813 335563
rect 234847 335560 234859 335563
rect 240410 335560 240416 335572
rect 234847 335532 240416 335560
rect 234847 335529 234859 335532
rect 234801 335523 234859 335529
rect 240410 335520 240416 335532
rect 240468 335520 240474 335572
rect 242345 335563 242403 335569
rect 242345 335529 242357 335563
rect 242391 335560 242403 335563
rect 243924 335560 243952 335600
rect 244461 335597 244473 335600
rect 244507 335597 244519 335631
rect 257890 335628 257896 335640
rect 257851 335600 257896 335628
rect 244461 335591 244519 335597
rect 257890 335588 257896 335600
rect 257948 335588 257954 335640
rect 260742 335588 260748 335640
rect 260800 335628 260806 335640
rect 260800 335600 262168 335628
rect 260800 335588 260806 335600
rect 247218 335560 247224 335572
rect 242391 335532 243952 335560
rect 244016 335532 247224 335560
rect 242391 335529 242403 335532
rect 242345 335523 242403 335529
rect 232866 335452 232872 335504
rect 232924 335492 232930 335504
rect 232924 335464 236408 335492
rect 232924 335452 232930 335464
rect 231210 335384 231216 335436
rect 231268 335424 231274 335436
rect 234801 335427 234859 335433
rect 234801 335424 234813 335427
rect 231268 335396 234813 335424
rect 231268 335384 231274 335396
rect 234801 335393 234813 335396
rect 234847 335393 234859 335427
rect 234801 335387 234859 335393
rect 234982 335384 234988 335436
rect 235040 335424 235046 335436
rect 235905 335427 235963 335433
rect 235905 335424 235917 335427
rect 235040 335396 235917 335424
rect 235040 335384 235046 335396
rect 235905 335393 235917 335396
rect 235951 335393 235963 335427
rect 236380 335424 236408 335464
rect 237926 335452 237932 335504
rect 237984 335492 237990 335504
rect 241609 335495 241667 335501
rect 241609 335492 241621 335495
rect 237984 335464 241621 335492
rect 237984 335452 237990 335464
rect 241609 335461 241621 335464
rect 241655 335461 241667 335495
rect 241609 335455 241667 335461
rect 242158 335452 242164 335504
rect 242216 335492 242222 335504
rect 243354 335492 243360 335504
rect 242216 335464 243360 335492
rect 242216 335452 242222 335464
rect 243354 335452 243360 335464
rect 243412 335452 243418 335504
rect 242066 335424 242072 335436
rect 236380 335396 242072 335424
rect 235905 335387 235963 335393
rect 242066 335384 242072 335396
rect 242124 335384 242130 335436
rect 242250 335384 242256 335436
rect 242308 335424 242314 335436
rect 244016 335424 244044 335532
rect 247218 335520 247224 335532
rect 247276 335520 247282 335572
rect 244182 335452 244188 335504
rect 244240 335492 244246 335504
rect 245565 335495 245623 335501
rect 245565 335492 245577 335495
rect 244240 335464 245577 335492
rect 244240 335452 244246 335464
rect 245565 335461 245577 335464
rect 245611 335461 245623 335495
rect 245565 335455 245623 335461
rect 260558 335452 260564 335504
rect 260616 335492 260622 335504
rect 260742 335492 260748 335504
rect 260616 335464 260748 335492
rect 260616 335452 260622 335464
rect 260742 335452 260748 335464
rect 260800 335452 260806 335504
rect 242308 335396 244044 335424
rect 242308 335384 242314 335396
rect 244458 335384 244464 335436
rect 244516 335424 244522 335436
rect 244829 335427 244887 335433
rect 244829 335424 244841 335427
rect 244516 335396 244841 335424
rect 244516 335384 244522 335396
rect 244829 335393 244841 335396
rect 244875 335393 244887 335427
rect 244829 335387 244887 335393
rect 6822 335316 6828 335368
rect 6880 335356 6886 335368
rect 234709 335359 234767 335365
rect 234709 335356 234721 335359
rect 6880 335328 234721 335356
rect 6880 335316 6886 335328
rect 234709 335325 234721 335328
rect 234755 335325 234767 335359
rect 234709 335319 234767 335325
rect 238018 335316 238024 335368
rect 238076 335356 238082 335368
rect 239861 335359 239919 335365
rect 239861 335356 239873 335359
rect 238076 335328 239873 335356
rect 238076 335316 238082 335328
rect 239861 335325 239873 335328
rect 239907 335325 239919 335359
rect 239861 335319 239919 335325
rect 241238 335316 241244 335368
rect 241296 335356 241302 335368
rect 255682 335356 255688 335368
rect 241296 335328 255688 335356
rect 241296 335316 241302 335328
rect 255682 335316 255688 335328
rect 255740 335316 255746 335368
rect 256878 335316 256884 335368
rect 256936 335356 256942 335368
rect 257338 335356 257344 335368
rect 256936 335328 257344 335356
rect 256936 335316 256942 335328
rect 257338 335316 257344 335328
rect 257396 335316 257402 335368
rect 260374 335316 260380 335368
rect 260432 335356 260438 335368
rect 260558 335356 260564 335368
rect 260432 335328 260564 335356
rect 260432 335316 260438 335328
rect 260558 335316 260564 335328
rect 260616 335316 260622 335368
rect 261018 335316 261024 335368
rect 261076 335356 261082 335368
rect 261478 335356 261484 335368
rect 261076 335328 261484 335356
rect 261076 335316 261082 335328
rect 261478 335316 261484 335328
rect 261536 335316 261542 335368
rect 261754 335316 261760 335368
rect 261812 335356 261818 335368
rect 261938 335356 261944 335368
rect 261812 335328 261944 335356
rect 261812 335316 261818 335328
rect 261938 335316 261944 335328
rect 261996 335316 262002 335368
rect 262140 335356 262168 335600
rect 262398 335588 262404 335640
rect 262456 335628 262462 335640
rect 263134 335628 263140 335640
rect 262456 335600 263140 335628
rect 262456 335588 262462 335600
rect 263134 335588 263140 335600
rect 263192 335588 263198 335640
rect 263229 335631 263287 335637
rect 263229 335597 263241 335631
rect 263275 335628 263287 335631
rect 268289 335631 268347 335637
rect 268289 335628 268301 335631
rect 263275 335600 268301 335628
rect 263275 335597 263287 335600
rect 263229 335591 263287 335597
rect 268289 335597 268301 335600
rect 268335 335597 268347 335631
rect 300210 335628 300216 335640
rect 268289 335591 268347 335597
rect 268396 335600 300216 335628
rect 262861 335563 262919 335569
rect 262861 335529 262873 335563
rect 262907 335560 262919 335563
rect 268396 335560 268424 335600
rect 300210 335588 300216 335600
rect 300268 335588 300274 335640
rect 262907 335532 268424 335560
rect 268841 335563 268899 335569
rect 262907 335529 262919 335532
rect 262861 335523 262919 335529
rect 268841 335529 268853 335563
rect 268887 335560 268899 335563
rect 271966 335560 271972 335572
rect 268887 335532 271972 335560
rect 268887 335529 268899 335532
rect 268841 335523 268899 335529
rect 271966 335520 271972 335532
rect 272024 335520 272030 335572
rect 273717 335563 273775 335569
rect 273717 335529 273729 335563
rect 273763 335560 273775 335563
rect 274450 335560 274456 335572
rect 273763 335532 274456 335560
rect 273763 335529 273775 335532
rect 273717 335523 273775 335529
rect 274450 335520 274456 335532
rect 274508 335520 274514 335572
rect 274818 335520 274824 335572
rect 274876 335560 274882 335572
rect 275462 335560 275468 335572
rect 274876 335532 275468 335560
rect 274876 335520 274882 335532
rect 275462 335520 275468 335532
rect 275520 335520 275526 335572
rect 277946 335520 277952 335572
rect 278004 335560 278010 335572
rect 278498 335560 278504 335572
rect 278004 335532 278504 335560
rect 278004 335520 278010 335532
rect 278498 335520 278504 335532
rect 278556 335520 278562 335572
rect 281810 335520 281816 335572
rect 281868 335560 281874 335572
rect 282546 335560 282552 335572
rect 281868 335532 282552 335560
rect 281868 335520 281874 335532
rect 282546 335520 282552 335532
rect 282604 335520 282610 335572
rect 283466 335560 283472 335572
rect 283427 335532 283472 335560
rect 283466 335520 283472 335532
rect 283524 335520 283530 335572
rect 283742 335520 283748 335572
rect 283800 335560 283806 335572
rect 283800 335532 284248 335560
rect 283800 335520 283806 335532
rect 268102 335452 268108 335504
rect 268160 335492 268166 335504
rect 268289 335495 268347 335501
rect 268289 335492 268301 335495
rect 268160 335464 268301 335492
rect 268160 335452 268166 335464
rect 268289 335461 268301 335464
rect 268335 335461 268347 335495
rect 268289 335455 268347 335461
rect 268473 335495 268531 335501
rect 268473 335461 268485 335495
rect 268519 335492 268531 335495
rect 269758 335492 269764 335504
rect 268519 335464 269764 335492
rect 268519 335461 268531 335464
rect 268473 335455 268531 335461
rect 269758 335452 269764 335464
rect 269816 335452 269822 335504
rect 272058 335452 272064 335504
rect 272116 335492 272122 335504
rect 272794 335492 272800 335504
rect 272116 335464 272800 335492
rect 272116 335452 272122 335464
rect 272794 335452 272800 335464
rect 272852 335452 272858 335504
rect 273073 335495 273131 335501
rect 273073 335461 273085 335495
rect 273119 335492 273131 335495
rect 273809 335495 273867 335501
rect 273809 335492 273821 335495
rect 273119 335464 273821 335492
rect 273119 335461 273131 335464
rect 273073 335455 273131 335461
rect 273809 335461 273821 335464
rect 273855 335461 273867 335495
rect 273809 335455 273867 335461
rect 273898 335452 273904 335504
rect 273956 335492 273962 335504
rect 274542 335492 274548 335504
rect 273956 335464 274548 335492
rect 273956 335452 273962 335464
rect 274542 335452 274548 335464
rect 274600 335452 274606 335504
rect 275741 335495 275799 335501
rect 275741 335461 275753 335495
rect 275787 335492 275799 335495
rect 278317 335495 278375 335501
rect 278317 335492 278329 335495
rect 275787 335464 278329 335492
rect 275787 335461 275799 335464
rect 275741 335455 275799 335461
rect 278317 335461 278329 335464
rect 278363 335461 278375 335495
rect 281350 335492 281356 335504
rect 281311 335464 281356 335492
rect 278317 335455 278375 335461
rect 281350 335452 281356 335464
rect 281408 335452 281414 335504
rect 281994 335492 282000 335504
rect 281955 335464 282000 335492
rect 281994 335452 282000 335464
rect 282052 335452 282058 335504
rect 282086 335452 282092 335504
rect 282144 335492 282150 335504
rect 282638 335492 282644 335504
rect 282144 335464 282644 335492
rect 282144 335452 282150 335464
rect 282638 335452 282644 335464
rect 282696 335452 282702 335504
rect 262858 335384 262864 335436
rect 262916 335424 262922 335436
rect 263318 335424 263324 335436
rect 262916 335396 263324 335424
rect 262916 335384 262922 335396
rect 263318 335384 263324 335396
rect 263376 335384 263382 335436
rect 263778 335384 263784 335436
rect 263836 335424 263842 335436
rect 268749 335427 268807 335433
rect 268749 335424 268761 335427
rect 263836 335396 268761 335424
rect 263836 335384 263842 335396
rect 268749 335393 268761 335396
rect 268795 335393 268807 335427
rect 268749 335387 268807 335393
rect 270678 335384 270684 335436
rect 270736 335424 270742 335436
rect 271782 335424 271788 335436
rect 270736 335396 271788 335424
rect 270736 335384 270742 335396
rect 271782 335384 271788 335396
rect 271840 335384 271846 335436
rect 272981 335427 273039 335433
rect 272981 335393 272993 335427
rect 273027 335424 273039 335427
rect 273027 335396 278084 335424
rect 273027 335393 273039 335396
rect 272981 335387 273039 335393
rect 262140 335328 262444 335356
rect 201402 335248 201408 335300
rect 201460 335288 201466 335300
rect 244182 335288 244188 335300
rect 201460 335260 244188 335288
rect 201460 335248 201466 335260
rect 244182 335248 244188 335260
rect 244240 335248 244246 335300
rect 245010 335248 245016 335300
rect 245068 335288 245074 335300
rect 254210 335288 254216 335300
rect 245068 335260 254216 335288
rect 245068 335248 245074 335260
rect 254210 335248 254216 335260
rect 254268 335248 254274 335300
rect 262416 335288 262444 335328
rect 263870 335316 263876 335368
rect 263928 335356 263934 335368
rect 264330 335356 264336 335368
rect 263928 335328 264336 335356
rect 263928 335316 263934 335328
rect 264330 335316 264336 335328
rect 264388 335316 264394 335368
rect 267734 335316 267740 335368
rect 267792 335356 267798 335368
rect 267918 335356 267924 335368
rect 267792 335328 267924 335356
rect 267792 335316 267798 335328
rect 267918 335316 267924 335328
rect 267976 335316 267982 335368
rect 269942 335316 269948 335368
rect 270000 335356 270006 335368
rect 270402 335356 270408 335368
rect 270000 335328 270408 335356
rect 270000 335316 270006 335328
rect 270402 335316 270408 335328
rect 270460 335316 270466 335368
rect 274726 335316 274732 335368
rect 274784 335356 274790 335368
rect 274910 335356 274916 335368
rect 274784 335328 274916 335356
rect 274784 335316 274790 335328
rect 274910 335316 274916 335328
rect 274968 335316 274974 335368
rect 275462 335356 275468 335368
rect 275423 335328 275468 335356
rect 275462 335316 275468 335328
rect 275520 335316 275526 335368
rect 275554 335316 275560 335368
rect 275612 335356 275618 335368
rect 275738 335356 275744 335368
rect 275612 335328 275744 335356
rect 275612 335316 275618 335328
rect 275738 335316 275744 335328
rect 275796 335316 275802 335368
rect 277394 335316 277400 335368
rect 277452 335356 277458 335368
rect 277762 335356 277768 335368
rect 277452 335328 277768 335356
rect 277452 335316 277458 335328
rect 277762 335316 277768 335328
rect 277820 335316 277826 335368
rect 277857 335359 277915 335365
rect 277857 335325 277869 335359
rect 277903 335356 277915 335359
rect 277946 335356 277952 335368
rect 277903 335328 277952 335356
rect 277903 335325 277915 335328
rect 277857 335319 277915 335325
rect 277946 335316 277952 335328
rect 278004 335316 278010 335368
rect 278056 335356 278084 335396
rect 278222 335384 278228 335436
rect 278280 335424 278286 335436
rect 278406 335424 278412 335436
rect 278280 335396 278412 335424
rect 278280 335384 278286 335396
rect 278406 335384 278412 335396
rect 278464 335384 278470 335436
rect 278501 335427 278559 335433
rect 278501 335393 278513 335427
rect 278547 335424 278559 335427
rect 278547 335396 283512 335424
rect 278547 335393 278559 335396
rect 278501 335387 278559 335393
rect 283484 335356 283512 335396
rect 283558 335384 283564 335436
rect 283616 335424 283622 335436
rect 284018 335424 284024 335436
rect 283616 335396 284024 335424
rect 283616 335384 283622 335396
rect 284018 335384 284024 335396
rect 284076 335384 284082 335436
rect 278056 335328 283420 335356
rect 283484 335328 283696 335356
rect 262582 335288 262588 335300
rect 262416 335260 262588 335288
rect 262582 335248 262588 335260
rect 262640 335248 262646 335300
rect 268289 335291 268347 335297
rect 268289 335257 268301 335291
rect 268335 335288 268347 335291
rect 268746 335288 268752 335300
rect 268335 335260 268752 335288
rect 268335 335257 268347 335260
rect 268289 335251 268347 335257
rect 268746 335248 268752 335260
rect 268804 335248 268810 335300
rect 282270 335288 282276 335300
rect 276354 335260 282276 335288
rect 208302 335180 208308 335232
rect 208360 335220 208366 335232
rect 251453 335223 251511 335229
rect 251453 335220 251465 335223
rect 208360 335192 251465 335220
rect 208360 335180 208366 335192
rect 251453 335189 251465 335192
rect 251499 335189 251511 335223
rect 251453 335183 251511 335189
rect 258905 335223 258963 335229
rect 258905 335189 258917 335223
rect 258951 335220 258963 335223
rect 276354 335220 276382 335260
rect 282270 335248 282276 335260
rect 282328 335248 282334 335300
rect 282546 335288 282552 335300
rect 282507 335260 282552 335288
rect 282546 335248 282552 335260
rect 282604 335248 282610 335300
rect 282733 335291 282791 335297
rect 282733 335257 282745 335291
rect 282779 335288 282791 335291
rect 282779 335260 283190 335288
rect 282779 335257 282791 335260
rect 282733 335251 282791 335257
rect 282638 335220 282644 335232
rect 258951 335192 276382 335220
rect 276446 335192 282644 335220
rect 258951 335189 258963 335192
rect 258905 335183 258963 335189
rect 197262 335112 197268 335164
rect 197320 335152 197326 335164
rect 250990 335152 250996 335164
rect 197320 335124 250996 335152
rect 197320 335112 197326 335124
rect 250990 335112 250996 335124
rect 251048 335112 251054 335164
rect 276446 335152 276474 335192
rect 282638 335180 282644 335192
rect 282696 335180 282702 335232
rect 282917 335155 282975 335161
rect 282917 335152 282929 335155
rect 268396 335124 276474 335152
rect 276538 335124 282929 335152
rect 194502 335044 194508 335096
rect 194560 335084 194566 335096
rect 250533 335087 250591 335093
rect 250533 335084 250545 335087
rect 194560 335056 250545 335084
rect 194560 335044 194566 335056
rect 250533 335053 250545 335056
rect 250579 335053 250591 335087
rect 250533 335047 250591 335053
rect 251266 335044 251272 335096
rect 251324 335084 251330 335096
rect 255130 335084 255136 335096
rect 251324 335056 255136 335084
rect 251324 335044 251330 335056
rect 255130 335044 255136 335056
rect 255188 335044 255194 335096
rect 261754 335084 261760 335096
rect 261715 335056 261760 335084
rect 261754 335044 261760 335056
rect 261812 335044 261818 335096
rect 190362 334976 190368 335028
rect 190420 335016 190426 335028
rect 250438 335016 250444 335028
rect 190420 334988 250444 335016
rect 190420 334976 190426 334988
rect 250438 334976 250444 334988
rect 250496 334976 250502 335028
rect 183462 334908 183468 334960
rect 183520 334948 183526 334960
rect 242897 334951 242955 334957
rect 242897 334948 242909 334951
rect 183520 334920 242909 334948
rect 183520 334908 183526 334920
rect 242897 334917 242909 334920
rect 242943 334917 242955 334951
rect 242897 334911 242955 334917
rect 243262 334908 243268 334960
rect 243320 334948 243326 334960
rect 243998 334948 244004 334960
rect 243320 334920 244004 334948
rect 243320 334908 243326 334920
rect 243998 334908 244004 334920
rect 244056 334908 244062 334960
rect 245470 334948 245476 334960
rect 245431 334920 245476 334948
rect 245470 334908 245476 334920
rect 245528 334908 245534 334960
rect 186222 334840 186228 334892
rect 186280 334880 186286 334892
rect 250073 334883 250131 334889
rect 250073 334880 250085 334883
rect 186280 334852 250085 334880
rect 186280 334840 186286 334852
rect 250073 334849 250085 334852
rect 250119 334849 250131 334883
rect 250073 334843 250131 334849
rect 252738 334840 252744 334892
rect 252796 334880 252802 334892
rect 253290 334880 253296 334892
rect 252796 334852 253296 334880
rect 252796 334840 252802 334852
rect 253290 334840 253296 334852
rect 253348 334840 253354 334892
rect 258353 334883 258411 334889
rect 258353 334849 258365 334883
rect 258399 334880 258411 334883
rect 268396 334880 268424 335124
rect 276538 335084 276566 335124
rect 282917 335121 282929 335124
rect 282963 335121 282975 335155
rect 283162 335152 283190 335260
rect 283392 335220 283420 335328
rect 283668 335288 283696 335328
rect 284110 335316 284116 335368
rect 284168 335356 284174 335368
rect 284220 335356 284248 335532
rect 284294 335452 284300 335504
rect 284352 335492 284358 335504
rect 285398 335492 285404 335504
rect 284352 335464 285404 335492
rect 284352 335452 284358 335464
rect 285398 335452 285404 335464
rect 285456 335452 285462 335504
rect 284570 335384 284576 335436
rect 284628 335424 284634 335436
rect 285306 335424 285312 335436
rect 284628 335396 285312 335424
rect 284628 335384 284634 335396
rect 285306 335384 285312 335396
rect 285364 335384 285370 335436
rect 284168 335328 284248 335356
rect 284168 335316 284174 335328
rect 284662 335316 284668 335368
rect 284720 335356 284726 335368
rect 284846 335356 284852 335368
rect 284720 335328 284852 335356
rect 284720 335316 284726 335328
rect 284846 335316 284852 335328
rect 284904 335316 284910 335368
rect 285030 335288 285036 335300
rect 283668 335260 285036 335288
rect 285030 335248 285036 335260
rect 285088 335248 285094 335300
rect 285122 335220 285128 335232
rect 283392 335192 285128 335220
rect 285122 335180 285128 335192
rect 285180 335180 285186 335232
rect 285217 335223 285275 335229
rect 285217 335189 285229 335223
rect 285263 335220 285275 335223
rect 288434 335220 288440 335232
rect 285263 335192 288440 335220
rect 285263 335189 285275 335192
rect 285217 335183 285275 335189
rect 288434 335180 288440 335192
rect 288492 335180 288498 335232
rect 286410 335152 286416 335164
rect 283162 335124 286416 335152
rect 282917 335115 282975 335121
rect 286410 335112 286416 335124
rect 286468 335112 286474 335164
rect 258399 334852 268424 334880
rect 268488 335056 276566 335084
rect 277029 335087 277087 335093
rect 258399 334849 258411 334852
rect 258353 334843 258411 334849
rect 179322 334772 179328 334824
rect 179380 334812 179386 334824
rect 249518 334812 249524 334824
rect 179380 334784 249524 334812
rect 179380 334772 179386 334784
rect 249518 334772 249524 334784
rect 249576 334772 249582 334824
rect 258810 334772 258816 334824
rect 258868 334812 258874 334824
rect 268488 334812 268516 335056
rect 277029 335053 277041 335087
rect 277075 335084 277087 335087
rect 283006 335084 283012 335096
rect 277075 335056 283012 335084
rect 277075 335053 277087 335056
rect 277029 335047 277087 335053
rect 283006 335044 283012 335056
rect 283064 335044 283070 335096
rect 283101 335087 283159 335093
rect 283101 335053 283113 335087
rect 283147 335084 283159 335087
rect 289354 335084 289360 335096
rect 283147 335056 289360 335084
rect 283147 335053 283159 335056
rect 283101 335047 283159 335053
rect 289354 335044 289360 335056
rect 289412 335044 289418 335096
rect 273714 335016 273720 335028
rect 273675 334988 273720 335016
rect 273714 334976 273720 334988
rect 273772 334976 273778 335028
rect 276293 335019 276351 335025
rect 276293 334985 276305 335019
rect 276339 335016 276351 335019
rect 316034 335016 316040 335028
rect 276339 334988 316040 335016
rect 276339 334985 276351 334988
rect 276293 334979 276351 334985
rect 316034 334976 316040 334988
rect 316092 334976 316098 335028
rect 268933 334951 268991 334957
rect 268933 334917 268945 334951
rect 268979 334948 268991 334951
rect 369854 334948 369860 334960
rect 268979 334920 369860 334948
rect 268979 334917 268991 334920
rect 268933 334911 268991 334917
rect 369854 334908 369860 334920
rect 369912 334908 369918 334960
rect 276753 334883 276811 334889
rect 276753 334849 276765 334883
rect 276799 334880 276811 334883
rect 277026 334880 277032 334892
rect 276799 334852 277032 334880
rect 276799 334849 276811 334852
rect 276753 334843 276811 334849
rect 277026 334840 277032 334852
rect 277084 334840 277090 334892
rect 277949 334883 278007 334889
rect 277949 334849 277961 334883
rect 277995 334880 278007 334883
rect 401594 334880 401600 334892
rect 277995 334852 401600 334880
rect 277995 334849 278007 334852
rect 277949 334843 278007 334849
rect 401594 334840 401600 334852
rect 401652 334840 401658 334892
rect 271782 334812 271788 334824
rect 258868 334784 268516 334812
rect 271743 334784 271788 334812
rect 258868 334772 258874 334784
rect 271782 334772 271788 334784
rect 271840 334772 271846 334824
rect 271966 334772 271972 334824
rect 272024 334812 272030 334824
rect 276293 334815 276351 334821
rect 276293 334812 276305 334815
rect 272024 334784 276305 334812
rect 272024 334772 272030 334784
rect 276293 334781 276305 334784
rect 276339 334781 276351 334815
rect 276293 334775 276351 334781
rect 278041 334815 278099 334821
rect 278041 334781 278053 334815
rect 278087 334812 278099 334815
rect 415486 334812 415492 334824
rect 278087 334784 415492 334812
rect 278087 334781 278099 334784
rect 278041 334775 278099 334781
rect 415486 334772 415492 334784
rect 415544 334772 415550 334824
rect 169662 334704 169668 334756
rect 169720 334744 169726 334756
rect 240226 334744 240232 334756
rect 169720 334716 240232 334744
rect 169720 334704 169726 334716
rect 240226 334704 240232 334716
rect 240284 334704 240290 334756
rect 240321 334747 240379 334753
rect 240321 334713 240333 334747
rect 240367 334744 240379 334747
rect 248322 334744 248328 334756
rect 240367 334716 248328 334744
rect 240367 334713 240379 334716
rect 240321 334707 240379 334713
rect 248322 334704 248328 334716
rect 248380 334704 248386 334756
rect 272518 334704 272524 334756
rect 272576 334744 272582 334756
rect 438118 334744 438124 334756
rect 272576 334716 438124 334744
rect 272576 334704 272582 334716
rect 438118 334704 438124 334716
rect 438176 334704 438182 334756
rect 176562 334636 176568 334688
rect 176620 334676 176626 334688
rect 248966 334676 248972 334688
rect 176620 334648 248972 334676
rect 176620 334636 176626 334648
rect 248966 334636 248972 334648
rect 249024 334636 249030 334688
rect 257617 334679 257675 334685
rect 257617 334645 257629 334679
rect 257663 334676 257675 334679
rect 260006 334676 260012 334688
rect 257663 334648 260012 334676
rect 257663 334645 257675 334648
rect 257617 334639 257675 334645
rect 260006 334636 260012 334648
rect 260064 334636 260070 334688
rect 265526 334636 265532 334688
rect 265584 334676 265590 334688
rect 373994 334676 374000 334688
rect 265584 334648 374000 334676
rect 265584 334636 265590 334648
rect 373994 334636 374000 334648
rect 374052 334636 374058 334688
rect 395338 334636 395344 334688
rect 395396 334676 395402 334688
rect 580718 334676 580724 334688
rect 395396 334648 580724 334676
rect 395396 334636 395402 334648
rect 580718 334636 580724 334648
rect 580776 334636 580782 334688
rect 165522 334568 165528 334620
rect 165580 334608 165586 334620
rect 234617 334611 234675 334617
rect 234617 334608 234629 334611
rect 165580 334580 234629 334608
rect 165580 334568 165586 334580
rect 234617 334577 234629 334580
rect 234663 334577 234675 334611
rect 234617 334571 234675 334577
rect 235629 334611 235687 334617
rect 235629 334577 235641 334611
rect 235675 334608 235687 334611
rect 238754 334608 238760 334620
rect 235675 334580 238760 334608
rect 235675 334577 235687 334580
rect 235629 334571 235687 334577
rect 238754 334568 238760 334580
rect 238812 334568 238818 334620
rect 239033 334611 239091 334617
rect 239033 334577 239045 334611
rect 239079 334608 239091 334611
rect 240321 334611 240379 334617
rect 240321 334608 240333 334611
rect 239079 334580 240333 334608
rect 239079 334577 239091 334580
rect 239033 334571 239091 334577
rect 240321 334577 240333 334580
rect 240367 334577 240379 334611
rect 240321 334571 240379 334577
rect 240410 334568 240416 334620
rect 240468 334608 240474 334620
rect 240468 334580 240513 334608
rect 240468 334568 240474 334580
rect 240870 334568 240876 334620
rect 240928 334608 240934 334620
rect 241238 334608 241244 334620
rect 240928 334580 241244 334608
rect 240928 334568 240934 334580
rect 241238 334568 241244 334580
rect 241296 334568 241302 334620
rect 243538 334568 243544 334620
rect 243596 334608 243602 334620
rect 243722 334608 243728 334620
rect 243596 334580 243728 334608
rect 243596 334568 243602 334580
rect 243722 334568 243728 334580
rect 243780 334568 243786 334620
rect 244642 334568 244648 334620
rect 244700 334608 244706 334620
rect 245194 334608 245200 334620
rect 244700 334580 245200 334608
rect 244700 334568 244706 334580
rect 245194 334568 245200 334580
rect 245252 334568 245258 334620
rect 251818 334568 251824 334620
rect 251876 334608 251882 334620
rect 252094 334608 252100 334620
rect 251876 334580 252100 334608
rect 251876 334568 251882 334580
rect 252094 334568 252100 334580
rect 252152 334568 252158 334620
rect 254302 334608 254308 334620
rect 254263 334580 254308 334608
rect 254302 334568 254308 334580
rect 254360 334568 254366 334620
rect 274634 334568 274640 334620
rect 274692 334608 274698 334620
rect 280982 334608 280988 334620
rect 274692 334580 280988 334608
rect 274692 334568 274698 334580
rect 280982 334568 280988 334580
rect 281040 334568 281046 334620
rect 281813 334611 281871 334617
rect 281813 334577 281825 334611
rect 281859 334608 281871 334611
rect 554774 334608 554780 334620
rect 281859 334580 554780 334608
rect 281859 334577 281871 334580
rect 281813 334571 281871 334577
rect 554774 334568 554780 334580
rect 554832 334568 554838 334620
rect 204162 334500 204168 334552
rect 204220 334540 204226 334552
rect 244458 334540 244464 334552
rect 204220 334512 244464 334540
rect 204220 334500 204226 334512
rect 244458 334500 244464 334512
rect 244516 334500 244522 334552
rect 265894 334500 265900 334552
rect 265952 334540 265958 334552
rect 268197 334543 268255 334549
rect 268197 334540 268209 334543
rect 265952 334512 268209 334540
rect 265952 334500 265958 334512
rect 268197 334509 268209 334512
rect 268243 334509 268255 334543
rect 268197 334503 268255 334509
rect 276290 334500 276296 334552
rect 276348 334540 276354 334552
rect 283101 334543 283159 334549
rect 283101 334540 283113 334543
rect 276348 334512 283113 334540
rect 276348 334500 276354 334512
rect 283101 334509 283113 334512
rect 283147 334509 283159 334543
rect 283101 334503 283159 334509
rect 283190 334500 283196 334552
rect 283248 334540 283254 334552
rect 286594 334540 286600 334552
rect 283248 334512 286600 334540
rect 283248 334500 283254 334512
rect 286594 334500 286600 334512
rect 286652 334500 286658 334552
rect 210970 334432 210976 334484
rect 211028 334472 211034 334484
rect 252186 334472 252192 334484
rect 211028 334444 252192 334472
rect 211028 334432 211034 334444
rect 252186 334432 252192 334444
rect 252244 334432 252250 334484
rect 277397 334475 277455 334481
rect 277397 334441 277409 334475
rect 277443 334472 277455 334475
rect 282733 334475 282791 334481
rect 277443 334444 282684 334472
rect 277443 334441 277455 334444
rect 277397 334435 277455 334441
rect 215202 334364 215208 334416
rect 215260 334404 215266 334416
rect 252465 334407 252523 334413
rect 252465 334404 252477 334407
rect 215260 334376 252477 334404
rect 215260 334364 215266 334376
rect 252465 334373 252477 334376
rect 252511 334373 252523 334407
rect 252465 334367 252523 334373
rect 272150 334364 272156 334416
rect 272208 334404 272214 334416
rect 272886 334404 272892 334416
rect 272208 334376 272892 334404
rect 272208 334364 272214 334376
rect 272886 334364 272892 334376
rect 272944 334364 272950 334416
rect 276934 334364 276940 334416
rect 276992 334404 276998 334416
rect 279973 334407 280031 334413
rect 276992 334376 278176 334404
rect 276992 334364 276998 334376
rect 222102 334296 222108 334348
rect 222160 334336 222166 334348
rect 253014 334336 253020 334348
rect 222160 334308 253020 334336
rect 222160 334296 222166 334308
rect 253014 334296 253020 334308
rect 253072 334296 253078 334348
rect 269025 334339 269083 334345
rect 269025 334305 269037 334339
rect 269071 334336 269083 334339
rect 278041 334339 278099 334345
rect 278041 334336 278053 334339
rect 269071 334308 278053 334336
rect 269071 334305 269083 334308
rect 269025 334299 269083 334305
rect 278041 334305 278053 334308
rect 278087 334305 278099 334339
rect 278148 334336 278176 334376
rect 279973 334373 279985 334407
rect 280019 334404 280031 334407
rect 282273 334407 282331 334413
rect 282273 334404 282285 334407
rect 280019 334376 282285 334404
rect 280019 334373 280031 334376
rect 279973 334367 280031 334373
rect 282273 334373 282285 334376
rect 282319 334373 282331 334407
rect 282656 334404 282684 334444
rect 282733 334441 282745 334475
rect 282779 334472 282791 334475
rect 287882 334472 287888 334484
rect 282779 334444 287888 334472
rect 282779 334441 282791 334444
rect 282733 334435 282791 334441
rect 287882 334432 287888 334444
rect 287940 334432 287946 334484
rect 283745 334407 283803 334413
rect 283745 334404 283757 334407
rect 282656 334376 283757 334404
rect 282273 334367 282331 334373
rect 283745 334373 283757 334376
rect 283791 334373 283803 334407
rect 289262 334404 289268 334416
rect 283745 334367 283803 334373
rect 283852 334376 289268 334404
rect 283852 334336 283880 334376
rect 289262 334364 289268 334376
rect 289320 334364 289326 334416
rect 289078 334336 289084 334348
rect 278148 334308 283880 334336
rect 283944 334308 289084 334336
rect 278041 334299 278099 334305
rect 226242 334228 226248 334280
rect 226300 334268 226306 334280
rect 253382 334268 253388 334280
rect 226300 334240 253388 334268
rect 226300 334228 226306 334240
rect 253382 334228 253388 334240
rect 253440 334228 253446 334280
rect 269666 334228 269672 334280
rect 269724 334268 269730 334280
rect 274913 334271 274971 334277
rect 269724 334240 273254 334268
rect 269724 334228 269730 334240
rect 229002 334160 229008 334212
rect 229060 334200 229066 334212
rect 253566 334200 253572 334212
rect 229060 334172 253572 334200
rect 229060 334160 229066 334172
rect 253566 334160 253572 334172
rect 253624 334160 253630 334212
rect 273226 334200 273254 334240
rect 274913 334237 274925 334271
rect 274959 334268 274971 334271
rect 275370 334268 275376 334280
rect 274959 334240 275376 334268
rect 274959 334237 274971 334240
rect 274913 334231 274971 334237
rect 275370 334228 275376 334240
rect 275428 334228 275434 334280
rect 276569 334271 276627 334277
rect 276569 334237 276581 334271
rect 276615 334268 276627 334271
rect 283944 334268 283972 334308
rect 289078 334296 289084 334308
rect 289136 334296 289142 334348
rect 276615 334240 283972 334268
rect 284021 334271 284079 334277
rect 276615 334237 276627 334240
rect 276569 334231 276627 334237
rect 284021 334237 284033 334271
rect 284067 334268 284079 334271
rect 289170 334268 289176 334280
rect 284067 334240 289176 334268
rect 284067 334237 284079 334240
rect 284021 334231 284079 334237
rect 289170 334228 289176 334240
rect 289228 334228 289234 334280
rect 282270 334200 282276 334212
rect 273226 334172 282276 334200
rect 282270 334160 282276 334172
rect 282328 334160 282334 334212
rect 282362 334160 282368 334212
rect 282420 334200 282426 334212
rect 282420 334172 284156 334200
rect 282420 334160 282426 334172
rect 219342 334092 219348 334144
rect 219400 334132 219406 334144
rect 234617 334135 234675 334141
rect 234617 334132 234629 334135
rect 219400 334104 234629 334132
rect 219400 334092 219406 334104
rect 234617 334101 234629 334104
rect 234663 334101 234675 334135
rect 234617 334095 234675 334101
rect 234709 334135 234767 334141
rect 234709 334101 234721 334135
rect 234755 334132 234767 334135
rect 239033 334135 239091 334141
rect 239033 334132 239045 334135
rect 234755 334104 239045 334132
rect 234755 334101 234767 334104
rect 234709 334095 234767 334101
rect 239033 334101 239045 334104
rect 239079 334101 239091 334135
rect 239033 334095 239091 334101
rect 239122 334092 239128 334144
rect 239180 334132 239186 334144
rect 240042 334132 240048 334144
rect 239180 334104 240048 334132
rect 239180 334092 239186 334104
rect 240042 334092 240048 334104
rect 240100 334092 240106 334144
rect 240686 334092 240692 334144
rect 240744 334132 240750 334144
rect 240962 334132 240968 334144
rect 240744 334104 240968 334132
rect 240744 334092 240750 334104
rect 240962 334092 240968 334104
rect 241020 334092 241026 334144
rect 242066 334092 242072 334144
rect 242124 334132 242130 334144
rect 242526 334132 242532 334144
rect 242124 334104 242532 334132
rect 242124 334092 242130 334104
rect 242526 334092 242532 334104
rect 242584 334092 242590 334144
rect 242989 334135 243047 334141
rect 242989 334101 243001 334135
rect 243035 334132 243047 334135
rect 243814 334132 243820 334144
rect 243035 334104 243820 334132
rect 243035 334101 243047 334104
rect 242989 334095 243047 334101
rect 243814 334092 243820 334104
rect 243872 334092 243878 334144
rect 245194 334132 245200 334144
rect 245155 334104 245200 334132
rect 245194 334092 245200 334104
rect 245252 334092 245258 334144
rect 272702 334092 272708 334144
rect 272760 334132 272766 334144
rect 272889 334135 272947 334141
rect 272889 334132 272901 334135
rect 272760 334104 272901 334132
rect 272760 334092 272766 334104
rect 272889 334101 272901 334104
rect 272935 334101 272947 334135
rect 272889 334095 272947 334101
rect 276014 334092 276020 334144
rect 276072 334132 276078 334144
rect 276937 334135 276995 334141
rect 276937 334132 276949 334135
rect 276072 334104 276949 334132
rect 276072 334092 276078 334104
rect 276937 334101 276949 334104
rect 276983 334101 276995 334135
rect 276937 334095 276995 334101
rect 278590 334092 278596 334144
rect 278648 334132 278654 334144
rect 284021 334135 284079 334141
rect 284021 334132 284033 334135
rect 278648 334104 284033 334132
rect 278648 334092 278654 334104
rect 284021 334101 284033 334104
rect 284067 334101 284079 334135
rect 284128 334132 284156 334172
rect 285582 334160 285588 334212
rect 285640 334200 285646 334212
rect 287974 334200 287980 334212
rect 285640 334172 287980 334200
rect 285640 334160 285646 334172
rect 287974 334160 287980 334172
rect 288032 334160 288038 334212
rect 287790 334132 287796 334144
rect 284128 334104 287796 334132
rect 284021 334095 284079 334101
rect 287790 334092 287796 334104
rect 287848 334092 287854 334144
rect 231394 334024 231400 334076
rect 231452 334064 231458 334076
rect 248874 334064 248880 334076
rect 231452 334036 248880 334064
rect 231452 334024 231458 334036
rect 248874 334024 248880 334036
rect 248932 334024 248938 334076
rect 250346 334024 250352 334076
rect 250404 334064 250410 334076
rect 254670 334064 254676 334076
rect 250404 334036 254676 334064
rect 250404 334024 250410 334036
rect 254670 334024 254676 334036
rect 254728 334024 254734 334076
rect 268746 334024 268752 334076
rect 268804 334064 268810 334076
rect 277949 334067 278007 334073
rect 277949 334064 277961 334067
rect 268804 334036 277961 334064
rect 268804 334024 268810 334036
rect 277949 334033 277961 334036
rect 277995 334033 278007 334067
rect 277949 334027 278007 334033
rect 278869 334067 278927 334073
rect 278869 334033 278881 334067
rect 278915 334064 278927 334067
rect 282362 334064 282368 334076
rect 278915 334036 282368 334064
rect 278915 334033 278927 334036
rect 278869 334027 278927 334033
rect 282362 334024 282368 334036
rect 282420 334024 282426 334076
rect 282457 334067 282515 334073
rect 282457 334033 282469 334067
rect 282503 334064 282515 334067
rect 287698 334064 287704 334076
rect 282503 334036 287704 334064
rect 282503 334033 282515 334036
rect 282457 334027 282515 334033
rect 287698 334024 287704 334036
rect 287756 334024 287762 334076
rect 232498 333956 232504 334008
rect 232556 333996 232562 334008
rect 247313 333999 247371 334005
rect 247313 333996 247325 333999
rect 232556 333968 247325 333996
rect 232556 333956 232562 333968
rect 247313 333965 247325 333968
rect 247359 333965 247371 333999
rect 247313 333959 247371 333965
rect 250530 333956 250536 334008
rect 250588 333996 250594 334008
rect 254486 333996 254492 334008
rect 250588 333968 254492 333996
rect 250588 333956 250594 333968
rect 254486 333956 254492 333968
rect 254544 333956 254550 334008
rect 271414 333956 271420 334008
rect 271472 333996 271478 334008
rect 278038 333996 278044 334008
rect 271472 333968 278044 333996
rect 271472 333956 271478 333968
rect 278038 333956 278044 333968
rect 278096 333956 278102 334008
rect 278317 333999 278375 334005
rect 278317 333965 278329 333999
rect 278363 333996 278375 333999
rect 282733 333999 282791 334005
rect 282733 333996 282745 333999
rect 278363 333968 282745 333996
rect 278363 333965 278375 333968
rect 278317 333959 278375 333965
rect 282733 333965 282745 333968
rect 282779 333965 282791 333999
rect 282733 333959 282791 333965
rect 282914 333956 282920 334008
rect 282972 333996 282978 334008
rect 284386 333996 284392 334008
rect 282972 333968 284392 333996
rect 282972 333956 282978 333968
rect 284386 333956 284392 333968
rect 284444 333956 284450 334008
rect 284481 333999 284539 334005
rect 284481 333965 284493 333999
rect 284527 333996 284539 333999
rect 290642 333996 290648 334008
rect 284527 333968 290648 333996
rect 284527 333965 284539 333968
rect 284481 333959 284539 333965
rect 290642 333956 290648 333968
rect 290700 333956 290706 334008
rect 180702 333888 180708 333940
rect 180760 333928 180766 333940
rect 249613 333931 249671 333937
rect 249613 333928 249625 333931
rect 180760 333900 249625 333928
rect 180760 333888 180766 333900
rect 249613 333897 249625 333900
rect 249659 333897 249671 333931
rect 249613 333891 249671 333897
rect 258537 333931 258595 333937
rect 258537 333897 258549 333931
rect 258583 333928 258595 333931
rect 258810 333928 258816 333940
rect 258583 333900 258816 333928
rect 258583 333897 258595 333900
rect 258537 333891 258595 333897
rect 258810 333888 258816 333900
rect 258868 333888 258874 333940
rect 264790 333888 264796 333940
rect 264848 333928 264854 333940
rect 362954 333928 362960 333940
rect 264848 333900 362960 333928
rect 264848 333888 264854 333900
rect 362954 333888 362960 333900
rect 363012 333888 363018 333940
rect 177942 333820 177948 333872
rect 178000 333860 178006 333872
rect 249426 333860 249432 333872
rect 178000 333832 249432 333860
rect 178000 333820 178006 333832
rect 249426 333820 249432 333832
rect 249484 333820 249490 333872
rect 266357 333863 266415 333869
rect 266357 333829 266369 333863
rect 266403 333860 266415 333863
rect 365714 333860 365720 333872
rect 266403 333832 365720 333860
rect 266403 333829 266415 333832
rect 266357 333823 266415 333829
rect 365714 333820 365720 333832
rect 365772 333820 365778 333872
rect 173802 333752 173808 333804
rect 173860 333792 173866 333804
rect 249150 333792 249156 333804
rect 173860 333764 249156 333792
rect 173860 333752 173866 333764
rect 249150 333752 249156 333764
rect 249208 333752 249214 333804
rect 265710 333752 265716 333804
rect 265768 333792 265774 333804
rect 376754 333792 376760 333804
rect 265768 333764 376760 333792
rect 265768 333752 265774 333764
rect 376754 333752 376760 333764
rect 376812 333752 376818 333804
rect 169570 333684 169576 333736
rect 169628 333724 169634 333736
rect 248785 333727 248843 333733
rect 248785 333724 248797 333727
rect 169628 333696 248797 333724
rect 169628 333684 169634 333696
rect 248785 333693 248797 333696
rect 248831 333693 248843 333727
rect 248785 333687 248843 333693
rect 266078 333684 266084 333736
rect 266136 333724 266142 333736
rect 380894 333724 380900 333736
rect 266136 333696 380900 333724
rect 266136 333684 266142 333696
rect 380894 333684 380900 333696
rect 380952 333684 380958 333736
rect 166902 333616 166908 333668
rect 166960 333656 166966 333668
rect 248509 333659 248567 333665
rect 248509 333656 248521 333659
rect 166960 333628 248521 333656
rect 166960 333616 166966 333628
rect 248509 333625 248521 333628
rect 248555 333625 248567 333659
rect 248509 333619 248567 333625
rect 266633 333659 266691 333665
rect 266633 333625 266645 333659
rect 266679 333656 266691 333659
rect 387794 333656 387800 333668
rect 266679 333628 387800 333656
rect 266679 333625 266691 333628
rect 266633 333619 266691 333625
rect 387794 333616 387800 333628
rect 387852 333616 387858 333668
rect 162762 333548 162768 333600
rect 162820 333588 162826 333600
rect 244737 333591 244795 333597
rect 244737 333588 244749 333591
rect 162820 333560 244749 333588
rect 162820 333548 162826 333560
rect 244737 333557 244749 333560
rect 244783 333557 244795 333591
rect 244737 333551 244795 333557
rect 244918 333548 244924 333600
rect 244976 333588 244982 333600
rect 245746 333588 245752 333600
rect 244976 333560 245752 333588
rect 244976 333548 244982 333560
rect 245746 333548 245752 333560
rect 245804 333548 245810 333600
rect 266446 333548 266452 333600
rect 266504 333588 266510 333600
rect 383654 333588 383660 333600
rect 266504 333560 383660 333588
rect 266504 333548 266510 333560
rect 383654 333548 383660 333560
rect 383712 333548 383718 333600
rect 151722 333480 151728 333532
rect 151780 333520 151786 333532
rect 242250 333520 242256 333532
rect 151780 333492 242256 333520
rect 151780 333480 151786 333492
rect 242250 333480 242256 333492
rect 242308 333480 242314 333532
rect 245381 333523 245439 333529
rect 245381 333489 245393 333523
rect 245427 333520 245439 333523
rect 247126 333520 247132 333532
rect 245427 333492 247132 333520
rect 245427 333489 245439 333492
rect 245381 333483 245439 333489
rect 247126 333480 247132 333492
rect 247184 333480 247190 333532
rect 266909 333523 266967 333529
rect 266909 333489 266921 333523
rect 266955 333520 266967 333523
rect 390646 333520 390652 333532
rect 266955 333492 390652 333520
rect 266955 333489 266967 333492
rect 266909 333483 266967 333489
rect 390646 333480 390652 333492
rect 390704 333480 390710 333532
rect 154482 333412 154488 333464
rect 154540 333452 154546 333464
rect 247494 333452 247500 333464
rect 154540 333424 247500 333452
rect 154540 333412 154546 333424
rect 247494 333412 247500 333424
rect 247552 333412 247558 333464
rect 267737 333455 267795 333461
rect 267737 333421 267749 333455
rect 267783 333452 267795 333455
rect 394694 333452 394700 333464
rect 267783 333424 394700 333452
rect 267783 333421 267795 333424
rect 267737 333415 267795 333421
rect 394694 333412 394700 333424
rect 394752 333412 394758 333464
rect 148962 333344 148968 333396
rect 149020 333384 149026 333396
rect 245381 333387 245439 333393
rect 245381 333384 245393 333387
rect 149020 333356 245393 333384
rect 149020 333344 149026 333356
rect 245381 333353 245393 333356
rect 245427 333353 245439 333387
rect 245930 333384 245936 333396
rect 245381 333347 245439 333353
rect 245580 333356 245936 333384
rect 147582 333276 147588 333328
rect 147640 333316 147646 333328
rect 245580 333316 245608 333356
rect 245930 333344 245936 333356
rect 245988 333344 245994 333396
rect 253382 333344 253388 333396
rect 253440 333384 253446 333396
rect 255314 333384 255320 333396
rect 253440 333356 255320 333384
rect 253440 333344 253446 333356
rect 255314 333344 255320 333356
rect 255372 333344 255378 333396
rect 267550 333344 267556 333396
rect 267608 333384 267614 333396
rect 398834 333384 398840 333396
rect 267608 333356 398840 333384
rect 267608 333344 267614 333356
rect 398834 333344 398840 333356
rect 398892 333344 398898 333396
rect 147640 333288 245608 333316
rect 245657 333319 245715 333325
rect 147640 333276 147646 333288
rect 245657 333285 245669 333319
rect 245703 333316 245715 333319
rect 253934 333316 253940 333328
rect 245703 333288 253940 333316
rect 245703 333285 245715 333288
rect 245657 333279 245715 333285
rect 253934 333276 253940 333288
rect 253992 333276 253998 333328
rect 256970 333276 256976 333328
rect 257028 333316 257034 333328
rect 257982 333316 257988 333328
rect 257028 333288 257988 333316
rect 257028 333276 257034 333288
rect 257982 333276 257988 333288
rect 258040 333276 258046 333328
rect 258077 333319 258135 333325
rect 258077 333285 258089 333319
rect 258123 333316 258135 333319
rect 264422 333316 264428 333328
rect 258123 333288 264428 333316
rect 258123 333285 258135 333288
rect 258077 333279 258135 333285
rect 264422 333276 264428 333288
rect 264480 333276 264486 333328
rect 268105 333319 268163 333325
rect 268105 333285 268117 333319
rect 268151 333316 268163 333319
rect 405734 333316 405740 333328
rect 268151 333288 405740 333316
rect 268151 333285 268163 333288
rect 268105 333279 268163 333285
rect 405734 333276 405740 333288
rect 405792 333276 405798 333328
rect 131022 333208 131028 333260
rect 131080 333248 131086 333260
rect 245562 333248 245568 333260
rect 131080 333220 245568 333248
rect 131080 333208 131086 333220
rect 245562 333208 245568 333220
rect 245620 333208 245626 333260
rect 248509 333251 248567 333257
rect 248509 333217 248521 333251
rect 248555 333248 248567 333251
rect 252922 333248 252928 333260
rect 248555 333220 252928 333248
rect 248555 333217 248567 333220
rect 248509 333211 248567 333217
rect 252922 333208 252928 333220
rect 252980 333208 252986 333260
rect 255222 333248 255228 333260
rect 255183 333220 255228 333248
rect 255222 333208 255228 333220
rect 255280 333208 255286 333260
rect 256050 333208 256056 333260
rect 256108 333248 256114 333260
rect 256602 333248 256608 333260
rect 256108 333220 256608 333248
rect 256108 333208 256114 333220
rect 256602 333208 256608 333220
rect 256660 333208 256666 333260
rect 256881 333251 256939 333257
rect 256881 333217 256893 333251
rect 256927 333248 256939 333251
rect 264698 333248 264704 333260
rect 256927 333220 264704 333248
rect 256927 333217 256939 333220
rect 256881 333211 256939 333217
rect 264698 333208 264704 333220
rect 264756 333208 264762 333260
rect 268565 333251 268623 333257
rect 268565 333217 268577 333251
rect 268611 333248 268623 333251
rect 408494 333248 408500 333260
rect 268611 333220 408500 333248
rect 268611 333217 268623 333220
rect 268565 333211 268623 333217
rect 408494 333208 408500 333220
rect 408552 333208 408558 333260
rect 184842 333140 184848 333192
rect 184900 333180 184906 333192
rect 249886 333180 249892 333192
rect 184900 333152 249892 333180
rect 184900 333140 184906 333152
rect 249886 333140 249892 333152
rect 249944 333140 249950 333192
rect 251910 333140 251916 333192
rect 251968 333180 251974 333192
rect 254946 333180 254952 333192
rect 251968 333152 254952 333180
rect 251968 333140 251974 333152
rect 254946 333140 254952 333152
rect 255004 333140 255010 333192
rect 257062 333140 257068 333192
rect 257120 333180 257126 333192
rect 257433 333183 257491 333189
rect 257433 333180 257445 333183
rect 257120 333152 257445 333180
rect 257120 333140 257126 333152
rect 257433 333149 257445 333152
rect 257479 333149 257491 333183
rect 257433 333143 257491 333149
rect 259546 333140 259552 333192
rect 259604 333180 259610 333192
rect 260561 333183 260619 333189
rect 260561 333180 260573 333183
rect 259604 333152 260573 333180
rect 259604 333140 259610 333152
rect 260561 333149 260573 333152
rect 260607 333149 260619 333183
rect 260561 333143 260619 333149
rect 261202 333140 261208 333192
rect 261260 333180 261266 333192
rect 262125 333183 262183 333189
rect 262125 333180 262137 333183
rect 261260 333152 262137 333180
rect 261260 333140 261266 333152
rect 262125 333149 262137 333152
rect 262171 333149 262183 333183
rect 262125 333143 262183 333149
rect 262858 333140 262864 333192
rect 262916 333180 262922 333192
rect 263686 333180 263692 333192
rect 262916 333152 263692 333180
rect 262916 333140 262922 333152
rect 263686 333140 263692 333152
rect 263744 333140 263750 333192
rect 264517 333183 264575 333189
rect 264517 333149 264529 333183
rect 264563 333180 264575 333183
rect 358814 333180 358820 333192
rect 264563 333152 358820 333180
rect 264563 333149 264575 333152
rect 264517 333143 264575 333149
rect 358814 333140 358820 333152
rect 358872 333140 358878 333192
rect 187602 333072 187608 333124
rect 187660 333112 187666 333124
rect 250162 333112 250168 333124
rect 187660 333084 250168 333112
rect 187660 333072 187666 333084
rect 250162 333072 250168 333084
rect 250220 333072 250226 333124
rect 259457 333115 259515 333121
rect 259457 333081 259469 333115
rect 259503 333112 259515 333115
rect 268381 333115 268439 333121
rect 268381 333112 268393 333115
rect 259503 333084 268393 333112
rect 259503 333081 259515 333084
rect 259457 333075 259515 333081
rect 268381 333081 268393 333084
rect 268427 333081 268439 333115
rect 268381 333075 268439 333081
rect 268841 333115 268899 333121
rect 268841 333081 268853 333115
rect 268887 333112 268899 333115
rect 356054 333112 356060 333124
rect 268887 333084 356060 333112
rect 268887 333081 268899 333084
rect 268841 333075 268899 333081
rect 356054 333072 356060 333084
rect 356112 333072 356118 333124
rect 191742 333004 191748 333056
rect 191800 333044 191806 333056
rect 250438 333044 250444 333056
rect 191800 333016 250444 333044
rect 191800 333004 191806 333016
rect 250438 333004 250444 333016
rect 250496 333004 250502 333056
rect 261113 333047 261171 333053
rect 261113 333013 261125 333047
rect 261159 333044 261171 333047
rect 320174 333044 320180 333056
rect 261159 333016 320180 333044
rect 261159 333013 261171 333016
rect 261113 333007 261171 333013
rect 320174 333004 320180 333016
rect 320232 333004 320238 333056
rect 194410 332936 194416 332988
rect 194468 332976 194474 332988
rect 250806 332976 250812 332988
rect 194468 332948 250812 332976
rect 194468 332936 194474 332948
rect 250806 332936 250812 332948
rect 250864 332936 250870 332988
rect 262677 332979 262735 332985
rect 262677 332945 262689 332979
rect 262723 332976 262735 332979
rect 263226 332976 263232 332988
rect 262723 332948 263232 332976
rect 262723 332945 262735 332948
rect 262677 332939 262735 332945
rect 263226 332936 263232 332948
rect 263284 332936 263290 332988
rect 264146 332936 264152 332988
rect 264204 332976 264210 332988
rect 268657 332979 268715 332985
rect 268657 332976 268669 332979
rect 264204 332948 268669 332976
rect 264204 332936 264210 332948
rect 268657 332945 268669 332948
rect 268703 332945 268715 332979
rect 268657 332939 268715 332945
rect 268749 332979 268807 332985
rect 268749 332945 268761 332979
rect 268795 332976 268807 332979
rect 351914 332976 351920 332988
rect 268795 332948 351920 332976
rect 268795 332945 268807 332948
rect 268749 332939 268807 332945
rect 351914 332936 351920 332948
rect 351972 332936 351978 332988
rect 202782 332868 202788 332920
rect 202840 332908 202846 332920
rect 251361 332911 251419 332917
rect 251361 332908 251373 332911
rect 202840 332880 251373 332908
rect 202840 332868 202846 332880
rect 251361 332877 251373 332880
rect 251407 332877 251419 332911
rect 251361 332871 251419 332877
rect 260469 332911 260527 332917
rect 260469 332877 260481 332911
rect 260515 332908 260527 332911
rect 309134 332908 309140 332920
rect 260515 332880 309140 332908
rect 260515 332877 260527 332880
rect 260469 332871 260527 332877
rect 309134 332868 309140 332880
rect 309192 332868 309198 332920
rect 205542 332800 205548 332852
rect 205600 332840 205606 332852
rect 251637 332843 251695 332849
rect 251637 332840 251649 332843
rect 205600 332812 251649 332840
rect 205600 332800 205606 332812
rect 251637 332809 251649 332812
rect 251683 332809 251695 332843
rect 251637 332803 251695 332809
rect 260742 332800 260748 332852
rect 260800 332840 260806 332852
rect 306374 332840 306380 332852
rect 260800 332812 306380 332840
rect 260800 332800 260806 332812
rect 306374 332800 306380 332812
rect 306432 332800 306438 332852
rect 216582 332732 216588 332784
rect 216640 332772 216646 332784
rect 252554 332772 252560 332784
rect 216640 332744 252560 332772
rect 216640 332732 216646 332744
rect 252554 332732 252560 332744
rect 252612 332732 252618 332784
rect 259730 332732 259736 332784
rect 259788 332772 259794 332784
rect 302234 332772 302240 332784
rect 259788 332744 302240 332772
rect 259788 332732 259794 332744
rect 302234 332732 302240 332744
rect 302292 332732 302298 332784
rect 219250 332664 219256 332716
rect 219308 332704 219314 332716
rect 248509 332707 248567 332713
rect 248509 332704 248521 332707
rect 219308 332676 248521 332704
rect 219308 332664 219314 332676
rect 248509 332673 248521 332676
rect 248555 332673 248567 332707
rect 248509 332667 248567 332673
rect 249150 332664 249156 332716
rect 249208 332704 249214 332716
rect 254210 332704 254216 332716
rect 249208 332676 254216 332704
rect 249208 332664 249214 332676
rect 254210 332664 254216 332676
rect 254268 332664 254274 332716
rect 268381 332707 268439 332713
rect 268381 332673 268393 332707
rect 268427 332704 268439 332707
rect 299474 332704 299480 332716
rect 268427 332676 299480 332704
rect 268427 332673 268439 332676
rect 268381 332667 268439 332673
rect 299474 332664 299480 332676
rect 299532 332664 299538 332716
rect 234522 332596 234528 332648
rect 234580 332636 234586 332648
rect 245657 332639 245715 332645
rect 245657 332636 245669 332639
rect 234580 332608 245669 332636
rect 234580 332596 234586 332608
rect 245657 332605 245669 332608
rect 245703 332605 245715 332639
rect 245657 332599 245715 332605
rect 249978 332596 249984 332648
rect 250036 332636 250042 332648
rect 254854 332636 254860 332648
rect 250036 332608 254860 332636
rect 250036 332596 250042 332608
rect 254854 332596 254860 332608
rect 254912 332596 254918 332648
rect 271046 332596 271052 332648
rect 271104 332636 271110 332648
rect 271509 332639 271567 332645
rect 271509 332636 271521 332639
rect 271104 332608 271521 332636
rect 271104 332596 271110 332608
rect 271509 332605 271521 332608
rect 271555 332605 271567 332639
rect 271509 332599 271567 332605
rect 272334 332596 272340 332648
rect 272392 332636 272398 332648
rect 272886 332636 272892 332648
rect 272392 332608 272892 332636
rect 272392 332596 272398 332608
rect 272886 332596 272892 332608
rect 272944 332596 272950 332648
rect 276474 332596 276480 332648
rect 276532 332636 276538 332648
rect 277210 332636 277216 332648
rect 276532 332608 277216 332636
rect 276532 332596 276538 332608
rect 277210 332596 277216 332608
rect 277268 332596 277274 332648
rect 279602 332596 279608 332648
rect 279660 332636 279666 332648
rect 280249 332639 280307 332645
rect 280249 332636 280261 332639
rect 279660 332608 280261 332636
rect 279660 332596 279666 332608
rect 280249 332605 280261 332608
rect 280295 332605 280307 332639
rect 280249 332599 280307 332605
rect 280341 332639 280399 332645
rect 280341 332605 280353 332639
rect 280387 332636 280399 332639
rect 283558 332636 283564 332648
rect 280387 332608 283564 332636
rect 280387 332605 280399 332608
rect 280341 332599 280399 332605
rect 283558 332596 283564 332608
rect 283616 332596 283622 332648
rect 283742 332596 283748 332648
rect 283800 332636 283806 332648
rect 283926 332636 283932 332648
rect 283800 332608 283932 332636
rect 283800 332596 283806 332608
rect 283926 332596 283932 332608
rect 283984 332596 283990 332648
rect 284110 332596 284116 332648
rect 284168 332636 284174 332648
rect 286686 332636 286692 332648
rect 284168 332608 286692 332636
rect 284168 332596 284174 332608
rect 286686 332596 286692 332608
rect 286744 332596 286750 332648
rect 160002 332528 160008 332580
rect 160060 332568 160066 332580
rect 247954 332568 247960 332580
rect 160060 332540 247960 332568
rect 160060 332528 160066 332540
rect 247954 332528 247960 332540
rect 248012 332528 248018 332580
rect 252462 332528 252468 332580
rect 252520 332568 252526 332580
rect 255406 332568 255412 332580
rect 252520 332540 255412 332568
rect 252520 332528 252526 332540
rect 255406 332528 255412 332540
rect 255464 332528 255470 332580
rect 263689 332571 263747 332577
rect 263689 332537 263701 332571
rect 263735 332568 263747 332571
rect 269482 332568 269488 332580
rect 263735 332540 269488 332568
rect 263735 332537 263747 332540
rect 263689 332531 263747 332537
rect 269482 332528 269488 332540
rect 269540 332528 269546 332580
rect 270405 332571 270463 332577
rect 270405 332537 270417 332571
rect 270451 332568 270463 332571
rect 429838 332568 429844 332580
rect 270451 332540 429844 332568
rect 270451 332537 270463 332540
rect 270405 332531 270463 332537
rect 429838 332528 429844 332540
rect 429896 332528 429902 332580
rect 155862 332460 155868 332512
rect 155920 332500 155926 332512
rect 247678 332500 247684 332512
rect 155920 332472 247684 332500
rect 155920 332460 155926 332472
rect 247678 332460 247684 332472
rect 247736 332460 247742 332512
rect 269390 332460 269396 332512
rect 269448 332500 269454 332512
rect 430574 332500 430580 332512
rect 269448 332472 430580 332500
rect 269448 332460 269454 332472
rect 430574 332460 430580 332472
rect 430632 332460 430638 332512
rect 153102 332392 153108 332444
rect 153160 332432 153166 332444
rect 247402 332432 247408 332444
rect 153160 332404 247408 332432
rect 153160 332392 153166 332404
rect 247402 332392 247408 332404
rect 247460 332392 247466 332444
rect 272978 332392 272984 332444
rect 273036 332432 273042 332444
rect 276382 332432 276388 332444
rect 273036 332404 276388 332432
rect 273036 332392 273042 332404
rect 276382 332392 276388 332404
rect 276440 332392 276446 332444
rect 276566 332392 276572 332444
rect 276624 332432 276630 332444
rect 276845 332435 276903 332441
rect 276845 332432 276857 332435
rect 276624 332404 276857 332432
rect 276624 332392 276630 332404
rect 276845 332401 276857 332404
rect 276891 332401 276903 332435
rect 276845 332395 276903 332401
rect 277305 332435 277363 332441
rect 277305 332401 277317 332435
rect 277351 332432 277363 332435
rect 434714 332432 434720 332444
rect 277351 332404 434720 332432
rect 277351 332401 277363 332404
rect 277305 332395 277363 332401
rect 434714 332392 434720 332404
rect 434772 332392 434778 332444
rect 144822 332324 144828 332376
rect 144880 332364 144886 332376
rect 246758 332364 246764 332376
rect 144880 332336 246764 332364
rect 144880 332324 144886 332336
rect 246758 332324 246764 332336
rect 246816 332324 246822 332376
rect 271049 332367 271107 332373
rect 271049 332333 271061 332367
rect 271095 332364 271107 332367
rect 439590 332364 439596 332376
rect 271095 332336 439596 332364
rect 271095 332333 271107 332336
rect 271049 332327 271107 332333
rect 439590 332324 439596 332336
rect 439648 332324 439654 332376
rect 142062 332256 142068 332308
rect 142120 332296 142126 332308
rect 246482 332296 246488 332308
rect 142120 332268 246488 332296
rect 142120 332256 142126 332268
rect 246482 332256 246488 332268
rect 246540 332256 246546 332308
rect 256786 332256 256792 332308
rect 256844 332296 256850 332308
rect 436830 332296 436836 332308
rect 256844 332268 270494 332296
rect 256844 332256 256850 332268
rect 137922 332188 137928 332240
rect 137980 332228 137986 332240
rect 246206 332228 246212 332240
rect 137980 332200 246212 332228
rect 137980 332188 137986 332200
rect 246206 332188 246212 332200
rect 246264 332188 246270 332240
rect 270466 332228 270494 332268
rect 274192 332268 436836 332296
rect 274192 332228 274220 332268
rect 436830 332256 436836 332268
rect 436888 332256 436894 332308
rect 270466 332200 274220 332228
rect 276201 332231 276259 332237
rect 276201 332197 276213 332231
rect 276247 332228 276259 332231
rect 276934 332228 276940 332240
rect 276247 332200 276940 332228
rect 276247 332197 276259 332200
rect 276201 332191 276259 332197
rect 276934 332188 276940 332200
rect 276992 332188 276998 332240
rect 287793 332231 287851 332237
rect 287793 332197 287805 332231
rect 287839 332228 287851 332231
rect 536926 332228 536932 332240
rect 287839 332200 536932 332228
rect 287839 332197 287851 332200
rect 287793 332191 287851 332197
rect 536926 332188 536932 332200
rect 536984 332188 536990 332240
rect 135162 332120 135168 332172
rect 135220 332160 135226 332172
rect 245749 332163 245807 332169
rect 245749 332160 245761 332163
rect 135220 332132 245761 332160
rect 135220 332120 135226 332132
rect 245749 332129 245761 332132
rect 245795 332129 245807 332163
rect 245749 332123 245807 332129
rect 274174 332120 274180 332172
rect 274232 332160 274238 332172
rect 279602 332160 279608 332172
rect 274232 332132 279608 332160
rect 274232 332120 274238 332132
rect 279602 332120 279608 332132
rect 279660 332120 279666 332172
rect 282181 332163 282239 332169
rect 282181 332129 282193 332163
rect 282227 332160 282239 332163
rect 282362 332160 282368 332172
rect 282227 332132 282368 332160
rect 282227 332129 282239 332132
rect 282181 332123 282239 332129
rect 282362 332120 282368 332132
rect 282420 332120 282426 332172
rect 540330 332160 540336 332172
rect 282886 332132 540336 332160
rect 128170 332052 128176 332104
rect 128228 332092 128234 332104
rect 245289 332095 245347 332101
rect 245289 332092 245301 332095
rect 128228 332064 245301 332092
rect 128228 332052 128234 332064
rect 245289 332061 245301 332064
rect 245335 332061 245347 332095
rect 245289 332055 245347 332061
rect 276385 332095 276443 332101
rect 276385 332061 276397 332095
rect 276431 332092 276443 332095
rect 276842 332092 276848 332104
rect 276431 332064 276848 332092
rect 276431 332061 276443 332064
rect 276385 332055 276443 332061
rect 276842 332052 276848 332064
rect 276900 332052 276906 332104
rect 279234 332052 279240 332104
rect 279292 332092 279298 332104
rect 282886 332092 282914 332132
rect 540330 332120 540336 332132
rect 540388 332120 540394 332172
rect 279292 332064 282914 332092
rect 283101 332095 283159 332101
rect 279292 332052 279298 332064
rect 283101 332061 283113 332095
rect 283147 332092 283159 332095
rect 286597 332095 286655 332101
rect 286597 332092 286609 332095
rect 283147 332064 286609 332092
rect 283147 332061 283159 332064
rect 283101 332055 283159 332061
rect 286597 332061 286609 332064
rect 286643 332061 286655 332095
rect 286597 332055 286655 332061
rect 286689 332095 286747 332101
rect 286689 332061 286701 332095
rect 286735 332092 286747 332095
rect 542998 332092 543004 332104
rect 286735 332064 543004 332092
rect 286735 332061 286747 332064
rect 286689 332055 286747 332061
rect 542998 332052 543004 332064
rect 543056 332052 543062 332104
rect 230382 331984 230388 332036
rect 230440 332024 230446 332036
rect 253569 332027 253627 332033
rect 253569 332024 253581 332027
rect 230440 331996 253581 332024
rect 230440 331984 230446 331996
rect 253569 331993 253581 331996
rect 253615 331993 253627 332027
rect 253569 331987 253627 331993
rect 273901 332027 273959 332033
rect 273901 331993 273913 332027
rect 273947 332024 273959 332027
rect 274174 332024 274180 332036
rect 273947 331996 274180 332024
rect 273947 331993 273959 331996
rect 273901 331987 273959 331993
rect 274174 331984 274180 331996
rect 274232 331984 274238 332036
rect 279326 331984 279332 332036
rect 279384 332024 279390 332036
rect 547138 332024 547144 332036
rect 279384 331996 547144 332024
rect 279384 331984 279390 331996
rect 547138 331984 547144 331996
rect 547196 331984 547202 332036
rect 88242 331916 88248 331968
rect 88300 331956 88306 331968
rect 232866 331956 232872 331968
rect 88300 331928 232872 331956
rect 88300 331916 88306 331928
rect 232866 331916 232872 331928
rect 232924 331916 232930 331968
rect 234706 331916 234712 331968
rect 234764 331956 234770 331968
rect 235810 331956 235816 331968
rect 234764 331928 235816 331956
rect 234764 331916 234770 331928
rect 235810 331916 235816 331928
rect 235868 331916 235874 331968
rect 236454 331916 236460 331968
rect 236512 331956 236518 331968
rect 236917 331959 236975 331965
rect 236917 331956 236929 331959
rect 236512 331928 236929 331956
rect 236512 331916 236518 331928
rect 236917 331925 236929 331928
rect 236963 331925 236975 331959
rect 236917 331919 236975 331925
rect 238110 331916 238116 331968
rect 238168 331956 238174 331968
rect 238665 331959 238723 331965
rect 238665 331956 238677 331959
rect 238168 331928 238677 331956
rect 238168 331916 238174 331928
rect 238665 331925 238677 331928
rect 238711 331925 238723 331959
rect 238665 331919 238723 331925
rect 239398 331916 239404 331968
rect 239456 331956 239462 331968
rect 242805 331959 242863 331965
rect 242805 331956 242817 331959
rect 239456 331928 242817 331956
rect 239456 331916 239462 331928
rect 242805 331925 242817 331928
rect 242851 331925 242863 331959
rect 279234 331956 279240 331968
rect 279195 331928 279240 331956
rect 242805 331919 242863 331925
rect 279234 331916 279240 331928
rect 279292 331916 279298 331968
rect 279789 331959 279847 331965
rect 279789 331925 279801 331959
rect 279835 331956 279847 331959
rect 548518 331956 548524 331968
rect 279835 331928 548524 331956
rect 279835 331925 279847 331928
rect 279789 331919 279847 331925
rect 548518 331916 548524 331928
rect 548576 331916 548582 331968
rect 43530 331848 43536 331900
rect 43588 331888 43594 331900
rect 237834 331888 237840 331900
rect 43588 331860 237840 331888
rect 43588 331848 43594 331860
rect 237834 331848 237840 331860
rect 237892 331848 237898 331900
rect 248325 331891 248383 331897
rect 248325 331888 248337 331891
rect 239416 331860 248337 331888
rect 164142 331780 164148 331832
rect 164200 331820 164206 331832
rect 239416 331820 239444 331860
rect 248325 331857 248337 331860
rect 248371 331857 248383 331891
rect 248325 331851 248383 331857
rect 260834 331848 260840 331900
rect 260892 331888 260898 331900
rect 280154 331888 280160 331900
rect 260892 331860 280160 331888
rect 260892 331848 260898 331860
rect 280154 331848 280160 331860
rect 280212 331848 280218 331900
rect 280249 331891 280307 331897
rect 280249 331857 280261 331891
rect 280295 331888 280307 331891
rect 286689 331891 286747 331897
rect 286689 331888 286701 331891
rect 280295 331860 286701 331888
rect 280295 331857 280307 331860
rect 280249 331851 280307 331857
rect 286689 331857 286701 331860
rect 286735 331857 286747 331891
rect 286689 331851 286747 331857
rect 286870 331848 286876 331900
rect 286928 331888 286934 331900
rect 556154 331888 556160 331900
rect 286928 331860 556160 331888
rect 286928 331848 286934 331860
rect 556154 331848 556160 331860
rect 556212 331848 556218 331900
rect 164200 331792 239444 331820
rect 164200 331780 164206 331792
rect 239490 331780 239496 331832
rect 239548 331820 239554 331832
rect 246298 331820 246304 331832
rect 239548 331792 246304 331820
rect 239548 331780 239554 331792
rect 246298 331780 246304 331792
rect 246356 331780 246362 331832
rect 265342 331780 265348 331832
rect 265400 331820 265406 331832
rect 371234 331820 371240 331832
rect 265400 331792 371240 331820
rect 265400 331780 265406 331792
rect 371234 331780 371240 331792
rect 371292 331780 371298 331832
rect 168282 331712 168288 331764
rect 168340 331752 168346 331764
rect 248506 331752 248512 331764
rect 168340 331724 248512 331752
rect 168340 331712 168346 331724
rect 248506 331712 248512 331724
rect 248564 331712 248570 331764
rect 265069 331755 265127 331761
rect 265069 331721 265081 331755
rect 265115 331752 265127 331755
rect 367094 331752 367100 331764
rect 265115 331724 367100 331752
rect 265115 331721 265127 331724
rect 265069 331715 265127 331721
rect 367094 331712 367100 331724
rect 367152 331712 367158 331764
rect 186130 331644 186136 331696
rect 186188 331684 186194 331696
rect 249886 331684 249892 331696
rect 186188 331656 249892 331684
rect 186188 331644 186194 331656
rect 249886 331644 249892 331656
rect 249944 331644 249950 331696
rect 259638 331644 259644 331696
rect 259696 331684 259702 331696
rect 299566 331684 299572 331696
rect 259696 331656 299572 331684
rect 259696 331644 259702 331656
rect 299566 331644 299572 331656
rect 299624 331644 299630 331696
rect 200022 331576 200028 331628
rect 200080 331616 200086 331628
rect 251174 331616 251180 331628
rect 200080 331588 251180 331616
rect 200080 331576 200086 331588
rect 251174 331576 251180 331588
rect 251232 331576 251238 331628
rect 261110 331576 261116 331628
rect 261168 331616 261174 331628
rect 298094 331616 298100 331628
rect 261168 331588 298100 331616
rect 261168 331576 261174 331588
rect 298094 331576 298100 331588
rect 298152 331576 298158 331628
rect 212442 331508 212448 331560
rect 212500 331548 212506 331560
rect 252278 331548 252284 331560
rect 212500 331520 252284 331548
rect 212500 331508 212506 331520
rect 252278 331508 252284 331520
rect 252336 331508 252342 331560
rect 258629 331551 258687 331557
rect 258629 331517 258641 331551
rect 258675 331548 258687 331551
rect 258675 331520 283236 331548
rect 258675 331517 258687 331520
rect 258629 331511 258687 331517
rect 217962 331440 217968 331492
rect 218020 331480 218026 331492
rect 252646 331480 252652 331492
rect 218020 331452 252652 331480
rect 218020 331440 218026 331452
rect 252646 331440 252652 331452
rect 252704 331440 252710 331492
rect 263502 331440 263508 331492
rect 263560 331480 263566 331492
rect 283101 331483 283159 331489
rect 283101 331480 283113 331483
rect 263560 331452 283113 331480
rect 263560 331440 263566 331452
rect 283101 331449 283113 331452
rect 283147 331449 283159 331483
rect 283208 331480 283236 331520
rect 289814 331480 289820 331492
rect 283208 331452 289820 331480
rect 283101 331443 283159 331449
rect 289814 331440 289820 331452
rect 289872 331440 289878 331492
rect 223482 331372 223488 331424
rect 223540 331412 223546 331424
rect 253198 331412 253204 331424
rect 223540 331384 253204 331412
rect 223540 331372 223546 331384
rect 253198 331372 253204 331384
rect 253256 331372 253262 331424
rect 258442 331372 258448 331424
rect 258500 331412 258506 331424
rect 285674 331412 285680 331424
rect 258500 331384 285680 331412
rect 258500 331372 258506 331384
rect 285674 331372 285680 331384
rect 285732 331372 285738 331424
rect 286597 331415 286655 331421
rect 286597 331381 286609 331415
rect 286643 331412 286655 331415
rect 291194 331412 291200 331424
rect 286643 331384 291200 331412
rect 286643 331381 286655 331384
rect 286597 331375 286655 331381
rect 291194 331372 291200 331384
rect 291252 331372 291258 331424
rect 227622 331304 227628 331356
rect 227680 331344 227686 331356
rect 236641 331347 236699 331353
rect 227680 331316 234614 331344
rect 227680 331304 227686 331316
rect 110322 331236 110328 331288
rect 110380 331276 110386 331288
rect 233602 331276 233608 331288
rect 110380 331248 233608 331276
rect 110380 331236 110386 331248
rect 233602 331236 233608 331248
rect 233660 331236 233666 331288
rect 234586 331276 234614 331316
rect 236641 331313 236653 331347
rect 236687 331344 236699 331347
rect 237282 331344 237288 331356
rect 236687 331316 237288 331344
rect 236687 331313 236699 331316
rect 236641 331307 236699 331313
rect 237282 331304 237288 331316
rect 237340 331304 237346 331356
rect 238938 331304 238944 331356
rect 238996 331344 239002 331356
rect 239858 331344 239864 331356
rect 238996 331316 239864 331344
rect 238996 331304 239002 331316
rect 239858 331304 239864 331316
rect 239916 331304 239922 331356
rect 240686 331304 240692 331356
rect 240744 331344 240750 331356
rect 241057 331347 241115 331353
rect 241057 331344 241069 331347
rect 240744 331316 241069 331344
rect 240744 331304 240750 331316
rect 241057 331313 241069 331316
rect 241103 331313 241115 331347
rect 241057 331307 241115 331313
rect 274361 331347 274419 331353
rect 274361 331313 274373 331347
rect 274407 331344 274419 331347
rect 294598 331344 294604 331356
rect 274407 331316 294604 331344
rect 274407 331313 274419 331316
rect 274361 331307 274419 331313
rect 294598 331304 294604 331316
rect 294656 331304 294662 331356
rect 252738 331276 252744 331288
rect 234586 331248 252744 331276
rect 252738 331236 252744 331248
rect 252796 331236 252802 331288
rect 253198 331236 253204 331288
rect 253256 331276 253262 331288
rect 254029 331279 254087 331285
rect 254029 331276 254041 331279
rect 253256 331248 254041 331276
rect 253256 331236 253262 331248
rect 254029 331245 254041 331248
rect 254075 331245 254087 331279
rect 254029 331239 254087 331245
rect 256513 331279 256571 331285
rect 256513 331245 256525 331279
rect 256559 331276 256571 331279
rect 258258 331276 258264 331288
rect 256559 331248 258264 331276
rect 256559 331245 256571 331248
rect 256513 331239 256571 331245
rect 258258 331236 258264 331248
rect 258316 331236 258322 331288
rect 278774 331236 278780 331288
rect 278832 331276 278838 331288
rect 287793 331279 287851 331285
rect 287793 331276 287805 331279
rect 278832 331248 287805 331276
rect 278832 331236 278838 331248
rect 287793 331245 287805 331248
rect 287839 331245 287851 331279
rect 287793 331239 287851 331245
rect 175182 331168 175188 331220
rect 175240 331208 175246 331220
rect 249334 331208 249340 331220
rect 175240 331180 249340 331208
rect 175240 331168 175246 331180
rect 249334 331168 249340 331180
rect 249392 331168 249398 331220
rect 265618 331168 265624 331220
rect 265676 331208 265682 331220
rect 374086 331208 374092 331220
rect 265676 331180 374092 331208
rect 265676 331168 265682 331180
rect 374086 331168 374092 331180
rect 374144 331168 374150 331220
rect 171042 331100 171048 331152
rect 171100 331140 171106 331152
rect 248969 331143 249027 331149
rect 248969 331140 248981 331143
rect 171100 331112 248981 331140
rect 171100 331100 171106 331112
rect 248969 331109 248981 331112
rect 249015 331109 249027 331143
rect 248969 331103 249027 331109
rect 268197 331143 268255 331149
rect 268197 331109 268209 331143
rect 268243 331140 268255 331143
rect 378134 331140 378140 331152
rect 268243 331112 378140 331140
rect 268243 331109 268255 331112
rect 268197 331103 268255 331109
rect 378134 331100 378140 331112
rect 378192 331100 378198 331152
rect 157242 331032 157248 331084
rect 157300 331072 157306 331084
rect 247586 331072 247592 331084
rect 157300 331044 247592 331072
rect 157300 331032 157306 331044
rect 247586 331032 247592 331044
rect 247644 331032 247650 331084
rect 266170 331032 266176 331084
rect 266228 331072 266234 331084
rect 382366 331072 382372 331084
rect 266228 331044 382372 331072
rect 266228 331032 266234 331044
rect 382366 331032 382372 331044
rect 382424 331032 382430 331084
rect 153010 330964 153016 331016
rect 153068 331004 153074 331016
rect 247310 331004 247316 331016
rect 153068 330976 247316 331004
rect 153068 330964 153074 330976
rect 247310 330964 247316 330976
rect 247368 330964 247374 331016
rect 266541 331007 266599 331013
rect 266541 330973 266553 331007
rect 266587 331004 266599 331007
rect 385034 331004 385040 331016
rect 266587 330976 385040 331004
rect 266587 330973 266599 330976
rect 266541 330967 266599 330973
rect 385034 330964 385040 330976
rect 385092 330964 385098 331016
rect 150342 330896 150348 330948
rect 150400 330936 150406 330948
rect 247034 330936 247040 330948
rect 150400 330908 247040 330936
rect 150400 330896 150406 330908
rect 247034 330896 247040 330908
rect 247092 330896 247098 330948
rect 256694 330896 256700 330948
rect 256752 330936 256758 330948
rect 266354 330936 266360 330948
rect 256752 330908 266360 330936
rect 256752 330896 256758 330908
rect 266354 330896 266360 330908
rect 266412 330896 266418 330948
rect 266817 330939 266875 330945
rect 266817 330905 266829 330939
rect 266863 330936 266875 330939
rect 389174 330936 389180 330948
rect 266863 330908 389180 330936
rect 266863 330905 266875 330908
rect 266817 330899 266875 330905
rect 389174 330896 389180 330908
rect 389232 330896 389238 330948
rect 143442 330828 143448 330880
rect 143500 330868 143506 330880
rect 246666 330868 246672 330880
rect 143500 330840 246672 330868
rect 143500 330828 143506 330840
rect 246666 330828 246672 330840
rect 246724 330828 246730 330880
rect 267090 330828 267096 330880
rect 267148 330868 267154 330880
rect 391934 330868 391940 330880
rect 267148 330840 391940 330868
rect 267148 330828 267154 330840
rect 391934 330828 391940 330840
rect 391992 330828 391998 330880
rect 139302 330760 139308 330812
rect 139360 330800 139366 330812
rect 243170 330800 243176 330812
rect 139360 330772 243176 330800
rect 139360 330760 139366 330772
rect 243170 330760 243176 330772
rect 243228 330760 243234 330812
rect 267369 330803 267427 330809
rect 267369 330769 267381 330803
rect 267415 330800 267427 330803
rect 396074 330800 396080 330812
rect 267415 330772 396080 330800
rect 267415 330769 267427 330772
rect 267369 330763 267427 330769
rect 396074 330760 396080 330772
rect 396132 330760 396138 330812
rect 132402 330692 132408 330744
rect 132460 330732 132466 330744
rect 245654 330732 245660 330744
rect 132460 330704 245660 330732
rect 132460 330692 132466 330704
rect 245654 330692 245660 330704
rect 245712 330692 245718 330744
rect 267642 330692 267648 330744
rect 267700 330732 267706 330744
rect 398926 330732 398932 330744
rect 267700 330704 398932 330732
rect 267700 330692 267706 330704
rect 398926 330692 398932 330704
rect 398984 330692 398990 330744
rect 102042 330624 102048 330676
rect 102100 330664 102106 330676
rect 243265 330667 243323 330673
rect 243265 330664 243277 330667
rect 102100 330636 243277 330664
rect 102100 330624 102106 330636
rect 243265 330633 243277 330636
rect 243311 330633 243323 330667
rect 243265 330627 243323 330633
rect 274269 330667 274327 330673
rect 274269 330633 274281 330667
rect 274315 330664 274327 330667
rect 277305 330667 277363 330673
rect 274315 330636 277256 330664
rect 274315 330633 274327 330636
rect 274269 330627 274327 330633
rect 84102 330556 84108 330608
rect 84160 330596 84166 330608
rect 241698 330596 241704 330608
rect 84160 330568 241704 330596
rect 84160 330556 84166 330568
rect 241698 330556 241704 330568
rect 241756 330556 241762 330608
rect 268654 330556 268660 330608
rect 268712 330596 268718 330608
rect 277228 330596 277256 330636
rect 277305 330633 277317 330667
rect 277351 330664 277363 330667
rect 402974 330664 402980 330676
rect 277351 330636 402980 330664
rect 277351 330633 277363 330636
rect 277305 330627 277363 330633
rect 402974 330624 402980 330636
rect 403032 330624 403038 330676
rect 407206 330596 407212 330608
rect 268712 330568 277164 330596
rect 277228 330568 407212 330596
rect 268712 330556 268718 330568
rect 73062 330488 73068 330540
rect 73120 330528 73126 330540
rect 241238 330528 241244 330540
rect 73120 330500 241244 330528
rect 73120 330488 73126 330500
rect 241238 330488 241244 330500
rect 241296 330488 241302 330540
rect 264609 330531 264667 330537
rect 264609 330497 264621 330531
rect 264655 330497 264667 330531
rect 264609 330491 264667 330497
rect 177850 330420 177856 330472
rect 177908 330460 177914 330472
rect 248417 330463 248475 330469
rect 248417 330460 248429 330463
rect 177908 330432 248429 330460
rect 177908 330420 177914 330432
rect 248417 330429 248429 330432
rect 248463 330429 248475 330463
rect 264624 330460 264652 330491
rect 268286 330488 268292 330540
rect 268344 330528 268350 330540
rect 274269 330531 274327 330537
rect 274269 330528 274281 330531
rect 268344 330500 274281 330528
rect 268344 330488 268350 330500
rect 274269 330497 274281 330500
rect 274315 330497 274327 330531
rect 277136 330528 277164 330568
rect 407206 330556 407212 330568
rect 407264 330556 407270 330608
rect 409874 330528 409880 330540
rect 277136 330500 409880 330528
rect 274269 330491 274327 330497
rect 409874 330488 409880 330500
rect 409932 330488 409938 330540
rect 364334 330460 364340 330472
rect 264624 330432 364340 330460
rect 248417 330423 248475 330429
rect 364334 330420 364340 330432
rect 364392 330420 364398 330472
rect 188982 330352 188988 330404
rect 189040 330392 189046 330404
rect 250254 330392 250260 330404
rect 189040 330364 250260 330392
rect 189040 330352 189046 330364
rect 250254 330352 250260 330364
rect 250312 330352 250318 330404
rect 264606 330352 264612 330404
rect 264664 330392 264670 330404
rect 360194 330392 360200 330404
rect 264664 330364 360200 330392
rect 264664 330352 264670 330364
rect 360194 330352 360200 330364
rect 360252 330352 360258 330404
rect 193122 330284 193128 330336
rect 193180 330324 193186 330336
rect 249981 330327 250039 330333
rect 249981 330324 249993 330327
rect 193180 330296 249993 330324
rect 193180 330284 193186 330296
rect 249981 330293 249993 330296
rect 250027 330293 250039 330327
rect 249981 330287 250039 330293
rect 264241 330327 264299 330333
rect 264241 330293 264253 330327
rect 264287 330324 264299 330327
rect 357434 330324 357440 330336
rect 264287 330296 357440 330324
rect 264287 330293 264299 330296
rect 264241 330287 264299 330293
rect 357434 330284 357440 330296
rect 357492 330284 357498 330336
rect 202690 330216 202696 330268
rect 202748 330256 202754 330268
rect 251545 330259 251603 330265
rect 251545 330256 251557 330259
rect 202748 330228 251557 330256
rect 202748 330216 202754 330228
rect 251545 330225 251557 330228
rect 251591 330225 251603 330259
rect 251545 330219 251603 330225
rect 264330 330216 264336 330268
rect 264388 330256 264394 330268
rect 353294 330256 353300 330268
rect 264388 330228 353300 330256
rect 264388 330216 264394 330228
rect 353294 330216 353300 330228
rect 353352 330216 353358 330268
rect 206922 330148 206928 330200
rect 206980 330188 206986 330200
rect 252094 330188 252100 330200
rect 206980 330160 252100 330188
rect 206980 330148 206986 330160
rect 252094 330148 252100 330160
rect 252152 330148 252158 330200
rect 253290 330148 253296 330200
rect 253348 330188 253354 330200
rect 254394 330188 254400 330200
rect 253348 330160 254400 330188
rect 253348 330148 253354 330160
rect 254394 330148 254400 330160
rect 254452 330148 254458 330200
rect 262582 330148 262588 330200
rect 262640 330188 262646 330200
rect 316126 330188 316132 330200
rect 262640 330160 316132 330188
rect 262640 330148 262646 330160
rect 316126 330148 316132 330160
rect 316184 330148 316190 330200
rect 213822 330080 213828 330132
rect 213880 330120 213886 330132
rect 252370 330120 252376 330132
rect 213880 330092 252376 330120
rect 213880 330080 213886 330092
rect 252370 330080 252376 330092
rect 252428 330080 252434 330132
rect 260558 330080 260564 330132
rect 260616 330120 260622 330132
rect 310514 330120 310520 330132
rect 260616 330092 310520 330120
rect 260616 330080 260622 330092
rect 310514 330080 310520 330092
rect 310572 330080 310578 330132
rect 220722 330012 220728 330064
rect 220780 330052 220786 330064
rect 252830 330052 252836 330064
rect 220780 330024 252836 330052
rect 220780 330012 220786 330024
rect 252830 330012 252836 330024
rect 252888 330012 252894 330064
rect 259822 330012 259828 330064
rect 259880 330052 259886 330064
rect 303614 330052 303620 330064
rect 259880 330024 303620 330052
rect 259880 330012 259886 330024
rect 303614 330012 303620 330024
rect 303672 330012 303678 330064
rect 224862 329944 224868 329996
rect 224920 329984 224926 329996
rect 252649 329987 252707 329993
rect 252649 329984 252661 329987
rect 224920 329956 252661 329984
rect 224920 329944 224926 329956
rect 252649 329953 252661 329956
rect 252695 329953 252707 329987
rect 252649 329947 252707 329953
rect 258994 329944 259000 329996
rect 259052 329984 259058 329996
rect 292666 329984 292672 329996
rect 259052 329956 292672 329984
rect 259052 329944 259058 329956
rect 292666 329944 292672 329956
rect 292724 329944 292730 329996
rect 227530 329876 227536 329928
rect 227588 329916 227594 329928
rect 253385 329919 253443 329925
rect 253385 329916 253397 329919
rect 227588 329888 253397 329916
rect 227588 329876 227594 329888
rect 253385 329885 253397 329888
rect 253431 329885 253443 329919
rect 253385 329879 253443 329885
rect 273346 329876 273352 329928
rect 273404 329916 273410 329928
rect 273714 329916 273720 329928
rect 273404 329888 273720 329916
rect 273404 329876 273410 329888
rect 273714 329876 273720 329888
rect 273772 329876 273778 329928
rect 277670 329876 277676 329928
rect 277728 329916 277734 329928
rect 278314 329916 278320 329928
rect 277728 329888 278320 329916
rect 277728 329876 277734 329888
rect 278314 329876 278320 329888
rect 278372 329876 278378 329928
rect 284294 329876 284300 329928
rect 284352 329916 284358 329928
rect 284938 329916 284944 329928
rect 284352 329888 284944 329916
rect 284352 329876 284358 329888
rect 284938 329876 284944 329888
rect 284996 329876 285002 329928
rect 285490 329876 285496 329928
rect 285548 329916 285554 329928
rect 288342 329916 288348 329928
rect 285548 329888 288348 329916
rect 285548 329876 285554 329888
rect 288342 329876 288348 329888
rect 288400 329876 288406 329928
rect 235258 329808 235264 329860
rect 235316 329848 235322 329860
rect 236457 329851 236515 329857
rect 236457 329848 236469 329851
rect 235316 329820 236469 329848
rect 235316 329808 235322 329820
rect 236457 329817 236469 329820
rect 236503 329817 236515 329851
rect 236457 329811 236515 329817
rect 267734 329808 267740 329860
rect 267792 329848 267798 329860
rect 267792 329820 276152 329848
rect 267792 329808 267798 329820
rect 97902 329740 97908 329792
rect 97960 329780 97966 329792
rect 242894 329780 242900 329792
rect 97960 329752 242900 329780
rect 97960 329740 97966 329752
rect 242894 329740 242900 329752
rect 242952 329740 242958 329792
rect 272061 329783 272119 329789
rect 272061 329749 272073 329783
rect 272107 329780 272119 329783
rect 273898 329780 273904 329792
rect 272107 329752 273904 329780
rect 272107 329749 272119 329752
rect 272061 329743 272119 329749
rect 273898 329740 273904 329752
rect 273956 329740 273962 329792
rect 95050 329672 95056 329724
rect 95108 329712 95114 329724
rect 242618 329712 242624 329724
rect 95108 329684 242624 329712
rect 95108 329672 95114 329684
rect 242618 329672 242624 329684
rect 242676 329672 242682 329724
rect 276124 329712 276152 329820
rect 276290 329740 276296 329792
rect 276348 329780 276354 329792
rect 277302 329780 277308 329792
rect 276348 329752 277308 329780
rect 276348 329740 276354 329752
rect 277302 329740 277308 329752
rect 277360 329740 277366 329792
rect 279142 329740 279148 329792
rect 279200 329780 279206 329792
rect 542354 329780 542360 329792
rect 279200 329752 542360 329780
rect 279200 329740 279206 329752
rect 542354 329740 542360 329752
rect 542412 329740 542418 329792
rect 277213 329715 277271 329721
rect 277213 329712 277225 329715
rect 276124 329684 277225 329712
rect 277213 329681 277225 329684
rect 277259 329681 277271 329715
rect 277213 329675 277271 329681
rect 277578 329672 277584 329724
rect 277636 329712 277642 329724
rect 277946 329712 277952 329724
rect 277636 329684 277952 329712
rect 277636 329672 277642 329684
rect 277946 329672 277952 329684
rect 278004 329672 278010 329724
rect 279970 329672 279976 329724
rect 280028 329712 280034 329724
rect 544378 329712 544384 329724
rect 280028 329684 544384 329712
rect 280028 329672 280034 329684
rect 544378 329672 544384 329684
rect 544436 329672 544442 329724
rect 91002 329604 91008 329656
rect 91060 329644 91066 329656
rect 241793 329647 241851 329653
rect 241793 329644 241805 329647
rect 91060 329616 241805 329644
rect 91060 329604 91066 329616
rect 241793 329613 241805 329616
rect 241839 329613 241851 329647
rect 241793 329607 241851 329613
rect 272705 329647 272763 329653
rect 272705 329613 272717 329647
rect 272751 329644 272763 329647
rect 279694 329644 279700 329656
rect 272751 329616 279700 329644
rect 272751 329613 272763 329616
rect 272705 329607 272763 329613
rect 279694 329604 279700 329616
rect 279752 329604 279758 329656
rect 279786 329604 279792 329656
rect 279844 329644 279850 329656
rect 546494 329644 546500 329656
rect 279844 329616 546500 329644
rect 279844 329604 279850 329616
rect 546494 329604 546500 329616
rect 546552 329604 546558 329656
rect 86862 329536 86868 329588
rect 86920 329576 86926 329588
rect 241882 329576 241888 329588
rect 86920 329548 241888 329576
rect 86920 329536 86926 329548
rect 241882 329536 241888 329548
rect 241940 329536 241946 329588
rect 284478 329536 284484 329588
rect 284536 329576 284542 329588
rect 289630 329576 289636 329588
rect 284536 329548 289636 329576
rect 284536 329536 284542 329548
rect 289630 329536 289636 329548
rect 289688 329536 289694 329588
rect 291749 329579 291807 329585
rect 291749 329545 291761 329579
rect 291795 329576 291807 329579
rect 553394 329576 553400 329588
rect 291795 329548 553400 329576
rect 291795 329545 291807 329548
rect 291749 329539 291807 329545
rect 553394 329536 553400 329548
rect 553452 329536 553458 329588
rect 79962 329468 79968 329520
rect 80020 329508 80026 329520
rect 241422 329508 241428 329520
rect 80020 329480 241428 329508
rect 80020 329468 80026 329480
rect 241422 329468 241428 329480
rect 241480 329468 241486 329520
rect 291841 329511 291899 329517
rect 291841 329477 291853 329511
rect 291887 329508 291899 329511
rect 560294 329508 560300 329520
rect 291887 329480 560300 329508
rect 291887 329477 291899 329480
rect 291841 329471 291899 329477
rect 560294 329468 560300 329480
rect 560352 329468 560358 329520
rect 77202 329400 77208 329452
rect 77260 329440 77266 329452
rect 233234 329440 233240 329452
rect 77260 329412 233240 329440
rect 77260 329400 77266 329412
rect 233234 329400 233240 329412
rect 233292 329400 233298 329452
rect 280522 329400 280528 329452
rect 280580 329440 280586 329452
rect 556246 329440 556252 329452
rect 280580 329412 556252 329440
rect 280580 329400 280586 329412
rect 556246 329400 556252 329412
rect 556304 329400 556310 329452
rect 50338 329332 50344 329384
rect 50396 329372 50402 329384
rect 239030 329372 239036 329384
rect 50396 329344 239036 329372
rect 50396 329332 50402 329344
rect 239030 329332 239036 329344
rect 239088 329332 239094 329384
rect 281074 329332 281080 329384
rect 281132 329372 281138 329384
rect 564526 329372 564532 329384
rect 281132 329344 564532 329372
rect 281132 329332 281138 329344
rect 564526 329332 564532 329344
rect 564584 329332 564590 329384
rect 46198 329264 46204 329316
rect 46256 329304 46262 329316
rect 239493 329307 239551 329313
rect 239493 329304 239505 329307
rect 46256 329276 239505 329304
rect 46256 329264 46262 329276
rect 239493 329273 239505 329276
rect 239539 329273 239551 329307
rect 239493 329267 239551 329273
rect 258166 329264 258172 329316
rect 258224 329304 258230 329316
rect 258442 329304 258448 329316
rect 258224 329276 258448 329304
rect 258224 329264 258230 329276
rect 258442 329264 258448 329276
rect 258500 329264 258506 329316
rect 281258 329264 281264 329316
rect 281316 329304 281322 329316
rect 566458 329304 566464 329316
rect 281316 329276 566464 329304
rect 281316 329264 281322 329276
rect 566458 329264 566464 329276
rect 566516 329264 566522 329316
rect 44818 329196 44824 329248
rect 44876 329236 44882 329248
rect 237466 329236 237472 329248
rect 44876 329208 237472 329236
rect 44876 329196 44882 329208
rect 237466 329196 237472 329208
rect 237524 329196 237530 329248
rect 281721 329239 281779 329245
rect 281721 329205 281733 329239
rect 281767 329236 281779 329239
rect 571334 329236 571340 329248
rect 281767 329208 571340 329236
rect 281767 329205 281779 329208
rect 281721 329199 281779 329205
rect 571334 329196 571340 329208
rect 571392 329196 571398 329248
rect 22738 329128 22744 329180
rect 22796 329168 22802 329180
rect 235994 329168 236000 329180
rect 22796 329140 236000 329168
rect 22796 329128 22802 329140
rect 235994 329128 236000 329140
rect 236052 329128 236058 329180
rect 282822 329128 282828 329180
rect 282880 329168 282886 329180
rect 574094 329168 574100 329180
rect 282880 329140 574100 329168
rect 282880 329128 282886 329140
rect 574094 329128 574100 329140
rect 574152 329128 574158 329180
rect 14458 329060 14464 329112
rect 14516 329100 14522 329112
rect 235902 329100 235908 329112
rect 14516 329072 235908 329100
rect 14516 329060 14522 329072
rect 235902 329060 235908 329072
rect 235960 329060 235966 329112
rect 272889 329103 272947 329109
rect 272889 329069 272901 329103
rect 272935 329100 272947 329103
rect 281074 329100 281080 329112
rect 272935 329072 281080 329100
rect 272935 329069 272947 329072
rect 272889 329063 272947 329069
rect 281074 329060 281080 329072
rect 281132 329060 281138 329112
rect 282454 329060 282460 329112
rect 282512 329100 282518 329112
rect 576118 329100 576124 329112
rect 282512 329072 576124 329100
rect 282512 329060 282518 329072
rect 576118 329060 576124 329072
rect 576176 329060 576182 329112
rect 104802 328992 104808 329044
rect 104860 329032 104866 329044
rect 243722 329032 243728 329044
rect 104860 329004 243728 329032
rect 104860 328992 104866 329004
rect 243722 328992 243728 329004
rect 243780 328992 243786 329044
rect 269206 328992 269212 329044
rect 269264 329032 269270 329044
rect 416774 329032 416780 329044
rect 269264 329004 416780 329032
rect 269264 328992 269270 329004
rect 416774 328992 416780 329004
rect 416832 328992 416838 329044
rect 108942 328924 108948 328976
rect 109000 328964 109006 328976
rect 242529 328967 242587 328973
rect 242529 328964 242541 328967
rect 109000 328936 242541 328964
rect 109000 328924 109006 328936
rect 242529 328933 242541 328936
rect 242575 328933 242587 328967
rect 242529 328927 242587 328933
rect 261386 328924 261392 328976
rect 261444 328924 261450 328976
rect 269577 328967 269635 328973
rect 269577 328933 269589 328967
rect 269623 328964 269635 328967
rect 414014 328964 414020 328976
rect 269623 328936 414020 328964
rect 269623 328933 269635 328936
rect 269577 328927 269635 328933
rect 414014 328924 414020 328936
rect 414072 328924 414078 328976
rect 111702 328856 111708 328908
rect 111760 328896 111766 328908
rect 244090 328896 244096 328908
rect 111760 328868 244096 328896
rect 111760 328856 111766 328868
rect 244090 328856 244096 328868
rect 244148 328856 244154 328908
rect 261404 328896 261432 328924
rect 322934 328896 322940 328908
rect 261404 328868 322940 328896
rect 322934 328856 322940 328868
rect 322992 328856 322998 328908
rect 115842 328788 115848 328840
rect 115900 328828 115906 328840
rect 244366 328828 244372 328840
rect 115900 328800 244372 328828
rect 115900 328788 115906 328800
rect 244366 328788 244372 328800
rect 244424 328788 244430 328840
rect 261389 328831 261447 328837
rect 261389 328797 261401 328831
rect 261435 328828 261447 328831
rect 293954 328828 293960 328840
rect 261435 328800 293960 328828
rect 261435 328797 261447 328800
rect 261389 328791 261447 328797
rect 293954 328788 293960 328800
rect 294012 328788 294018 328840
rect 119890 328720 119896 328772
rect 119948 328760 119954 328772
rect 244734 328760 244740 328772
rect 119948 328732 244740 328760
rect 119948 328720 119954 328732
rect 244734 328720 244740 328732
rect 244792 328720 244798 328772
rect 280614 328720 280620 328772
rect 280672 328760 280678 328772
rect 291841 328763 291899 328769
rect 291841 328760 291853 328763
rect 280672 328732 291853 328760
rect 280672 328720 280678 328732
rect 291841 328729 291853 328732
rect 291887 328729 291899 328763
rect 291841 328723 291899 328729
rect 122742 328652 122748 328704
rect 122800 328692 122806 328704
rect 244921 328695 244979 328701
rect 244921 328692 244933 328695
rect 122800 328664 244933 328692
rect 122800 328652 122806 328664
rect 244921 328661 244933 328664
rect 244967 328661 244979 328695
rect 244921 328655 244979 328661
rect 280433 328695 280491 328701
rect 280433 328661 280445 328695
rect 280479 328692 280491 328695
rect 291749 328695 291807 328701
rect 291749 328692 291761 328695
rect 280479 328664 291761 328692
rect 280479 328661 280491 328664
rect 280433 328655 280491 328661
rect 291749 328661 291761 328664
rect 291795 328661 291807 328695
rect 291749 328655 291807 328661
rect 161382 328584 161388 328636
rect 161440 328624 161446 328636
rect 248046 328624 248052 328636
rect 161440 328596 248052 328624
rect 161440 328584 161446 328596
rect 248046 328584 248052 328596
rect 248104 328584 248110 328636
rect 86218 328380 86224 328432
rect 86276 328420 86282 328432
rect 241790 328420 241796 328432
rect 86276 328392 241796 328420
rect 86276 328380 86282 328392
rect 241790 328380 241796 328392
rect 241848 328380 241854 328432
rect 80698 328312 80704 328364
rect 80756 328352 80762 328364
rect 240870 328352 240876 328364
rect 80756 328324 240876 328352
rect 80756 328312 80762 328324
rect 240870 328312 240876 328324
rect 240928 328312 240934 328364
rect 266630 328312 266636 328364
rect 266688 328352 266694 328364
rect 386414 328352 386420 328364
rect 266688 328324 386420 328352
rect 266688 328312 266694 328324
rect 386414 328312 386420 328324
rect 386472 328312 386478 328364
rect 75178 328244 75184 328296
rect 75236 328284 75242 328296
rect 241054 328284 241060 328296
rect 75236 328256 241060 328284
rect 75236 328244 75242 328256
rect 241054 328244 241060 328256
rect 241112 328244 241118 328296
rect 267182 328244 267188 328296
rect 267240 328284 267246 328296
rect 393314 328284 393320 328296
rect 267240 328256 393320 328284
rect 267240 328244 267246 328256
rect 393314 328244 393320 328256
rect 393372 328244 393378 328296
rect 70210 328176 70216 328228
rect 70268 328216 70274 328228
rect 240594 328216 240600 328228
rect 70268 328188 240600 328216
rect 70268 328176 70274 328188
rect 240594 328176 240600 328188
rect 240652 328176 240658 328228
rect 267826 328176 267832 328228
rect 267884 328216 267890 328228
rect 400214 328216 400220 328228
rect 267884 328188 400220 328216
rect 267884 328176 267890 328188
rect 400214 328176 400220 328188
rect 400272 328176 400278 328228
rect 68278 328108 68284 328160
rect 68336 328148 68342 328160
rect 240318 328148 240324 328160
rect 68336 328120 240324 328148
rect 68336 328108 68342 328120
rect 240318 328108 240324 328120
rect 240376 328108 240382 328160
rect 283466 328108 283472 328160
rect 283524 328148 283530 328160
rect 447042 328148 447048 328160
rect 283524 328120 447048 328148
rect 283524 328108 283530 328120
rect 447042 328108 447048 328120
rect 447100 328108 447106 328160
rect 62758 328040 62764 328092
rect 62816 328080 62822 328092
rect 238938 328080 238944 328092
rect 62816 328052 238944 328080
rect 62816 328040 62822 328052
rect 238938 328040 238944 328052
rect 238996 328040 239002 328092
rect 283834 328040 283840 328092
rect 283892 328080 283898 328092
rect 476022 328080 476028 328092
rect 283892 328052 476028 328080
rect 283892 328040 283898 328052
rect 476022 328040 476028 328052
rect 476080 328040 476086 328092
rect 57238 327972 57244 328024
rect 57296 328012 57302 328024
rect 238846 328012 238852 328024
rect 57296 327984 238852 328012
rect 57296 327972 57302 327984
rect 238846 327972 238852 327984
rect 238904 327972 238910 328024
rect 282546 327972 282552 328024
rect 282604 328012 282610 328024
rect 476574 328012 476580 328024
rect 282604 327984 476580 328012
rect 282604 327972 282610 327984
rect 476574 327972 476580 327984
rect 476632 327972 476638 328024
rect 51718 327904 51724 327956
rect 51776 327944 51782 327956
rect 237190 327944 237196 327956
rect 51776 327916 237196 327944
rect 51776 327904 51782 327916
rect 237190 327904 237196 327916
rect 237248 327904 237254 327956
rect 283374 327904 283380 327956
rect 283432 327944 283438 327956
rect 481726 327944 481732 327956
rect 283432 327916 481732 327944
rect 283432 327904 283438 327916
rect 481726 327904 481732 327916
rect 481784 327904 481790 327956
rect 53742 327836 53748 327888
rect 53800 327876 53806 327888
rect 239306 327876 239312 327888
rect 53800 327848 239312 327876
rect 53800 327836 53806 327848
rect 239306 327836 239312 327848
rect 239364 327836 239370 327888
rect 283650 327836 283656 327888
rect 283708 327876 283714 327888
rect 484854 327876 484860 327888
rect 283708 327848 484860 327876
rect 283708 327836 283714 327848
rect 484854 327836 484860 327848
rect 484912 327836 484918 327888
rect 11698 327768 11704 327820
rect 11756 327808 11762 327820
rect 234890 327808 234896 327820
rect 11756 327780 234896 327808
rect 11756 327768 11762 327780
rect 234890 327768 234896 327780
rect 234948 327768 234954 327820
rect 283926 327768 283932 327820
rect 283984 327808 283990 327820
rect 490558 327808 490564 327820
rect 283984 327780 490564 327808
rect 283984 327768 283990 327780
rect 490558 327768 490564 327780
rect 490616 327768 490622 327820
rect 10318 327700 10324 327752
rect 10376 327740 10382 327752
rect 235626 327740 235632 327752
rect 10376 327712 235632 327740
rect 10376 327700 10382 327712
rect 235626 327700 235632 327712
rect 235684 327700 235690 327752
rect 283742 327700 283748 327752
rect 283800 327740 283806 327752
rect 492674 327740 492680 327752
rect 283800 327712 492680 327740
rect 283800 327700 283806 327712
rect 492674 327700 492680 327712
rect 492732 327700 492738 327752
rect 93118 327632 93124 327684
rect 93176 327672 93182 327684
rect 242434 327672 242440 327684
rect 93176 327644 242440 327672
rect 93176 327632 93182 327644
rect 242434 327632 242440 327644
rect 242492 327632 242498 327684
rect 99282 327564 99288 327616
rect 99340 327604 99346 327616
rect 243814 327604 243820 327616
rect 99340 327576 243820 327604
rect 99340 327564 99346 327576
rect 243814 327564 243820 327576
rect 243872 327564 243878 327616
rect 195882 327496 195888 327548
rect 195940 327536 195946 327548
rect 250898 327536 250904 327548
rect 195940 327508 250904 327536
rect 195940 327496 195946 327508
rect 250898 327496 250904 327508
rect 250956 327496 250962 327548
rect 231762 327428 231768 327480
rect 231820 327468 231826 327480
rect 253750 327468 253756 327480
rect 231820 327440 253756 327468
rect 231820 327428 231826 327440
rect 253750 327428 253756 327440
rect 253808 327428 253814 327480
rect 215938 327360 215944 327412
rect 215996 327400 216002 327412
rect 236454 327400 236460 327412
rect 215996 327372 236460 327400
rect 215996 327360 216002 327372
rect 236454 327360 236460 327372
rect 236512 327360 236518 327412
rect 125502 327020 125508 327072
rect 125560 327060 125566 327072
rect 245102 327060 245108 327072
rect 125560 327032 245108 327060
rect 125560 327020 125566 327032
rect 245102 327020 245108 327032
rect 245160 327020 245166 327072
rect 124122 326952 124128 327004
rect 124180 326992 124186 327004
rect 243446 326992 243452 327004
rect 124180 326964 243452 326992
rect 124180 326952 124186 326964
rect 243446 326952 243452 326964
rect 243504 326952 243510 327004
rect 115198 326884 115204 326936
rect 115256 326924 115262 326936
rect 243262 326924 243268 326936
rect 115256 326896 243268 326924
rect 115256 326884 115262 326896
rect 243262 326884 243268 326896
rect 243320 326884 243326 326936
rect 106918 326816 106924 326868
rect 106976 326856 106982 326868
rect 238662 326856 238668 326868
rect 106976 326828 238668 326856
rect 106976 326816 106982 326828
rect 238662 326816 238668 326828
rect 238720 326816 238726 326868
rect 107562 326748 107568 326800
rect 107620 326788 107626 326800
rect 243630 326788 243636 326800
rect 107620 326760 243636 326788
rect 107620 326748 107626 326760
rect 243630 326748 243636 326760
rect 243688 326748 243694 326800
rect 106182 326680 106188 326732
rect 106240 326720 106246 326732
rect 242158 326720 242164 326732
rect 106240 326692 242164 326720
rect 106240 326680 106246 326692
rect 242158 326680 242164 326692
rect 242216 326680 242222 326732
rect 83458 326612 83464 326664
rect 83516 326652 83522 326664
rect 242710 326652 242716 326664
rect 83516 326624 242716 326652
rect 83516 326612 83522 326624
rect 242710 326612 242716 326624
rect 242768 326612 242774 326664
rect 63402 326544 63408 326596
rect 63460 326584 63466 326596
rect 239122 326584 239128 326596
rect 63460 326556 239128 326584
rect 63460 326544 63466 326556
rect 239122 326544 239128 326556
rect 239180 326544 239186 326596
rect 58618 326476 58624 326528
rect 58676 326516 58682 326528
rect 237742 326516 237748 326528
rect 58676 326488 237748 326516
rect 58676 326476 58682 326488
rect 237742 326476 237748 326488
rect 237800 326476 237806 326528
rect 255682 326476 255688 326528
rect 255740 326516 255746 326528
rect 255740 326488 263594 326516
rect 255740 326476 255746 326488
rect 47578 326408 47584 326460
rect 47636 326448 47642 326460
rect 237558 326448 237564 326460
rect 47636 326420 237564 326448
rect 47636 326408 47642 326420
rect 237558 326408 237564 326420
rect 237616 326408 237622 326460
rect 255406 326408 255412 326460
rect 255464 326448 255470 326460
rect 255590 326448 255596 326460
rect 255464 326420 255596 326448
rect 255464 326408 255470 326420
rect 255590 326408 255596 326420
rect 255648 326408 255654 326460
rect 255958 326408 255964 326460
rect 256016 326408 256022 326460
rect 257430 326408 257436 326460
rect 257488 326448 257494 326460
rect 257614 326448 257620 326460
rect 257488 326420 257620 326448
rect 257488 326408 257494 326420
rect 257614 326408 257620 326420
rect 257672 326408 257678 326460
rect 257890 326408 257896 326460
rect 257948 326408 257954 326460
rect 260006 326408 260012 326460
rect 260064 326448 260070 326460
rect 260190 326448 260196 326460
rect 260064 326420 260196 326448
rect 260064 326408 260070 326420
rect 260190 326408 260196 326420
rect 260248 326408 260254 326460
rect 26878 326340 26884 326392
rect 26936 326380 26942 326392
rect 234706 326380 234712 326392
rect 26936 326352 234712 326380
rect 26936 326340 26942 326352
rect 234706 326340 234712 326352
rect 234764 326340 234770 326392
rect 234982 326340 234988 326392
rect 235040 326380 235046 326392
rect 235350 326380 235356 326392
rect 235040 326352 235356 326380
rect 235040 326340 235046 326352
rect 235350 326340 235356 326352
rect 235408 326340 235414 326392
rect 236730 326340 236736 326392
rect 236788 326380 236794 326392
rect 237282 326380 237288 326392
rect 236788 326352 237288 326380
rect 236788 326340 236794 326352
rect 237282 326340 237288 326352
rect 237340 326340 237346 326392
rect 246022 326340 246028 326392
rect 246080 326380 246086 326392
rect 246206 326380 246212 326392
rect 246080 326352 246212 326380
rect 246080 326340 246086 326352
rect 246206 326340 246212 326352
rect 246264 326340 246270 326392
rect 248782 326340 248788 326392
rect 248840 326380 248846 326392
rect 249702 326380 249708 326392
rect 248840 326352 249708 326380
rect 248840 326340 248846 326352
rect 249702 326340 249708 326352
rect 249760 326340 249766 326392
rect 250162 326340 250168 326392
rect 250220 326380 250226 326392
rect 251082 326380 251088 326392
rect 250220 326352 251088 326380
rect 250220 326340 250226 326352
rect 251082 326340 251088 326352
rect 251140 326340 251146 326392
rect 254578 326204 254584 326256
rect 254636 326244 254642 326256
rect 255222 326244 255228 326256
rect 254636 326216 255228 326244
rect 254636 326204 254642 326216
rect 255222 326204 255228 326216
rect 255280 326204 255286 326256
rect 255866 326204 255872 326256
rect 255924 326244 255930 326256
rect 255976 326244 256004 326408
rect 256326 326340 256332 326392
rect 256384 326380 256390 326392
rect 256510 326380 256516 326392
rect 256384 326352 256516 326380
rect 256384 326340 256390 326352
rect 256510 326340 256516 326352
rect 256568 326340 256574 326392
rect 257908 326312 257936 326408
rect 262306 326340 262312 326392
rect 262364 326380 262370 326392
rect 263134 326380 263140 326392
rect 262364 326352 263140 326380
rect 262364 326340 262370 326352
rect 263134 326340 263140 326352
rect 263192 326340 263198 326392
rect 263566 326380 263594 326488
rect 267274 326476 267280 326528
rect 267332 326516 267338 326528
rect 267332 326488 273254 326516
rect 267332 326476 267338 326488
rect 269482 326408 269488 326460
rect 269540 326448 269546 326460
rect 269850 326448 269856 326460
rect 269540 326420 269856 326448
rect 269540 326408 269546 326420
rect 269850 326408 269856 326420
rect 269908 326408 269914 326460
rect 271414 326408 271420 326460
rect 271472 326448 271478 326460
rect 271690 326448 271696 326460
rect 271472 326420 271696 326448
rect 271472 326408 271478 326420
rect 271690 326408 271696 326420
rect 271748 326408 271754 326460
rect 272702 326448 272708 326460
rect 272663 326420 272708 326448
rect 272702 326408 272708 326420
rect 272760 326408 272766 326460
rect 273226 326448 273254 326488
rect 329834 326448 329840 326460
rect 273226 326420 329840 326448
rect 329834 326408 329840 326420
rect 329892 326408 329898 326460
rect 436922 326380 436928 326392
rect 263566 326352 436928 326380
rect 436922 326340 436928 326352
rect 436980 326340 436986 326392
rect 257724 326284 257936 326312
rect 257724 326256 257752 326284
rect 255924 326216 256004 326244
rect 255924 326204 255930 326216
rect 257706 326204 257712 326256
rect 257764 326204 257770 326256
rect 257798 326204 257804 326256
rect 257856 326244 257862 326256
rect 257982 326244 257988 326256
rect 257856 326216 257988 326244
rect 257856 326204 257862 326216
rect 257982 326204 257988 326216
rect 258040 326204 258046 326256
rect 260006 326204 260012 326256
rect 260064 326244 260070 326256
rect 260466 326244 260472 326256
rect 260064 326216 260472 326244
rect 260064 326204 260070 326216
rect 260466 326204 260472 326216
rect 260524 326204 260530 326256
rect 180150 325728 180156 325780
rect 180208 325768 180214 325780
rect 236730 325768 236736 325780
rect 180208 325740 236736 325768
rect 180208 325728 180214 325740
rect 236730 325728 236736 325740
rect 236788 325728 236794 325780
rect 50430 325660 50436 325712
rect 50488 325700 50494 325712
rect 235350 325700 235356 325712
rect 50488 325672 235356 325700
rect 50488 325660 50494 325672
rect 235350 325660 235356 325672
rect 235408 325660 235414 325712
rect 443638 325592 443644 325644
rect 443696 325632 443702 325644
rect 580166 325632 580172 325644
rect 443696 325604 580172 325632
rect 443696 325592 443702 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 5442 324912 5448 324964
rect 5500 324952 5506 324964
rect 235074 324952 235080 324964
rect 5500 324924 235080 324952
rect 5500 324912 5506 324924
rect 235074 324912 235080 324924
rect 235132 324912 235138 324964
rect 269666 324912 269672 324964
rect 269724 324952 269730 324964
rect 270034 324952 270040 324964
rect 269724 324924 270040 324952
rect 269724 324912 269730 324924
rect 270034 324912 270040 324924
rect 270092 324912 270098 324964
rect 113082 323552 113088 323604
rect 113140 323592 113146 323604
rect 240962 323592 240968 323604
rect 113140 323564 240968 323592
rect 113140 323552 113146 323564
rect 240962 323552 240968 323564
rect 241020 323552 241026 323604
rect 254486 323144 254492 323196
rect 254544 323184 254550 323196
rect 254762 323184 254768 323196
rect 254544 323156 254768 323184
rect 254544 323144 254550 323156
rect 254762 323144 254768 323156
rect 254820 323144 254826 323196
rect 255498 322940 255504 322992
rect 255556 322980 255562 322992
rect 255774 322980 255780 322992
rect 255556 322952 255780 322980
rect 255556 322940 255562 322952
rect 255774 322940 255780 322952
rect 255832 322940 255838 322992
rect 467098 322872 467104 322924
rect 467156 322912 467162 322924
rect 467156 322884 470594 322912
rect 467156 322872 467162 322884
rect 470566 322844 470594 322884
rect 471238 322872 471244 322924
rect 471296 322912 471302 322924
rect 474737 322915 474795 322921
rect 474737 322912 474749 322915
rect 471296 322884 474749 322912
rect 471296 322872 471302 322884
rect 474737 322881 474749 322884
rect 474783 322881 474795 322915
rect 474737 322875 474795 322881
rect 479518 322872 479524 322924
rect 479576 322912 479582 322924
rect 480622 322912 480628 322924
rect 479576 322884 480628 322912
rect 479576 322872 479582 322884
rect 480622 322872 480628 322884
rect 480680 322872 480686 322924
rect 472250 322844 472256 322856
rect 470566 322816 472256 322844
rect 472250 322804 472256 322816
rect 472308 322804 472314 322856
rect 473998 322804 474004 322856
rect 474056 322844 474062 322856
rect 479150 322844 479156 322856
rect 474056 322816 479156 322844
rect 474056 322804 474062 322816
rect 479150 322804 479156 322816
rect 479208 322804 479214 322856
rect 232682 322736 232688 322788
rect 232740 322776 232746 322788
rect 496814 322776 496820 322788
rect 232740 322748 496820 322776
rect 232740 322736 232746 322748
rect 496814 322736 496820 322748
rect 496872 322736 496878 322788
rect 232590 322668 232596 322720
rect 232648 322708 232654 322720
rect 494238 322708 494244 322720
rect 232648 322680 494244 322708
rect 232648 322668 232654 322680
rect 494238 322668 494244 322680
rect 494296 322668 494302 322720
rect 464338 322600 464344 322652
rect 464396 322640 464402 322652
rect 469398 322640 469404 322652
rect 464396 322612 469404 322640
rect 464396 322600 464402 322612
rect 469398 322600 469404 322612
rect 469456 322600 469462 322652
rect 472618 322600 472624 322652
rect 472676 322640 472682 322652
rect 474550 322640 474556 322652
rect 472676 322612 474556 322640
rect 472676 322600 472682 322612
rect 474550 322600 474556 322612
rect 474608 322600 474614 322652
rect 474737 322643 474795 322649
rect 474737 322609 474749 322643
rect 474783 322640 474795 322643
rect 506934 322640 506940 322652
rect 474783 322612 506940 322640
rect 474783 322609 474795 322612
rect 474737 322603 474795 322609
rect 506934 322600 506940 322612
rect 506992 322600 506998 322652
rect 468478 322532 468484 322584
rect 468536 322572 468542 322584
rect 504174 322572 504180 322584
rect 468536 322544 504180 322572
rect 468536 322532 468542 322544
rect 504174 322532 504180 322544
rect 504232 322532 504238 322584
rect 272702 322504 272708 322516
rect 272663 322476 272708 322504
rect 272702 322464 272708 322476
rect 272760 322464 272766 322516
rect 284754 322464 284760 322516
rect 284812 322504 284818 322516
rect 505462 322504 505468 322516
rect 284812 322476 505468 322504
rect 284812 322464 284818 322476
rect 505462 322464 505468 322476
rect 505520 322464 505526 322516
rect 285306 322396 285312 322448
rect 285364 322436 285370 322448
rect 498654 322436 498660 322448
rect 285364 322408 498660 322436
rect 285364 322396 285370 322408
rect 498654 322396 498660 322408
rect 498712 322396 498718 322448
rect 285398 322328 285404 322380
rect 285456 322368 285462 322380
rect 498194 322368 498200 322380
rect 285456 322340 498200 322368
rect 285456 322328 285462 322340
rect 498194 322328 498200 322340
rect 498252 322328 498258 322380
rect 287606 322260 287612 322312
rect 287664 322300 287670 322312
rect 484394 322300 484400 322312
rect 287664 322272 484400 322300
rect 287664 322260 287670 322272
rect 484394 322260 484400 322272
rect 484452 322260 484458 322312
rect 233142 322192 233148 322244
rect 233200 322232 233206 322244
rect 253014 322232 253020 322244
rect 233200 322204 253020 322232
rect 233200 322192 233206 322204
rect 253014 322192 253020 322204
rect 253072 322192 253078 322244
rect 447042 322192 447048 322244
rect 447100 322232 447106 322244
rect 495526 322232 495532 322244
rect 447100 322204 495532 322232
rect 447100 322192 447106 322204
rect 495526 322192 495532 322204
rect 495584 322192 495590 322244
rect 519538 322192 519544 322244
rect 519596 322232 519602 322244
rect 537110 322232 537116 322244
rect 519596 322204 537116 322232
rect 519596 322192 519602 322204
rect 537110 322192 537116 322204
rect 537168 322192 537174 322244
rect 465718 322124 465724 322176
rect 465776 322164 465782 322176
rect 501046 322164 501052 322176
rect 465776 322136 501052 322164
rect 465776 322124 465782 322136
rect 501046 322124 501052 322136
rect 501104 322124 501110 322176
rect 447778 322056 447784 322108
rect 447836 322096 447842 322108
rect 470686 322096 470692 322108
rect 447836 322068 470692 322096
rect 447836 322056 447842 322068
rect 470686 322056 470692 322068
rect 470744 322056 470750 322108
rect 476022 322056 476028 322108
rect 476080 322096 476086 322108
rect 492214 322096 492220 322108
rect 476080 322068 492220 322096
rect 476080 322056 476086 322068
rect 492214 322056 492220 322068
rect 492272 322056 492278 322108
rect 449158 321988 449164 322040
rect 449216 322028 449222 322040
rect 471974 322028 471980 322040
rect 449216 322000 471980 322028
rect 449216 321988 449222 322000
rect 471974 321988 471980 322000
rect 472032 321988 472038 322040
rect 233234 321920 233240 321972
rect 233292 321960 233298 321972
rect 503254 321960 503260 321972
rect 233292 321932 503260 321960
rect 233292 321920 233298 321932
rect 503254 321920 503260 321932
rect 503312 321920 503318 321972
rect 232774 321852 232780 321904
rect 232832 321892 232838 321904
rect 500678 321892 500684 321904
rect 232832 321864 500684 321892
rect 232832 321852 232838 321864
rect 500678 321852 500684 321864
rect 500736 321852 500742 321904
rect 232222 321784 232228 321836
rect 232280 321824 232286 321836
rect 475470 321824 475476 321836
rect 232280 321796 475476 321824
rect 232280 321784 232286 321796
rect 475470 321784 475476 321796
rect 475528 321784 475534 321836
rect 232406 321716 232412 321768
rect 232464 321756 232470 321768
rect 478230 321756 478236 321768
rect 232464 321728 478236 321756
rect 232464 321716 232470 321728
rect 478230 321716 478236 321728
rect 478288 321716 478294 321768
rect 481726 321580 481732 321632
rect 481784 321620 481790 321632
rect 488166 321620 488172 321632
rect 481784 321592 488172 321620
rect 481784 321580 481790 321592
rect 488166 321580 488172 321592
rect 488224 321580 488230 321632
rect 530026 321580 530032 321632
rect 530084 321620 530090 321632
rect 530670 321620 530676 321632
rect 530084 321592 530676 321620
rect 530084 321580 530090 321592
rect 530670 321580 530676 321592
rect 530728 321620 530734 321632
rect 537202 321620 537208 321632
rect 530728 321592 537208 321620
rect 530728 321580 530734 321592
rect 537202 321580 537208 321592
rect 537260 321580 537266 321632
rect 286778 320832 286784 320884
rect 286836 320872 286842 320884
rect 580994 320872 581000 320884
rect 286836 320844 581000 320872
rect 286836 320832 286842 320844
rect 580994 320832 581000 320844
rect 581052 320832 581058 320884
rect 251634 320152 251640 320204
rect 251692 320192 251698 320204
rect 252002 320192 252008 320204
rect 251692 320164 252008 320192
rect 251692 320152 251698 320164
rect 252002 320152 252008 320164
rect 252060 320152 252066 320204
rect 3510 320084 3516 320136
rect 3568 320124 3574 320136
rect 14642 320124 14648 320136
rect 3568 320096 14648 320124
rect 3568 320084 3574 320096
rect 14642 320084 14648 320096
rect 14700 320084 14706 320136
rect 547230 313216 547236 313268
rect 547288 313256 547294 313268
rect 580166 313256 580172 313268
rect 547288 313228 580172 313256
rect 547288 313216 547294 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3510 306280 3516 306332
rect 3568 306320 3574 306332
rect 35250 306320 35256 306332
rect 3568 306292 35256 306320
rect 3568 306280 3574 306292
rect 35250 306280 35256 306292
rect 35308 306280 35314 306332
rect 537478 299412 537484 299464
rect 537536 299452 537542 299464
rect 580166 299452 580172 299464
rect 537536 299424 580172 299452
rect 537536 299412 537542 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 3050 293904 3056 293956
rect 3108 293944 3114 293956
rect 33870 293944 33876 293956
rect 3108 293916 33876 293944
rect 3108 293904 3114 293916
rect 33870 293904 33876 293916
rect 33928 293904 33934 293956
rect 246298 274592 246304 274644
rect 246356 274632 246362 274644
rect 437474 274632 437480 274644
rect 246356 274604 437480 274632
rect 246356 274592 246362 274604
rect 437474 274592 437480 274604
rect 437532 274592 437538 274644
rect 540422 273164 540428 273216
rect 540480 273204 540486 273216
rect 579982 273204 579988 273216
rect 540480 273176 579988 273204
rect 540480 273164 540486 273176
rect 579982 273164 579988 273176
rect 580040 273164 580046 273216
rect 245194 272484 245200 272536
rect 245252 272524 245258 272536
rect 436646 272524 436652 272536
rect 245252 272496 436652 272524
rect 245252 272484 245258 272496
rect 436646 272484 436652 272496
rect 436704 272484 436710 272536
rect 248598 271804 248604 271856
rect 248656 271844 248662 271856
rect 436830 271844 436836 271856
rect 248656 271816 436836 271844
rect 248656 271804 248662 271816
rect 436830 271804 436836 271816
rect 436888 271804 436894 271856
rect 250714 270444 250720 270496
rect 250772 270484 250778 270496
rect 436830 270484 436836 270496
rect 250772 270456 436836 270484
rect 250772 270444 250778 270456
rect 436830 270444 436836 270456
rect 436888 270444 436894 270496
rect 268562 269764 268568 269816
rect 268620 269804 268626 269816
rect 357526 269804 357532 269816
rect 268620 269776 357532 269804
rect 268620 269764 268626 269776
rect 357526 269764 357532 269776
rect 357584 269764 357590 269816
rect 436922 269016 436928 269068
rect 436980 269056 436986 269068
rect 437290 269056 437296 269068
rect 436980 269028 437296 269056
rect 436980 269016 436986 269028
rect 437290 269016 437296 269028
rect 437348 269016 437354 269068
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 17310 267696 17316 267708
rect 3568 267668 17316 267696
rect 3568 267656 3574 267668
rect 17310 267656 17316 267668
rect 17368 267656 17374 267708
rect 245102 266976 245108 267028
rect 245160 267016 245166 267028
rect 436094 267016 436100 267028
rect 245160 266988 436100 267016
rect 245160 266976 245166 266988
rect 436094 266976 436100 266988
rect 436152 266976 436158 267028
rect 544470 259360 544476 259412
rect 544528 259400 544534 259412
rect 580166 259400 580172 259412
rect 544528 259372 580172 259400
rect 544528 259360 544534 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 36630 255252 36636 255264
rect 3200 255224 36636 255252
rect 3200 255212 3206 255224
rect 36630 255212 36636 255224
rect 36688 255212 36694 255264
rect 232038 248344 232044 248396
rect 232096 248384 232102 248396
rect 436094 248384 436100 248396
rect 232096 248356 436100 248384
rect 232096 248344 232102 248356
rect 436094 248344 436100 248356
rect 436152 248344 436158 248396
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 18690 241448 18696 241460
rect 3568 241420 18696 241448
rect 3568 241408 3574 241420
rect 18690 241408 18696 241420
rect 18748 241408 18754 241460
rect 282638 240728 282644 240780
rect 282696 240768 282702 240780
rect 439130 240768 439136 240780
rect 282696 240740 439136 240768
rect 282696 240728 282702 240740
rect 439130 240728 439136 240740
rect 439188 240728 439194 240780
rect 297726 239980 297732 240032
rect 297784 240020 297790 240032
rect 435913 240023 435971 240029
rect 297784 239992 431954 240020
rect 297784 239980 297790 239992
rect 431926 239952 431954 239992
rect 435913 239989 435925 240023
rect 435959 240020 435971 240023
rect 439866 240020 439872 240032
rect 435959 239992 439872 240020
rect 435959 239989 435971 239992
rect 435913 239983 435971 239989
rect 439866 239980 439872 239992
rect 439924 239980 439930 240032
rect 445662 239952 445668 239964
rect 431926 239924 445668 239952
rect 445662 239912 445668 239924
rect 445720 239912 445726 239964
rect 538490 239952 538496 239964
rect 445772 239924 538496 239952
rect 445772 239896 445800 239924
rect 538490 239912 538496 239924
rect 538548 239912 538554 239964
rect 438670 239844 438676 239896
rect 438728 239884 438734 239896
rect 445573 239887 445631 239893
rect 445573 239884 445585 239887
rect 438728 239856 445585 239884
rect 438728 239844 438734 239856
rect 445573 239853 445585 239856
rect 445619 239853 445631 239887
rect 445573 239847 445631 239853
rect 445754 239844 445760 239896
rect 445812 239844 445818 239896
rect 445849 239887 445907 239893
rect 445849 239853 445861 239887
rect 445895 239884 445907 239887
rect 522666 239884 522672 239896
rect 445895 239856 522672 239884
rect 445895 239853 445907 239856
rect 445849 239847 445907 239853
rect 522666 239844 522672 239856
rect 522724 239844 522730 239896
rect 438762 239776 438768 239828
rect 438820 239816 438826 239828
rect 445665 239819 445723 239825
rect 445665 239816 445677 239819
rect 438820 239788 445677 239816
rect 438820 239776 438826 239788
rect 445665 239785 445677 239788
rect 445711 239785 445723 239819
rect 445665 239779 445723 239785
rect 445941 239819 445999 239825
rect 445941 239785 445953 239819
rect 445987 239816 445999 239819
rect 523126 239816 523132 239828
rect 445987 239788 523132 239816
rect 445987 239785 445999 239788
rect 445941 239779 445999 239785
rect 523126 239776 523132 239788
rect 523184 239776 523190 239828
rect 438578 239708 438584 239760
rect 438636 239748 438642 239760
rect 523034 239748 523040 239760
rect 438636 239720 523040 239748
rect 438636 239708 438642 239720
rect 523034 239708 523040 239720
rect 523092 239708 523098 239760
rect 284846 239640 284852 239692
rect 284904 239680 284910 239692
rect 435913 239683 435971 239689
rect 435913 239680 435925 239683
rect 284904 239652 435925 239680
rect 284904 239640 284910 239652
rect 435913 239649 435925 239652
rect 435959 239649 435971 239683
rect 435913 239643 435971 239649
rect 436002 239640 436008 239692
rect 436060 239680 436066 239692
rect 445754 239680 445760 239692
rect 436060 239652 445760 239680
rect 436060 239640 436066 239652
rect 445754 239640 445760 239652
rect 445812 239640 445818 239692
rect 445846 239640 445852 239692
rect 445904 239680 445910 239692
rect 451090 239680 451096 239692
rect 445904 239652 451096 239680
rect 445904 239640 445910 239652
rect 451090 239640 451096 239652
rect 451148 239640 451154 239692
rect 451182 239640 451188 239692
rect 451240 239680 451246 239692
rect 456058 239680 456064 239692
rect 451240 239652 456064 239680
rect 451240 239640 451246 239652
rect 456058 239640 456064 239652
rect 456116 239640 456122 239692
rect 456153 239683 456211 239689
rect 456153 239649 456165 239683
rect 456199 239680 456211 239683
rect 537202 239680 537208 239692
rect 456199 239652 537208 239680
rect 456199 239649 456211 239652
rect 456153 239643 456211 239649
rect 537202 239640 537208 239652
rect 537260 239640 537266 239692
rect 437382 239572 437388 239624
rect 437440 239612 437446 239624
rect 505002 239612 505008 239624
rect 437440 239584 505008 239612
rect 437440 239572 437446 239584
rect 505002 239572 505008 239584
rect 505060 239572 505066 239624
rect 299014 239504 299020 239556
rect 299072 239544 299078 239556
rect 299072 239516 452700 239544
rect 299072 239504 299078 239516
rect 298922 239436 298928 239488
rect 298980 239476 298986 239488
rect 452562 239476 452568 239488
rect 298980 239448 452568 239476
rect 298980 239436 298986 239448
rect 452562 239436 452568 239448
rect 452620 239436 452626 239488
rect 452672 239476 452700 239516
rect 452746 239504 452752 239556
rect 452804 239544 452810 239556
rect 455969 239547 456027 239553
rect 455969 239544 455981 239547
rect 452804 239516 455981 239544
rect 452804 239504 452810 239516
rect 455969 239513 455981 239516
rect 456015 239513 456027 239547
rect 455969 239507 456027 239513
rect 456058 239504 456064 239556
rect 456116 239544 456122 239556
rect 460934 239544 460940 239556
rect 456116 239516 460940 239544
rect 456116 239504 456122 239516
rect 460934 239504 460940 239516
rect 460992 239504 460998 239556
rect 461026 239504 461032 239556
rect 461084 239544 461090 239556
rect 464709 239547 464767 239553
rect 464709 239544 464721 239547
rect 461084 239516 464721 239544
rect 461084 239504 461090 239516
rect 464709 239513 464721 239516
rect 464755 239513 464767 239547
rect 464709 239507 464767 239513
rect 464801 239547 464859 239553
rect 464801 239513 464813 239547
rect 464847 239544 464859 239547
rect 473170 239544 473176 239556
rect 464847 239516 473176 239544
rect 464847 239513 464859 239516
rect 464801 239507 464859 239513
rect 473170 239504 473176 239516
rect 473228 239504 473234 239556
rect 464985 239479 465043 239485
rect 452672 239448 464936 239476
rect 288158 239368 288164 239420
rect 288216 239408 288222 239420
rect 464801 239411 464859 239417
rect 464801 239408 464813 239411
rect 288216 239380 464813 239408
rect 288216 239368 288222 239380
rect 464801 239377 464813 239380
rect 464847 239377 464859 239411
rect 464908 239408 464936 239448
rect 464985 239445 464997 239479
rect 465031 239476 465043 239479
rect 479334 239476 479340 239488
rect 465031 239448 479340 239476
rect 465031 239445 465043 239448
rect 464985 239439 465043 239445
rect 479334 239436 479340 239448
rect 479392 239436 479398 239488
rect 471974 239408 471980 239420
rect 464908 239380 471980 239408
rect 464801 239371 464859 239377
rect 471974 239368 471980 239380
rect 472032 239368 472038 239420
rect 288066 239300 288072 239352
rect 288124 239340 288130 239352
rect 475654 239340 475660 239352
rect 288124 239312 475660 239340
rect 288124 239300 288130 239312
rect 475654 239300 475660 239312
rect 475712 239300 475718 239352
rect 297542 239232 297548 239284
rect 297600 239272 297606 239284
rect 487890 239272 487896 239284
rect 297600 239244 487896 239272
rect 297600 239232 297606 239244
rect 487890 239232 487896 239244
rect 487948 239232 487954 239284
rect 297450 239164 297456 239216
rect 297508 239204 297514 239216
rect 501874 239204 501880 239216
rect 297508 239176 501880 239204
rect 297508 239164 297514 239176
rect 501874 239164 501880 239176
rect 501932 239164 501938 239216
rect 297358 239096 297364 239148
rect 297416 239136 297422 239148
rect 503070 239136 503076 239148
rect 297416 239108 503076 239136
rect 297416 239096 297422 239108
rect 503070 239096 503076 239108
rect 503128 239096 503134 239148
rect 298738 239028 298744 239080
rect 298796 239068 298802 239080
rect 505554 239068 505560 239080
rect 298796 239040 505560 239068
rect 298796 239028 298802 239040
rect 505554 239028 505560 239040
rect 505612 239028 505618 239080
rect 292206 238960 292212 239012
rect 292264 239000 292270 239012
rect 506750 239000 506756 239012
rect 292264 238972 506756 239000
rect 292264 238960 292270 238972
rect 506750 238960 506756 238972
rect 506808 238960 506814 239012
rect 232958 238892 232964 238944
rect 233016 238932 233022 238944
rect 495618 238932 495624 238944
rect 233016 238904 495624 238932
rect 233016 238892 233022 238904
rect 495618 238892 495624 238904
rect 495676 238892 495682 238944
rect 233050 238824 233056 238876
rect 233108 238864 233114 238876
rect 496814 238864 496820 238876
rect 233108 238836 496820 238864
rect 233108 238824 233114 238836
rect 496814 238824 496820 238836
rect 496872 238824 496878 238876
rect 234430 238756 234436 238808
rect 234488 238796 234494 238808
rect 500494 238796 500500 238808
rect 234488 238768 500500 238796
rect 234488 238756 234494 238768
rect 500494 238756 500500 238768
rect 500552 238756 500558 238808
rect 296254 238688 296260 238740
rect 296312 238728 296318 238740
rect 485406 238728 485412 238740
rect 296312 238700 485412 238728
rect 296312 238688 296318 238700
rect 485406 238688 485412 238700
rect 485464 238688 485470 238740
rect 291838 238620 291844 238672
rect 291896 238660 291902 238672
rect 477678 238660 477684 238672
rect 291896 238632 477684 238660
rect 291896 238620 291902 238632
rect 477678 238620 477684 238632
rect 477736 238620 477742 238672
rect 296070 238552 296076 238604
rect 296128 238592 296134 238604
rect 484394 238592 484400 238604
rect 296128 238564 484400 238592
rect 296128 238552 296134 238564
rect 484394 238552 484400 238564
rect 484452 238552 484458 238604
rect 292022 238484 292028 238536
rect 292080 238524 292086 238536
rect 483382 238524 483388 238536
rect 292080 238496 483388 238524
rect 292080 238484 292086 238496
rect 483382 238484 483388 238496
rect 483440 238484 483446 238536
rect 290550 238416 290556 238468
rect 290608 238456 290614 238468
rect 482278 238456 482284 238468
rect 290608 238428 482284 238456
rect 290608 238416 290614 238428
rect 482278 238416 482284 238428
rect 482336 238416 482342 238468
rect 292298 238348 292304 238400
rect 292356 238388 292362 238400
rect 484854 238388 484860 238400
rect 292356 238360 484860 238388
rect 292356 238348 292362 238360
rect 484854 238348 484860 238360
rect 484912 238348 484918 238400
rect 293586 238280 293592 238332
rect 293644 238320 293650 238332
rect 488166 238320 488172 238332
rect 293644 238292 488172 238320
rect 293644 238280 293650 238292
rect 488166 238280 488172 238292
rect 488224 238280 488230 238332
rect 292114 238212 292120 238264
rect 292172 238252 292178 238264
rect 485958 238252 485964 238264
rect 292172 238224 485964 238252
rect 292172 238212 292178 238224
rect 485958 238212 485964 238224
rect 486016 238212 486022 238264
rect 293494 238144 293500 238196
rect 293552 238184 293558 238196
rect 491662 238184 491668 238196
rect 293552 238156 491668 238184
rect 293552 238144 293558 238156
rect 491662 238144 491668 238156
rect 491720 238144 491726 238196
rect 259086 238076 259092 238128
rect 259144 238116 259150 238128
rect 284386 238116 284392 238128
rect 259144 238088 284392 238116
rect 259144 238076 259150 238088
rect 284386 238076 284392 238088
rect 284444 238076 284450 238128
rect 294782 238076 294788 238128
rect 294840 238116 294846 238128
rect 495158 238116 495164 238128
rect 294840 238088 495164 238116
rect 294840 238076 294846 238088
rect 495158 238076 495164 238088
rect 495216 238076 495222 238128
rect 258810 238008 258816 238060
rect 258868 238048 258874 238060
rect 287054 238048 287060 238060
rect 258868 238020 287060 238048
rect 258868 238008 258874 238020
rect 287054 238008 287060 238020
rect 287112 238008 287118 238060
rect 293402 238008 293408 238060
rect 293460 238048 293466 238060
rect 492766 238048 492772 238060
rect 293460 238020 492772 238048
rect 293460 238008 293466 238020
rect 492766 238008 492772 238020
rect 492824 238008 492830 238060
rect 296346 237940 296352 237992
rect 296404 237980 296410 237992
rect 481726 237980 481732 237992
rect 296404 237952 481732 237980
rect 296404 237940 296410 237952
rect 481726 237940 481732 237952
rect 481784 237940 481790 237992
rect 291930 237872 291936 237924
rect 291988 237912 291994 237924
rect 476574 237912 476580 237924
rect 291988 237884 476580 237912
rect 291988 237872 291994 237884
rect 476574 237872 476580 237884
rect 476632 237872 476638 237924
rect 296438 237804 296444 237856
rect 296496 237844 296502 237856
rect 480622 237844 480628 237856
rect 296496 237816 480628 237844
rect 296496 237804 296502 237816
rect 480622 237804 480628 237816
rect 480680 237804 480686 237856
rect 294874 237736 294880 237788
rect 294932 237776 294938 237788
rect 467190 237776 467196 237788
rect 294932 237748 467196 237776
rect 294932 237736 294938 237748
rect 467190 237736 467196 237748
rect 467248 237736 467254 237788
rect 296530 237668 296536 237720
rect 296588 237708 296594 237720
rect 467834 237708 467840 237720
rect 296588 237680 467840 237708
rect 296588 237668 296594 237680
rect 467834 237668 467840 237680
rect 467892 237668 467898 237720
rect 294690 237600 294696 237652
rect 294748 237640 294754 237652
rect 465074 237640 465080 237652
rect 294748 237612 465080 237640
rect 294748 237600 294754 237612
rect 465074 237600 465080 237612
rect 465132 237600 465138 237652
rect 292390 237532 292396 237584
rect 292448 237572 292454 237584
rect 462314 237572 462320 237584
rect 292448 237544 462320 237572
rect 292448 237532 292454 237544
rect 462314 237532 462320 237544
rect 462372 237532 462378 237584
rect 295058 237464 295064 237516
rect 295116 237504 295122 237516
rect 463694 237504 463700 237516
rect 295116 237476 463700 237504
rect 295116 237464 295122 237476
rect 463694 237464 463700 237476
rect 463752 237464 463758 237516
rect 438302 237396 438308 237448
rect 438360 237436 438366 237448
rect 485774 237436 485780 237448
rect 438360 237408 485780 237436
rect 438360 237396 438366 237408
rect 485774 237396 485780 237408
rect 485832 237396 485838 237448
rect 233786 237328 233792 237380
rect 233844 237368 233850 237380
rect 470594 237368 470600 237380
rect 233844 237340 470600 237368
rect 233844 237328 233850 237340
rect 470594 237328 470600 237340
rect 470652 237328 470658 237380
rect 505002 237328 505008 237380
rect 505060 237368 505066 237380
rect 521654 237368 521660 237380
rect 505060 237340 521660 237368
rect 505060 237328 505066 237340
rect 521654 237328 521660 237340
rect 521712 237328 521718 237380
rect 233694 237260 233700 237312
rect 233752 237300 233758 237312
rect 467834 237300 467840 237312
rect 233752 237272 467840 237300
rect 233752 237260 233758 237272
rect 467834 237260 467840 237272
rect 467892 237260 467898 237312
rect 288342 237192 288348 237244
rect 288400 237232 288406 237244
rect 503714 237232 503720 237244
rect 288400 237204 503720 237232
rect 288400 237192 288406 237204
rect 503714 237192 503720 237204
rect 503772 237192 503778 237244
rect 289630 237124 289636 237176
rect 289688 237164 289694 237176
rect 498194 237164 498200 237176
rect 289688 237136 498200 237164
rect 289688 237124 289694 237136
rect 498194 237124 498200 237136
rect 498252 237124 498258 237176
rect 285214 237056 285220 237108
rect 285272 237096 285278 237108
rect 492674 237096 492680 237108
rect 285272 237068 492680 237096
rect 285272 237056 285278 237068
rect 492674 237056 492680 237068
rect 492732 237056 492738 237108
rect 288250 236988 288256 237040
rect 288308 237028 288314 237040
rect 494054 237028 494060 237040
rect 288308 237000 494060 237028
rect 288308 236988 288314 237000
rect 494054 236988 494060 237000
rect 494112 236988 494118 237040
rect 286686 236920 286692 236972
rect 286744 236960 286750 236972
rect 491294 236960 491300 236972
rect 286744 236932 491300 236960
rect 286744 236920 286750 236932
rect 491294 236920 491300 236932
rect 491352 236920 491358 236972
rect 286594 236852 286600 236904
rect 286652 236892 286658 236904
rect 490282 236892 490288 236904
rect 286652 236864 490288 236892
rect 286652 236852 286658 236864
rect 490282 236852 490288 236864
rect 490340 236852 490346 236904
rect 282086 236784 282092 236836
rect 282144 236824 282150 236836
rect 473354 236824 473360 236836
rect 282144 236796 473360 236824
rect 282144 236784 282150 236796
rect 473354 236784 473360 236796
rect 473412 236784 473418 236836
rect 258442 236716 258448 236768
rect 258500 236756 258506 236768
rect 282914 236756 282920 236768
rect 258500 236728 282920 236756
rect 258500 236716 258506 236728
rect 282914 236716 282920 236728
rect 282972 236716 282978 236768
rect 296162 236716 296168 236768
rect 296220 236756 296226 236768
rect 485774 236756 485780 236768
rect 296220 236728 485780 236756
rect 296220 236716 296226 236728
rect 485774 236716 485780 236728
rect 485832 236716 485838 236768
rect 281810 236648 281816 236700
rect 281868 236688 281874 236700
rect 469214 236688 469220 236700
rect 281868 236660 469220 236688
rect 281868 236648 281874 236660
rect 469214 236648 469220 236660
rect 469272 236648 469278 236700
rect 289446 236580 289452 236632
rect 289504 236620 289510 236632
rect 471974 236620 471980 236632
rect 289504 236592 471980 236620
rect 289504 236580 289510 236592
rect 471974 236580 471980 236592
rect 472032 236580 472038 236632
rect 298830 236512 298836 236564
rect 298888 236552 298894 236564
rect 476114 236552 476120 236564
rect 298888 236524 476120 236552
rect 298888 236512 298894 236524
rect 476114 236512 476120 236524
rect 476172 236512 476178 236564
rect 289538 236444 289544 236496
rect 289596 236484 289602 236496
rect 461118 236484 461124 236496
rect 289596 236456 461124 236484
rect 289596 236444 289602 236456
rect 461118 236444 461124 236456
rect 461176 236444 461182 236496
rect 294966 236376 294972 236428
rect 295024 236416 295030 236428
rect 465074 236416 465080 236428
rect 295024 236388 465080 236416
rect 295024 236376 295030 236388
rect 465074 236376 465080 236388
rect 465132 236376 465138 236428
rect 344554 236308 344560 236360
rect 344612 236348 344618 236360
rect 488534 236348 488540 236360
rect 344612 236320 488540 236348
rect 344612 236308 344618 236320
rect 488534 236308 488540 236320
rect 488592 236308 488598 236360
rect 344462 236240 344468 236292
rect 344520 236280 344526 236292
rect 474734 236280 474740 236292
rect 344520 236252 474740 236280
rect 344520 236240 344526 236252
rect 474734 236240 474740 236252
rect 474792 236240 474798 236292
rect 344370 236172 344376 236224
rect 344428 236212 344434 236224
rect 470870 236212 470876 236224
rect 344428 236184 470876 236212
rect 344428 236172 344434 236184
rect 470870 236172 470876 236184
rect 470928 236172 470934 236224
rect 440234 236104 440240 236156
rect 440292 236144 440298 236156
rect 495434 236144 495440 236156
rect 440292 236116 495440 236144
rect 440292 236104 440298 236116
rect 495434 236104 495440 236116
rect 495492 236104 495498 236156
rect 439130 236036 439136 236088
rect 439188 236076 439194 236088
rect 469214 236076 469220 236088
rect 439188 236048 469220 236076
rect 439188 236036 439194 236048
rect 469214 236036 469220 236048
rect 469272 236036 469278 236088
rect 275370 235900 275376 235952
rect 275428 235940 275434 235952
rect 488534 235940 488540 235952
rect 275428 235912 488540 235940
rect 275428 235900 275434 235912
rect 488534 235900 488540 235912
rect 488592 235900 488598 235952
rect 274818 235832 274824 235884
rect 274876 235872 274882 235884
rect 490558 235872 490564 235884
rect 274876 235844 490564 235872
rect 274876 235832 274882 235844
rect 490558 235832 490564 235844
rect 490616 235832 490622 235884
rect 275554 235764 275560 235816
rect 275612 235804 275618 235816
rect 493318 235804 493324 235816
rect 275612 235776 493324 235804
rect 275612 235764 275618 235776
rect 493318 235764 493324 235776
rect 493376 235764 493382 235816
rect 276658 235696 276664 235748
rect 276716 235736 276722 235748
rect 497458 235736 497464 235748
rect 276716 235708 497464 235736
rect 276716 235696 276722 235708
rect 497458 235696 497464 235708
rect 497516 235696 497522 235748
rect 276566 235628 276572 235680
rect 276624 235668 276630 235680
rect 500218 235668 500224 235680
rect 276624 235640 500224 235668
rect 276624 235628 276630 235640
rect 500218 235628 500224 235640
rect 500276 235628 500282 235680
rect 276474 235560 276480 235612
rect 276532 235600 276538 235612
rect 501598 235600 501604 235612
rect 276532 235572 501604 235600
rect 276532 235560 276538 235572
rect 501598 235560 501604 235572
rect 501656 235560 501662 235612
rect 276750 235492 276756 235544
rect 276808 235532 276814 235544
rect 502334 235532 502340 235544
rect 276808 235504 502340 235532
rect 276808 235492 276814 235504
rect 502334 235492 502340 235504
rect 502392 235492 502398 235544
rect 276842 235424 276848 235476
rect 276900 235464 276906 235476
rect 506474 235464 506480 235476
rect 276900 235436 506480 235464
rect 276900 235424 276906 235436
rect 506474 235424 506480 235436
rect 506532 235424 506538 235476
rect 277394 235356 277400 235408
rect 277452 235396 277458 235408
rect 508498 235396 508504 235408
rect 277452 235368 508504 235396
rect 277452 235356 277458 235368
rect 508498 235356 508504 235368
rect 508556 235356 508562 235408
rect 278130 235288 278136 235340
rect 278188 235328 278194 235340
rect 512638 235328 512644 235340
rect 278188 235300 512644 235328
rect 278188 235288 278194 235300
rect 512638 235288 512644 235300
rect 512696 235288 512702 235340
rect 277946 235220 277952 235272
rect 278004 235260 278010 235272
rect 520274 235260 520280 235272
rect 278004 235232 520280 235260
rect 278004 235220 278010 235232
rect 520274 235220 520280 235232
rect 520332 235220 520338 235272
rect 273990 235152 273996 235204
rect 274048 235192 274054 235204
rect 484394 235192 484400 235204
rect 274048 235164 484400 235192
rect 274048 235152 274054 235164
rect 484394 235152 484400 235164
rect 484452 235152 484458 235204
rect 275462 235084 275468 235136
rect 275520 235124 275526 235136
rect 483658 235124 483664 235136
rect 275520 235096 483664 235124
rect 275520 235084 275526 235096
rect 483658 235084 483664 235096
rect 483716 235084 483722 235136
rect 274082 235016 274088 235068
rect 274140 235056 274146 235068
rect 481726 235056 481732 235068
rect 274140 235028 481732 235056
rect 274140 235016 274146 235028
rect 481726 235016 481732 235028
rect 481784 235016 481790 235068
rect 274174 234948 274180 235000
rect 274232 234988 274238 235000
rect 475378 234988 475384 235000
rect 274232 234960 475384 234988
rect 274232 234948 274238 234960
rect 475378 234948 475384 234960
rect 475436 234948 475442 235000
rect 273254 234880 273260 234932
rect 273312 234920 273318 234932
rect 472618 234920 472624 234932
rect 273312 234892 472624 234920
rect 273312 234880 273318 234892
rect 472618 234880 472624 234892
rect 472676 234880 472682 234932
rect 272794 234812 272800 234864
rect 272852 234852 272858 234864
rect 459554 234852 459560 234864
rect 272852 234824 459560 234852
rect 272852 234812 272858 234824
rect 459554 234812 459560 234824
rect 459612 234812 459618 234864
rect 272886 234744 272892 234796
rect 272944 234784 272950 234796
rect 456886 234784 456892 234796
rect 272944 234756 456892 234784
rect 272944 234744 272950 234756
rect 456886 234744 456892 234756
rect 456944 234744 456950 234796
rect 271230 234676 271236 234728
rect 271288 234716 271294 234728
rect 441614 234716 441620 234728
rect 271288 234688 441620 234716
rect 271288 234676 271294 234688
rect 441614 234676 441620 234688
rect 441672 234676 441678 234728
rect 418890 234608 418896 234660
rect 418948 234648 418954 234660
rect 477494 234648 477500 234660
rect 418948 234620 477500 234648
rect 418948 234608 418954 234620
rect 477494 234608 477500 234620
rect 477552 234608 477558 234660
rect 272978 234540 272984 234592
rect 273036 234580 273042 234592
rect 466454 234580 466460 234592
rect 273036 234552 466460 234580
rect 273036 234540 273042 234552
rect 466454 234540 466460 234552
rect 466512 234540 466518 234592
rect 274358 234472 274364 234524
rect 274416 234512 274422 234524
rect 470594 234512 470600 234524
rect 274416 234484 470600 234512
rect 274416 234472 274422 234484
rect 470594 234472 470600 234484
rect 470652 234472 470658 234524
rect 274266 234404 274272 234456
rect 274324 234444 274330 234456
rect 472710 234444 472716 234456
rect 274324 234416 472716 234444
rect 274324 234404 274330 234416
rect 472710 234404 472716 234416
rect 472768 234404 472774 234456
rect 273622 234336 273628 234388
rect 273680 234376 273686 234388
rect 476758 234376 476764 234388
rect 273680 234348 476764 234376
rect 273680 234336 273686 234348
rect 476758 234336 476764 234348
rect 476816 234336 476822 234388
rect 273346 234268 273352 234320
rect 273404 234308 273410 234320
rect 479518 234308 479524 234320
rect 273404 234280 479524 234308
rect 273404 234268 273410 234280
rect 479518 234268 479524 234280
rect 479576 234268 479582 234320
rect 275738 234200 275744 234252
rect 275796 234240 275802 234252
rect 490006 234240 490012 234252
rect 275796 234212 490012 234240
rect 275796 234200 275802 234212
rect 490006 234200 490012 234212
rect 490064 234200 490070 234252
rect 275002 234132 275008 234184
rect 275060 234172 275066 234184
rect 492674 234172 492680 234184
rect 275060 234144 492680 234172
rect 275060 234132 275066 234144
rect 492674 234132 492680 234144
rect 492732 234132 492738 234184
rect 275646 234064 275652 234116
rect 275704 234104 275710 234116
rect 496814 234104 496820 234116
rect 275704 234076 496820 234104
rect 275704 234064 275710 234076
rect 496814 234064 496820 234076
rect 496872 234064 496878 234116
rect 276934 233996 276940 234048
rect 276992 234036 276998 234048
rect 503714 234036 503720 234048
rect 276992 234008 503720 234036
rect 276992 233996 276998 234008
rect 503714 233996 503720 234008
rect 503772 233996 503778 234048
rect 277026 233928 277032 233980
rect 277084 233968 277090 233980
rect 506566 233968 506572 233980
rect 277084 233940 506572 233968
rect 277084 233928 277090 233940
rect 506566 233928 506572 233940
rect 506624 233928 506630 233980
rect 278222 233860 278228 233912
rect 278280 233900 278286 233912
rect 519538 233900 519544 233912
rect 278280 233872 519544 233900
rect 278280 233860 278286 233872
rect 519538 233860 519544 233872
rect 519596 233860 519602 233912
rect 271874 233792 271880 233844
rect 271932 233832 271938 233844
rect 463694 233832 463700 233844
rect 271932 233804 463700 233832
rect 271932 233792 271938 233804
rect 463694 233792 463700 233804
rect 463752 233792 463758 233844
rect 271414 233724 271420 233776
rect 271472 233764 271478 233776
rect 448606 233764 448612 233776
rect 271472 233736 448612 233764
rect 271472 233724 271478 233736
rect 448606 233724 448612 233736
rect 448664 233724 448670 233776
rect 271322 233656 271328 233708
rect 271380 233696 271386 233708
rect 445754 233696 445760 233708
rect 271380 233668 445760 233696
rect 271380 233656 271386 233668
rect 445754 233656 445760 233668
rect 445812 233656 445818 233708
rect 270862 232908 270868 232960
rect 270920 232948 270926 232960
rect 440326 232948 440332 232960
rect 270920 232920 440332 232948
rect 270920 232908 270926 232920
rect 440326 232908 440332 232920
rect 440384 232908 440390 232960
rect 271506 232840 271512 232892
rect 271564 232880 271570 232892
rect 442994 232880 443000 232892
rect 271564 232852 443000 232880
rect 271564 232840 271570 232852
rect 442994 232840 443000 232852
rect 443052 232840 443058 232892
rect 272058 232772 272064 232824
rect 272116 232812 272122 232824
rect 465166 232812 465172 232824
rect 272116 232784 465172 232812
rect 272116 232772 272122 232784
rect 465166 232772 465172 232784
rect 465224 232772 465230 232824
rect 277118 232704 277124 232756
rect 277176 232744 277182 232756
rect 510614 232744 510620 232756
rect 277176 232716 510620 232744
rect 277176 232704 277182 232716
rect 510614 232704 510620 232716
rect 510672 232704 510678 232756
rect 278314 232636 278320 232688
rect 278372 232676 278378 232688
rect 521654 232676 521660 232688
rect 278372 232648 521660 232676
rect 278372 232636 278378 232648
rect 521654 232636 521660 232648
rect 521712 232636 521718 232688
rect 278498 232568 278504 232620
rect 278556 232608 278562 232620
rect 524414 232608 524420 232620
rect 278556 232580 524420 232608
rect 278556 232568 278562 232580
rect 524414 232568 524420 232580
rect 524472 232568 524478 232620
rect 260098 232500 260104 232552
rect 260156 232540 260162 232552
rect 276014 232540 276020 232552
rect 260156 232512 276020 232540
rect 260156 232500 260162 232512
rect 276014 232500 276020 232512
rect 276072 232500 276078 232552
rect 278406 232500 278412 232552
rect 278464 232540 278470 232552
rect 528554 232540 528560 232552
rect 278464 232512 528560 232540
rect 278464 232500 278470 232512
rect 528554 232500 528560 232512
rect 528612 232500 528618 232552
rect 274910 231140 274916 231192
rect 274968 231180 274974 231192
rect 499574 231180 499580 231192
rect 274968 231152 499580 231180
rect 274968 231140 274974 231152
rect 499574 231140 499580 231152
rect 499632 231140 499638 231192
rect 276106 231072 276112 231124
rect 276164 231112 276170 231124
rect 514754 231112 514760 231124
rect 276164 231084 514760 231112
rect 276164 231072 276170 231084
rect 514754 231072 514760 231084
rect 514812 231072 514818 231124
rect 286502 219376 286508 219428
rect 286560 219416 286566 219428
rect 580166 219416 580172 219428
rect 286560 219388 580172 219416
rect 286560 219376 286566 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 32490 215268 32496 215280
rect 3384 215240 32496 215268
rect 3384 215228 3390 215240
rect 32490 215228 32496 215240
rect 32548 215228 32554 215280
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 39390 202824 39396 202836
rect 3108 202796 39396 202824
rect 3108 202784 3114 202796
rect 39390 202784 39396 202796
rect 39448 202784 39454 202836
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 21450 189020 21456 189032
rect 3568 188992 21456 189020
rect 3568 188980 3574 188992
rect 21450 188980 21456 188992
rect 21508 188980 21514 189032
rect 543090 179324 543096 179376
rect 543148 179364 543154 179376
rect 579614 179364 579620 179376
rect 543148 179336 579620 179364
rect 543148 179324 543154 179336
rect 579614 179324 579620 179336
rect 579672 179324 579678 179376
rect 271046 177352 271052 177404
rect 271104 177392 271110 177404
rect 447134 177392 447140 177404
rect 271104 177364 447140 177392
rect 271104 177352 271110 177364
rect 447134 177352 447140 177364
rect 447192 177352 447198 177404
rect 276290 177284 276296 177336
rect 276348 177324 276354 177336
rect 517514 177324 517520 177336
rect 276348 177296 517520 177324
rect 276348 177284 276354 177296
rect 517514 177284 517520 177296
rect 517572 177284 517578 177336
rect 277670 175924 277676 175976
rect 277728 175964 277734 175976
rect 530578 175964 530584 175976
rect 277728 175936 530584 175964
rect 277728 175924 277734 175936
rect 530578 175924 530584 175936
rect 530636 175924 530642 175976
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 14550 164200 14556 164212
rect 3292 164172 14556 164200
rect 3292 164160 3298 164172
rect 14550 164160 14556 164172
rect 14608 164160 14614 164212
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 40770 150396 40776 150408
rect 3568 150368 40776 150396
rect 3568 150356 3574 150368
rect 40770 150356 40776 150368
rect 40828 150356 40834 150408
rect 573358 139340 573364 139392
rect 573416 139380 573422 139392
rect 580166 139380 580172 139392
rect 573416 139352 580172 139380
rect 573416 139340 573422 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 29638 137952 29644 137964
rect 3568 137924 29644 137952
rect 3568 137912 3574 137924
rect 29638 137912 29644 137924
rect 29696 137912 29702 137964
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 11790 111772 11796 111784
rect 3200 111744 11796 111772
rect 3200 111732 3206 111744
rect 11790 111732 11796 111744
rect 11848 111732 11854 111784
rect 569310 100648 569316 100700
rect 569368 100688 569374 100700
rect 580166 100688 580172 100700
rect 569368 100660 580172 100688
rect 569368 100648 569374 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 33778 97968 33784 97980
rect 3568 97940 33784 97968
rect 3568 97928 3574 97940
rect 33778 97928 33784 97940
rect 33836 97928 33842 97980
rect 264514 93100 264520 93152
rect 264572 93140 264578 93152
rect 273254 93140 273260 93152
rect 264572 93112 273260 93140
rect 264572 93100 264578 93112
rect 273254 93100 273260 93112
rect 273312 93100 273318 93152
rect 313918 86912 313924 86964
rect 313976 86952 313982 86964
rect 580166 86952 580172 86964
rect 313976 86924 580172 86952
rect 313976 86912 313982 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 17218 85524 17224 85536
rect 3568 85496 17224 85524
rect 3568 85484 3574 85496
rect 17218 85484 17224 85496
rect 17276 85484 17282 85536
rect 302878 73108 302884 73160
rect 302936 73148 302942 73160
rect 580166 73148 580172 73160
rect 302936 73120 580172 73148
rect 302936 73108 302942 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 2774 71612 2780 71664
rect 2832 71652 2838 71664
rect 4798 71652 4804 71664
rect 2832 71624 4804 71652
rect 2832 71612 2838 71624
rect 4798 71612 4804 71624
rect 4856 71612 4862 71664
rect 555418 60664 555424 60716
rect 555476 60704 555482 60716
rect 580166 60704 580172 60716
rect 555476 60676 580172 60704
rect 555476 60664 555482 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 35158 59344 35164 59356
rect 3108 59316 35164 59344
rect 3108 59304 3114 59316
rect 35158 59304 35164 59316
rect 35216 59304 35222 59356
rect 295978 46860 295984 46912
rect 296036 46900 296042 46912
rect 580166 46900 580172 46912
rect 296036 46872 580172 46900
rect 296036 46860 296042 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 18598 45540 18604 45552
rect 3568 45512 18604 45540
rect 3568 45500 3574 45512
rect 18598 45500 18604 45512
rect 18656 45500 18662 45552
rect 300118 33056 300124 33108
rect 300176 33096 300182 33108
rect 580166 33096 580172 33108
rect 300176 33068 580172 33096
rect 300176 33056 300182 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 152458 20652 152464 20664
rect 3476 20624 152464 20652
rect 3476 20612 3482 20624
rect 152458 20612 152464 20624
rect 152516 20612 152522 20664
rect 540238 20612 540244 20664
rect 540296 20652 540302 20664
rect 579982 20652 579988 20664
rect 540296 20624 579988 20652
rect 540296 20612 540302 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 265710 18572 265716 18624
rect 265768 18612 265774 18624
rect 372614 18612 372620 18624
rect 265768 18584 372620 18612
rect 265768 18572 265774 18584
rect 372614 18572 372620 18584
rect 372672 18572 372678 18624
rect 51810 13064 51816 13116
rect 51868 13104 51874 13116
rect 238570 13104 238576 13116
rect 51868 13076 238576 13104
rect 51868 13064 51874 13076
rect 238570 13064 238576 13076
rect 238628 13064 238634 13116
rect 357526 11704 357532 11756
rect 357584 11744 357590 11756
rect 358722 11744 358728 11756
rect 357584 11716 358728 11744
rect 357584 11704 357590 11716
rect 358722 11704 358728 11716
rect 358780 11704 358786 11756
rect 374086 11704 374092 11756
rect 374144 11744 374150 11756
rect 375282 11744 375288 11756
rect 374144 11716 375288 11744
rect 374144 11704 374150 11716
rect 375282 11704 375288 11716
rect 375340 11704 375346 11756
rect 398926 11704 398932 11756
rect 398984 11744 398990 11756
rect 400122 11744 400128 11756
rect 398984 11716 400128 11744
rect 398984 11704 398990 11716
rect 400122 11704 400128 11716
rect 400180 11704 400186 11756
rect 448606 11704 448612 11756
rect 448664 11744 448670 11756
rect 449802 11744 449808 11756
rect 448664 11716 449808 11744
rect 448664 11704 448670 11716
rect 449802 11704 449808 11716
rect 449860 11704 449866 11756
rect 260466 10956 260472 11008
rect 260524 10996 260530 11008
rect 314654 10996 314660 11008
rect 260524 10968 314660 10996
rect 260524 10956 260530 10968
rect 314654 10956 314660 10968
rect 314712 10956 314718 11008
rect 261570 10888 261576 10940
rect 261628 10928 261634 10940
rect 317966 10928 317972 10940
rect 261628 10900 317972 10928
rect 261628 10888 261634 10900
rect 317966 10888 317972 10900
rect 318024 10888 318030 10940
rect 261754 10820 261760 10872
rect 261812 10860 261818 10872
rect 322106 10860 322112 10872
rect 261812 10832 322112 10860
rect 261812 10820 261818 10832
rect 322106 10820 322112 10832
rect 322164 10820 322170 10872
rect 261662 10752 261668 10804
rect 261720 10792 261726 10804
rect 324314 10792 324320 10804
rect 261720 10764 324320 10792
rect 261720 10752 261726 10764
rect 324314 10752 324320 10764
rect 324372 10752 324378 10804
rect 261846 10684 261852 10736
rect 261904 10724 261910 10736
rect 328730 10724 328736 10736
rect 261904 10696 328736 10724
rect 261904 10684 261910 10696
rect 328730 10684 328736 10696
rect 328788 10684 328794 10736
rect 261478 10616 261484 10668
rect 261536 10656 261542 10668
rect 332686 10656 332692 10668
rect 261536 10628 332692 10656
rect 261536 10616 261542 10628
rect 332686 10616 332692 10628
rect 332744 10616 332750 10668
rect 262766 10548 262772 10600
rect 262824 10588 262830 10600
rect 336274 10588 336280 10600
rect 262824 10560 336280 10588
rect 262824 10548 262830 10560
rect 336274 10548 336280 10560
rect 336332 10548 336338 10600
rect 262674 10480 262680 10532
rect 262732 10520 262738 10532
rect 339494 10520 339500 10532
rect 262732 10492 339500 10520
rect 262732 10480 262738 10492
rect 339494 10480 339500 10492
rect 339552 10480 339558 10532
rect 263042 10412 263048 10464
rect 263100 10452 263106 10464
rect 342898 10452 342904 10464
rect 263100 10424 342904 10452
rect 263100 10412 263106 10424
rect 342898 10412 342904 10424
rect 342956 10412 342962 10464
rect 262950 10344 262956 10396
rect 263008 10384 263014 10396
rect 346946 10384 346952 10396
rect 263008 10356 346952 10384
rect 263008 10344 263014 10356
rect 346946 10344 346952 10356
rect 347004 10344 347010 10396
rect 245102 10276 245108 10328
rect 245160 10316 245166 10328
rect 254486 10316 254492 10328
rect 245160 10288 254492 10316
rect 245160 10276 245166 10288
rect 254486 10276 254492 10288
rect 254544 10276 254550 10328
rect 262858 10276 262864 10328
rect 262916 10316 262922 10328
rect 349154 10316 349160 10328
rect 262916 10288 349160 10316
rect 262916 10276 262922 10288
rect 349154 10276 349160 10288
rect 349212 10276 349218 10328
rect 252646 9528 252652 9580
rect 252704 9568 252710 9580
rect 254302 9568 254308 9580
rect 252704 9540 254308 9568
rect 252704 9528 252710 9540
rect 254302 9528 254308 9540
rect 254360 9528 254366 9580
rect 253474 8440 253480 8492
rect 253532 8480 253538 8492
rect 255590 8480 255596 8492
rect 253532 8452 255596 8480
rect 253532 8440 253538 8452
rect 255590 8440 255596 8452
rect 255648 8440 255654 8492
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 21358 6848 21364 6860
rect 3476 6820 21364 6848
rect 3476 6808 3482 6820
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 318058 6808 318064 6860
rect 318116 6848 318122 6860
rect 580166 6848 580172 6860
rect 318116 6820 580172 6848
rect 318116 6808 318122 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 259546 6672 259552 6724
rect 259604 6712 259610 6724
rect 313826 6712 313832 6724
rect 259604 6684 313832 6712
rect 259604 6672 259610 6684
rect 313826 6672 313832 6684
rect 313884 6672 313890 6724
rect 262030 6604 262036 6656
rect 262088 6644 262094 6656
rect 324406 6644 324412 6656
rect 262088 6616 324412 6644
rect 262088 6604 262094 6616
rect 324406 6604 324412 6616
rect 324464 6604 324470 6656
rect 261938 6536 261944 6588
rect 261996 6576 262002 6588
rect 327994 6576 328000 6588
rect 261996 6548 328000 6576
rect 261996 6536 262002 6548
rect 327994 6536 328000 6548
rect 328052 6536 328058 6588
rect 262122 6468 262128 6520
rect 262180 6508 262186 6520
rect 331582 6508 331588 6520
rect 262180 6480 331588 6508
rect 262180 6468 262186 6480
rect 331582 6468 331588 6480
rect 331640 6468 331646 6520
rect 263134 6400 263140 6452
rect 263192 6440 263198 6452
rect 335078 6440 335084 6452
rect 263192 6412 335084 6440
rect 263192 6400 263198 6412
rect 335078 6400 335084 6412
rect 335136 6400 335142 6452
rect 263226 6332 263232 6384
rect 263284 6372 263290 6384
rect 338666 6372 338672 6384
rect 263284 6344 338672 6372
rect 263284 6332 263290 6344
rect 338666 6332 338672 6344
rect 338724 6332 338730 6384
rect 263318 6264 263324 6316
rect 263376 6304 263382 6316
rect 342162 6304 342168 6316
rect 263376 6276 342168 6304
rect 263376 6264 263382 6276
rect 342162 6264 342168 6276
rect 342220 6264 342226 6316
rect 262398 6196 262404 6248
rect 262456 6236 262462 6248
rect 345750 6236 345756 6248
rect 262456 6208 345756 6236
rect 262456 6196 262462 6208
rect 345750 6196 345756 6208
rect 345808 6196 345814 6248
rect 74994 6128 75000 6180
rect 75052 6168 75058 6180
rect 240686 6168 240692 6180
rect 75052 6140 240692 6168
rect 75052 6128 75058 6140
rect 240686 6128 240692 6140
rect 240744 6128 240750 6180
rect 262214 6128 262220 6180
rect 262272 6168 262278 6180
rect 349246 6168 349252 6180
rect 262272 6140 349252 6168
rect 262272 6128 262278 6140
rect 349246 6128 349252 6140
rect 349304 6128 349310 6180
rect 257062 5448 257068 5500
rect 257120 5488 257126 5500
rect 272429 5491 272487 5497
rect 272429 5488 272441 5491
rect 257120 5460 272441 5488
rect 257120 5448 257126 5460
rect 272429 5457 272441 5460
rect 272475 5457 272487 5491
rect 272429 5451 272487 5457
rect 272521 5491 272579 5497
rect 272521 5457 272533 5491
rect 272567 5488 272579 5491
rect 278314 5488 278320 5500
rect 272567 5460 278320 5488
rect 272567 5457 272579 5460
rect 272521 5451 272579 5457
rect 278314 5448 278320 5460
rect 278372 5448 278378 5500
rect 286410 5448 286416 5500
rect 286468 5488 286474 5500
rect 411898 5488 411904 5500
rect 286468 5460 411904 5488
rect 286468 5448 286474 5460
rect 411898 5448 411904 5460
rect 411956 5448 411962 5500
rect 269298 5380 269304 5432
rect 269356 5420 269362 5432
rect 424962 5420 424968 5432
rect 269356 5392 424968 5420
rect 269356 5380 269362 5392
rect 424962 5380 424968 5392
rect 425020 5380 425026 5432
rect 256326 5312 256332 5364
rect 256384 5352 256390 5364
rect 264146 5352 264152 5364
rect 256384 5324 264152 5352
rect 256384 5312 256390 5324
rect 264146 5312 264152 5324
rect 264204 5312 264210 5364
rect 269666 5312 269672 5364
rect 269724 5352 269730 5364
rect 429654 5352 429660 5364
rect 269724 5324 429660 5352
rect 269724 5312 269730 5324
rect 429654 5312 429660 5324
rect 429712 5312 429718 5364
rect 257798 5244 257804 5296
rect 257856 5284 257862 5296
rect 268838 5284 268844 5296
rect 257856 5256 268844 5284
rect 257856 5244 257862 5256
rect 268838 5244 268844 5256
rect 268896 5244 268902 5296
rect 270218 5244 270224 5296
rect 270276 5284 270282 5296
rect 432046 5284 432052 5296
rect 270276 5256 432052 5284
rect 270276 5244 270282 5256
rect 432046 5244 432052 5256
rect 432104 5244 432110 5296
rect 257430 5176 257436 5228
rect 257488 5216 257494 5228
rect 272521 5219 272579 5225
rect 272521 5216 272533 5219
rect 257488 5188 272533 5216
rect 257488 5176 257494 5188
rect 272521 5185 272533 5188
rect 272567 5185 272579 5219
rect 272521 5179 272579 5185
rect 284938 5176 284944 5228
rect 284996 5216 285002 5228
rect 454494 5216 454500 5228
rect 284996 5188 454500 5216
rect 284996 5176 285002 5188
rect 454494 5176 454500 5188
rect 454552 5176 454558 5228
rect 234614 5108 234620 5160
rect 234672 5148 234678 5160
rect 249058 5148 249064 5160
rect 234672 5120 249064 5148
rect 234672 5108 234678 5120
rect 249058 5108 249064 5120
rect 249116 5108 249122 5160
rect 257614 5108 257620 5160
rect 257672 5148 257678 5160
rect 270586 5148 270592 5160
rect 257672 5120 270592 5148
rect 257672 5108 257678 5120
rect 270586 5108 270592 5120
rect 270644 5108 270650 5160
rect 270678 5108 270684 5160
rect 270736 5148 270742 5160
rect 450906 5148 450912 5160
rect 270736 5120 450912 5148
rect 270736 5108 270742 5120
rect 450906 5108 450912 5120
rect 450964 5108 450970 5160
rect 209774 5040 209780 5092
rect 209832 5080 209838 5092
rect 251634 5080 251640 5092
rect 209832 5052 251640 5080
rect 209832 5040 209838 5052
rect 251634 5040 251640 5052
rect 251692 5040 251698 5092
rect 257246 5040 257252 5092
rect 257304 5080 257310 5092
rect 281902 5080 281908 5092
rect 257304 5052 281908 5080
rect 257304 5040 257310 5052
rect 281902 5040 281908 5052
rect 281960 5040 281966 5092
rect 286318 5040 286324 5092
rect 286376 5080 286382 5092
rect 468662 5080 468668 5092
rect 286376 5052 468668 5080
rect 286376 5040 286382 5052
rect 468662 5040 468668 5052
rect 468720 5040 468726 5092
rect 181438 4972 181444 5024
rect 181496 5012 181502 5024
rect 248782 5012 248788 5024
rect 181496 4984 248788 5012
rect 181496 4972 181502 4984
rect 248782 4972 248788 4984
rect 248840 4972 248846 5024
rect 257706 4972 257712 5024
rect 257764 5012 257770 5024
rect 272426 5012 272432 5024
rect 257764 4984 272432 5012
rect 257764 4972 257770 4984
rect 272426 4972 272432 4984
rect 272484 4972 272490 5024
rect 273898 4972 273904 5024
rect 273956 5012 273962 5024
rect 455690 5012 455696 5024
rect 273956 4984 455696 5012
rect 273956 4972 273962 4984
rect 455690 4972 455696 4984
rect 455748 4972 455754 5024
rect 145926 4904 145932 4956
rect 145984 4944 145990 4956
rect 246666 4944 246672 4956
rect 145984 4916 246672 4944
rect 145984 4904 145990 4916
rect 246666 4904 246672 4916
rect 246724 4904 246730 4956
rect 257890 4904 257896 4956
rect 257948 4944 257954 4956
rect 279510 4944 279516 4956
rect 257948 4916 279516 4944
rect 257948 4904 257954 4916
rect 279510 4904 279516 4916
rect 279568 4904 279574 4956
rect 279602 4904 279608 4956
rect 279660 4944 279666 4956
rect 486418 4944 486424 4956
rect 279660 4916 486424 4944
rect 279660 4904 279666 4916
rect 486418 4904 486424 4916
rect 486476 4904 486482 4956
rect 135254 4836 135260 4888
rect 135312 4876 135318 4888
rect 246206 4876 246212 4888
rect 135312 4848 246212 4876
rect 135312 4836 135318 4848
rect 246206 4836 246212 4848
rect 246264 4836 246270 4888
rect 257338 4836 257344 4888
rect 257396 4876 257402 4888
rect 267734 4876 267740 4888
rect 257396 4848 267740 4876
rect 257396 4836 257402 4848
rect 267734 4836 267740 4848
rect 267792 4836 267798 4888
rect 272429 4879 272487 4885
rect 272429 4845 272441 4879
rect 272475 4876 272487 4879
rect 276014 4876 276020 4888
rect 272475 4848 276020 4876
rect 272475 4845 272487 4848
rect 272429 4839 272487 4845
rect 276014 4836 276020 4848
rect 276072 4836 276078 4888
rect 276109 4879 276167 4885
rect 276109 4845 276121 4879
rect 276155 4876 276167 4879
rect 301958 4876 301964 4888
rect 276155 4848 301964 4876
rect 276155 4845 276167 4848
rect 276109 4839 276167 4845
rect 301958 4836 301964 4848
rect 302016 4836 302022 4888
rect 304258 4836 304264 4888
rect 304316 4876 304322 4888
rect 582190 4876 582196 4888
rect 304316 4848 582196 4876
rect 304316 4836 304322 4848
rect 582190 4836 582196 4848
rect 582248 4836 582254 4888
rect 67910 4768 67916 4820
rect 67968 4808 67974 4820
rect 240594 4808 240600 4820
rect 67968 4780 240600 4808
rect 67968 4768 67974 4780
rect 240594 4768 240600 4780
rect 240652 4768 240658 4820
rect 258626 4768 258632 4820
rect 258684 4808 258690 4820
rect 297266 4808 297272 4820
rect 258684 4780 297272 4808
rect 258684 4768 258690 4780
rect 297266 4768 297272 4780
rect 297324 4768 297330 4820
rect 299566 4768 299572 4820
rect 299624 4808 299630 4820
rect 300762 4808 300768 4820
rect 299624 4780 300768 4808
rect 299624 4768 299630 4780
rect 300762 4768 300768 4780
rect 300820 4768 300826 4820
rect 304442 4768 304448 4820
rect 304500 4808 304506 4820
rect 583389 4811 583447 4817
rect 583389 4808 583401 4811
rect 304500 4780 583401 4808
rect 304500 4768 304506 4780
rect 583389 4777 583401 4780
rect 583435 4777 583447 4811
rect 583389 4771 583447 4777
rect 265802 4700 265808 4752
rect 265860 4740 265866 4752
rect 379974 4740 379980 4752
rect 265860 4712 379980 4740
rect 265860 4700 265866 4712
rect 379974 4700 379980 4712
rect 380032 4700 380038 4752
rect 268378 4632 268384 4684
rect 268436 4672 268442 4684
rect 276109 4675 276167 4681
rect 276109 4672 276121 4675
rect 268436 4644 276121 4672
rect 268436 4632 268442 4644
rect 276109 4641 276121 4644
rect 276155 4641 276167 4675
rect 276109 4635 276167 4641
rect 276201 4675 276259 4681
rect 276201 4641 276213 4675
rect 276247 4672 276259 4675
rect 276247 4644 354674 4672
rect 276247 4641 276259 4644
rect 276201 4635 276259 4641
rect 269850 4564 269856 4616
rect 269908 4604 269914 4616
rect 351638 4604 351644 4616
rect 269908 4576 351644 4604
rect 269908 4564 269914 4576
rect 351638 4564 351644 4576
rect 351696 4564 351702 4616
rect 354646 4604 354674 4644
rect 365806 4604 365812 4616
rect 354646 4576 365812 4604
rect 365806 4564 365812 4576
rect 365864 4564 365870 4616
rect 264238 4496 264244 4548
rect 264296 4536 264302 4548
rect 264296 4508 316034 4536
rect 264296 4496 264302 4508
rect 260006 4428 260012 4480
rect 260064 4468 260070 4480
rect 312630 4468 312636 4480
rect 260064 4440 312636 4468
rect 260064 4428 260070 4440
rect 312630 4428 312636 4440
rect 312688 4428 312694 4480
rect 316006 4468 316034 4508
rect 326798 4468 326804 4480
rect 316006 4440 326804 4468
rect 326798 4428 326804 4440
rect 326856 4428 326862 4480
rect 257522 4360 257528 4412
rect 257580 4400 257586 4412
rect 274818 4400 274824 4412
rect 257580 4372 274824 4400
rect 257580 4360 257586 4372
rect 274818 4360 274824 4372
rect 274876 4360 274882 4412
rect 285030 4360 285036 4412
rect 285088 4400 285094 4412
rect 333882 4400 333888 4412
rect 285088 4372 333888 4400
rect 285088 4360 285094 4372
rect 333882 4360 333888 4372
rect 333940 4360 333946 4412
rect 259914 4292 259920 4344
rect 259972 4332 259978 4344
rect 307938 4332 307944 4344
rect 259972 4304 307944 4332
rect 259972 4292 259978 4304
rect 307938 4292 307944 4304
rect 307996 4292 308002 4344
rect 269942 4224 269948 4276
rect 270000 4264 270006 4276
rect 309042 4264 309048 4276
rect 270000 4236 309048 4264
rect 270000 4224 270006 4236
rect 309042 4224 309048 4236
rect 309100 4224 309106 4276
rect 268470 4156 268476 4208
rect 268528 4196 268534 4208
rect 268528 4168 270540 4196
rect 268528 4156 268534 4168
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 22738 4128 22744 4140
rect 13596 4100 22744 4128
rect 13596 4088 13602 4100
rect 22738 4088 22744 4100
rect 22796 4088 22802 4140
rect 27706 4088 27712 4140
rect 27764 4128 27770 4140
rect 51718 4128 51724 4140
rect 27764 4100 51724 4128
rect 27764 4088 27770 4100
rect 51718 4088 51724 4100
rect 51776 4088 51782 4140
rect 99834 4088 99840 4140
rect 99892 4128 99898 4140
rect 233881 4131 233939 4137
rect 233881 4128 233893 4131
rect 99892 4100 233893 4128
rect 99892 4088 99898 4100
rect 233881 4097 233893 4100
rect 233927 4097 233939 4131
rect 233881 4091 233939 4097
rect 247586 4088 247592 4140
rect 247644 4128 247650 4140
rect 251174 4128 251180 4140
rect 247644 4100 251180 4128
rect 247644 4088 247650 4100
rect 251174 4088 251180 4100
rect 251232 4088 251238 4140
rect 270512 4128 270540 4168
rect 270586 4156 270592 4208
rect 270644 4196 270650 4208
rect 271230 4196 271236 4208
rect 270644 4168 271236 4196
rect 270644 4156 270650 4168
rect 271230 4156 271236 4168
rect 271288 4156 271294 4208
rect 276201 4199 276259 4205
rect 276201 4196 276213 4199
rect 271340 4168 276213 4196
rect 271340 4128 271368 4168
rect 276201 4165 276213 4168
rect 276247 4165 276259 4199
rect 276201 4159 276259 4165
rect 285122 4156 285128 4208
rect 285180 4196 285186 4208
rect 319714 4196 319720 4208
rect 285180 4168 319720 4196
rect 285180 4156 285186 4168
rect 319714 4156 319720 4168
rect 319772 4156 319778 4208
rect 324314 4156 324320 4208
rect 324372 4196 324378 4208
rect 325602 4196 325608 4208
rect 324372 4168 325608 4196
rect 324372 4156 324378 4168
rect 325602 4156 325608 4168
rect 325660 4156 325666 4208
rect 270512 4100 271368 4128
rect 279694 4088 279700 4140
rect 279752 4128 279758 4140
rect 475746 4128 475752 4140
rect 279752 4100 475752 4128
rect 279752 4088 279758 4100
rect 475746 4088 475752 4100
rect 475804 4088 475810 4140
rect 483658 4088 483664 4140
rect 483716 4128 483722 4140
rect 492306 4128 492312 4140
rect 483716 4100 492312 4128
rect 483716 4088 483722 4100
rect 492306 4088 492312 4100
rect 492364 4088 492370 4140
rect 547138 4088 547144 4140
rect 547196 4128 547202 4140
rect 549070 4128 549076 4140
rect 547196 4100 549076 4128
rect 547196 4088 547202 4100
rect 549070 4088 549076 4100
rect 549128 4088 549134 4140
rect 566458 4088 566464 4140
rect 566516 4128 566522 4140
rect 568022 4128 568028 4140
rect 566516 4100 568028 4128
rect 566516 4088 566522 4100
rect 568022 4088 568028 4100
rect 568080 4088 568086 4140
rect 566 4020 572 4072
rect 624 4060 630 4072
rect 32306 4060 32312 4072
rect 624 4032 32312 4060
rect 624 4020 630 4032
rect 32306 4020 32312 4032
rect 32364 4020 32370 4072
rect 34790 4020 34796 4072
rect 34848 4060 34854 4072
rect 58618 4060 58624 4072
rect 34848 4032 58624 4060
rect 34848 4020 34854 4032
rect 58618 4020 58624 4032
rect 58676 4020 58682 4072
rect 92750 4020 92756 4072
rect 92808 4060 92814 4072
rect 242066 4060 242072 4072
rect 92808 4032 242072 4060
rect 92808 4020 92814 4032
rect 242066 4020 242072 4032
rect 242124 4020 242130 4072
rect 257062 4020 257068 4072
rect 257120 4060 257126 4072
rect 259454 4060 259460 4072
rect 257120 4032 259460 4060
rect 257120 4020 257126 4032
rect 259454 4020 259460 4032
rect 259512 4020 259518 4072
rect 280798 4020 280804 4072
rect 280856 4060 280862 4072
rect 478233 4063 478291 4069
rect 478233 4060 478245 4063
rect 280856 4032 478245 4060
rect 280856 4020 280862 4032
rect 478233 4029 478245 4032
rect 478279 4029 478291 4063
rect 478233 4023 478291 4029
rect 544378 4020 544384 4072
rect 544436 4060 544442 4072
rect 550266 4060 550272 4072
rect 544436 4032 550272 4060
rect 544436 4020 544442 4032
rect 550266 4020 550272 4032
rect 550324 4020 550330 4072
rect 1670 3952 1676 4004
rect 1728 3992 1734 4004
rect 36538 3992 36544 4004
rect 1728 3964 36544 3992
rect 1728 3952 1734 3964
rect 36538 3952 36544 3964
rect 36596 3952 36602 4004
rect 44266 3952 44272 4004
rect 44324 3992 44330 4004
rect 46198 3992 46204 4004
rect 44324 3964 46204 3992
rect 44324 3952 44330 3964
rect 46198 3952 46204 3964
rect 46256 3952 46262 4004
rect 85666 3952 85672 4004
rect 85724 3992 85730 4004
rect 241974 3992 241980 4004
rect 85724 3964 241980 3992
rect 85724 3952 85730 3964
rect 241974 3952 241980 3964
rect 242032 3952 242038 4004
rect 245194 3952 245200 4004
rect 245252 3992 245258 4004
rect 251910 3992 251916 4004
rect 245252 3964 251916 3992
rect 245252 3952 245258 3964
rect 251910 3952 251916 3964
rect 251968 3952 251974 4004
rect 287974 3952 287980 4004
rect 288032 3992 288038 4004
rect 491110 3992 491116 4004
rect 288032 3964 491116 3992
rect 288032 3952 288038 3964
rect 491110 3952 491116 3964
rect 491168 3952 491174 4004
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 173069 3927 173127 3933
rect 173069 3924 173081 3927
rect 20680 3896 173081 3924
rect 20680 3884 20686 3896
rect 173069 3893 173081 3896
rect 173115 3893 173127 3927
rect 173069 3887 173127 3893
rect 173158 3884 173164 3936
rect 173216 3924 173222 3936
rect 173710 3924 173716 3936
rect 173216 3896 173716 3924
rect 173216 3884 173222 3896
rect 173710 3884 173716 3896
rect 173768 3884 173774 3936
rect 174262 3884 174268 3936
rect 174320 3924 174326 3936
rect 175182 3924 175188 3936
rect 174320 3896 175188 3924
rect 174320 3884 174326 3896
rect 175182 3884 175188 3896
rect 175240 3884 175246 3936
rect 175458 3884 175464 3936
rect 175516 3924 175522 3936
rect 176562 3924 176568 3936
rect 175516 3896 176568 3924
rect 175516 3884 175522 3896
rect 176562 3884 176568 3896
rect 176620 3884 176626 3936
rect 176654 3884 176660 3936
rect 176712 3924 176718 3936
rect 177942 3924 177948 3936
rect 176712 3896 177948 3924
rect 176712 3884 176718 3896
rect 177942 3884 177948 3896
rect 178000 3884 178006 3936
rect 180242 3884 180248 3936
rect 180300 3924 180306 3936
rect 180702 3924 180708 3936
rect 180300 3896 180708 3924
rect 180300 3884 180306 3896
rect 180702 3884 180708 3896
rect 180760 3884 180766 3936
rect 182542 3884 182548 3936
rect 182600 3924 182606 3936
rect 183462 3924 183468 3936
rect 182600 3896 183468 3924
rect 182600 3884 182606 3896
rect 183462 3884 183468 3896
rect 183520 3884 183526 3936
rect 183738 3884 183744 3936
rect 183796 3924 183802 3936
rect 184842 3924 184848 3936
rect 183796 3896 184848 3924
rect 183796 3884 183802 3896
rect 184842 3884 184848 3896
rect 184900 3884 184906 3936
rect 184934 3884 184940 3936
rect 184992 3924 184998 3936
rect 186038 3924 186044 3936
rect 184992 3896 186044 3924
rect 184992 3884 184998 3896
rect 186038 3884 186044 3896
rect 186096 3884 186102 3936
rect 188522 3884 188528 3936
rect 188580 3924 188586 3936
rect 188982 3924 188988 3936
rect 188580 3896 188988 3924
rect 188580 3884 188586 3896
rect 188982 3884 188988 3896
rect 189040 3884 189046 3936
rect 189718 3884 189724 3936
rect 189776 3924 189782 3936
rect 190362 3924 190368 3936
rect 189776 3896 190368 3924
rect 189776 3884 189782 3896
rect 190362 3884 190368 3896
rect 190420 3884 190426 3936
rect 190822 3884 190828 3936
rect 190880 3924 190886 3936
rect 191742 3924 191748 3936
rect 190880 3896 191748 3924
rect 190880 3884 190886 3896
rect 191742 3884 191748 3896
rect 191800 3884 191806 3936
rect 192018 3884 192024 3936
rect 192076 3924 192082 3936
rect 193122 3924 193128 3936
rect 192076 3896 193128 3924
rect 192076 3884 192082 3896
rect 193122 3884 193128 3896
rect 193180 3884 193186 3936
rect 193214 3884 193220 3936
rect 193272 3924 193278 3936
rect 194502 3924 194508 3936
rect 193272 3896 194508 3924
rect 193272 3884 193278 3896
rect 194502 3884 194508 3896
rect 194560 3884 194566 3936
rect 196802 3884 196808 3936
rect 196860 3924 196866 3936
rect 197262 3924 197268 3936
rect 196860 3896 197268 3924
rect 196860 3884 196866 3896
rect 197262 3884 197268 3896
rect 197320 3884 197326 3936
rect 199102 3884 199108 3936
rect 199160 3924 199166 3936
rect 200022 3924 200028 3936
rect 199160 3896 200028 3924
rect 199160 3884 199166 3896
rect 200022 3884 200028 3896
rect 200080 3884 200086 3936
rect 200298 3884 200304 3936
rect 200356 3924 200362 3936
rect 201402 3924 201408 3936
rect 200356 3896 201408 3924
rect 200356 3884 200362 3896
rect 201402 3884 201408 3896
rect 201460 3884 201466 3936
rect 201494 3884 201500 3936
rect 201552 3924 201558 3936
rect 202782 3924 202788 3936
rect 201552 3896 202788 3924
rect 201552 3884 201558 3896
rect 202782 3884 202788 3896
rect 202840 3884 202846 3936
rect 205082 3884 205088 3936
rect 205140 3924 205146 3936
rect 205542 3924 205548 3936
rect 205140 3896 205548 3924
rect 205140 3884 205146 3896
rect 205542 3884 205548 3896
rect 205600 3884 205606 3936
rect 206186 3884 206192 3936
rect 206244 3924 206250 3936
rect 206922 3924 206928 3936
rect 206244 3896 206928 3924
rect 206244 3884 206250 3896
rect 206922 3884 206928 3896
rect 206980 3884 206986 3936
rect 207382 3884 207388 3936
rect 207440 3924 207446 3936
rect 208302 3924 208308 3936
rect 207440 3896 208308 3924
rect 207440 3884 207446 3896
rect 208302 3884 208308 3896
rect 208360 3884 208366 3936
rect 208397 3927 208455 3933
rect 208397 3893 208409 3927
rect 208443 3924 208455 3927
rect 250162 3924 250168 3936
rect 208443 3896 250168 3924
rect 208443 3893 208455 3896
rect 208397 3887 208455 3893
rect 250162 3884 250168 3896
rect 250220 3884 250226 3936
rect 280982 3884 280988 3936
rect 281040 3924 281046 3936
rect 484026 3924 484032 3936
rect 281040 3896 484032 3924
rect 281040 3884 281046 3896
rect 484026 3884 484032 3896
rect 484084 3884 484090 3936
rect 497458 3884 497464 3936
rect 497516 3924 497522 3936
rect 510062 3924 510068 3936
rect 497516 3896 510068 3924
rect 497516 3884 497522 3896
rect 510062 3884 510068 3896
rect 510120 3884 510126 3936
rect 2866 3816 2872 3868
rect 2924 3856 2930 3868
rect 39298 3856 39304 3868
rect 2924 3828 39304 3856
rect 2924 3816 2930 3828
rect 39298 3816 39304 3828
rect 39356 3816 39362 3868
rect 43438 3856 43444 3868
rect 39684 3828 43444 3856
rect 7650 3748 7656 3800
rect 7708 3788 7714 3800
rect 39684 3788 39712 3828
rect 43438 3816 43444 3828
rect 43496 3816 43502 3868
rect 51810 3856 51816 3868
rect 45526 3828 51816 3856
rect 7708 3760 39712 3788
rect 7708 3748 7714 3760
rect 43070 3748 43076 3800
rect 43128 3788 43134 3800
rect 45526 3788 45554 3828
rect 51810 3816 51816 3828
rect 51868 3816 51874 3868
rect 69106 3816 69112 3868
rect 69164 3856 69170 3868
rect 70210 3856 70216 3868
rect 69164 3828 70216 3856
rect 69164 3816 69170 3828
rect 70210 3816 70216 3828
rect 70268 3816 70274 3868
rect 71498 3816 71504 3868
rect 71556 3856 71562 3868
rect 227717 3859 227775 3865
rect 227717 3856 227729 3859
rect 71556 3828 227729 3856
rect 71556 3816 71562 3828
rect 227717 3825 227729 3828
rect 227763 3825 227775 3859
rect 227717 3819 227775 3825
rect 235810 3816 235816 3868
rect 235868 3856 235874 3868
rect 245010 3856 245016 3868
rect 235868 3828 245016 3856
rect 235868 3816 235874 3828
rect 245010 3816 245016 3828
rect 245068 3816 245074 3868
rect 246390 3816 246396 3868
rect 246448 3856 246454 3868
rect 252646 3856 252652 3868
rect 246448 3828 252652 3856
rect 246448 3816 246454 3828
rect 252646 3816 252652 3828
rect 252704 3816 252710 3868
rect 280890 3816 280896 3868
rect 280948 3856 280954 3868
rect 487614 3856 487620 3868
rect 280948 3828 487620 3856
rect 280948 3816 280954 3828
rect 487614 3816 487620 3828
rect 487672 3816 487678 3868
rect 500310 3816 500316 3868
rect 500368 3856 500374 3868
rect 500368 3828 502104 3856
rect 500368 3816 500374 3828
rect 50430 3788 50436 3800
rect 43128 3760 45554 3788
rect 47964 3760 50436 3788
rect 43128 3748 43134 3760
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 47964 3720 47992 3760
rect 50430 3748 50436 3760
rect 50488 3748 50494 3800
rect 60826 3748 60832 3800
rect 60884 3788 60890 3800
rect 233881 3791 233939 3797
rect 60884 3760 233556 3788
rect 60884 3748 60890 3760
rect 11204 3692 47992 3720
rect 11204 3680 11210 3692
rect 50154 3680 50160 3732
rect 50212 3720 50218 3732
rect 50982 3720 50988 3732
rect 50212 3692 50988 3720
rect 50212 3680 50218 3692
rect 50982 3680 50988 3692
rect 51040 3680 51046 3732
rect 51350 3680 51356 3732
rect 51408 3720 51414 3732
rect 53098 3720 53104 3732
rect 51408 3692 53104 3720
rect 51408 3680 51414 3692
rect 53098 3680 53104 3692
rect 53156 3680 53162 3732
rect 53650 3680 53656 3732
rect 53708 3720 53714 3732
rect 233528 3720 233556 3760
rect 233881 3757 233893 3791
rect 233927 3788 233939 3791
rect 239398 3788 239404 3800
rect 233927 3760 239404 3788
rect 233927 3757 233939 3760
rect 233881 3751 233939 3757
rect 239398 3748 239404 3760
rect 239456 3748 239462 3800
rect 241698 3748 241704 3800
rect 241756 3788 241762 3800
rect 250438 3788 250444 3800
rect 241756 3760 250444 3788
rect 241756 3748 241762 3760
rect 250438 3748 250444 3760
rect 250496 3748 250502 3800
rect 287698 3748 287704 3800
rect 287756 3788 287762 3800
rect 494698 3788 494704 3800
rect 287756 3760 494704 3788
rect 287756 3748 287762 3760
rect 494698 3748 494704 3760
rect 494756 3748 494762 3800
rect 238018 3720 238024 3732
rect 53708 3692 233464 3720
rect 233528 3692 238024 3720
rect 53708 3680 53714 3692
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 26878 3652 26884 3664
rect 10008 3624 26884 3652
rect 10008 3612 10014 3624
rect 26878 3612 26884 3624
rect 26936 3612 26942 3664
rect 28902 3612 28908 3664
rect 28960 3652 28966 3664
rect 212813 3655 212871 3661
rect 212813 3652 212825 3655
rect 28960 3624 212825 3652
rect 28960 3612 28966 3624
rect 212813 3621 212825 3624
rect 212859 3621 212871 3655
rect 212813 3615 212871 3621
rect 213362 3612 213368 3664
rect 213420 3652 213426 3664
rect 213822 3652 213828 3664
rect 213420 3624 213828 3652
rect 213420 3612 213426 3624
rect 213822 3612 213828 3624
rect 213880 3612 213886 3664
rect 214466 3612 214472 3664
rect 214524 3652 214530 3664
rect 215202 3652 215208 3664
rect 214524 3624 215208 3652
rect 214524 3612 214530 3624
rect 215202 3612 215208 3624
rect 215260 3612 215266 3664
rect 215662 3612 215668 3664
rect 215720 3652 215726 3664
rect 216582 3652 216588 3664
rect 215720 3624 216588 3652
rect 215720 3612 215726 3624
rect 216582 3612 216588 3624
rect 216640 3612 216646 3664
rect 216858 3612 216864 3664
rect 216916 3652 216922 3664
rect 217962 3652 217968 3664
rect 216916 3624 217968 3652
rect 216916 3612 216922 3624
rect 217962 3612 217968 3624
rect 218020 3612 218026 3664
rect 218054 3612 218060 3664
rect 218112 3652 218118 3664
rect 219342 3652 219348 3664
rect 218112 3624 219348 3652
rect 218112 3612 218118 3624
rect 219342 3612 219348 3624
rect 219400 3612 219406 3664
rect 221550 3612 221556 3664
rect 221608 3652 221614 3664
rect 222102 3652 222108 3664
rect 221608 3624 222108 3652
rect 221608 3612 221614 3624
rect 222102 3612 222108 3624
rect 222160 3612 222166 3664
rect 222746 3612 222752 3664
rect 222804 3652 222810 3664
rect 223482 3652 223488 3664
rect 222804 3624 223488 3652
rect 222804 3612 222810 3624
rect 223482 3612 223488 3624
rect 223540 3612 223546 3664
rect 223942 3612 223948 3664
rect 224000 3652 224006 3664
rect 224862 3652 224868 3664
rect 224000 3624 224868 3652
rect 224000 3612 224006 3624
rect 224862 3612 224868 3624
rect 224920 3612 224926 3664
rect 225138 3612 225144 3664
rect 225196 3652 225202 3664
rect 226242 3652 226248 3664
rect 225196 3624 226248 3652
rect 225196 3612 225202 3624
rect 226242 3612 226248 3624
rect 226300 3612 226306 3664
rect 226334 3612 226340 3664
rect 226392 3652 226398 3664
rect 227622 3652 227628 3664
rect 226392 3624 227628 3652
rect 226392 3612 226398 3624
rect 227622 3612 227628 3624
rect 227680 3612 227686 3664
rect 227717 3655 227775 3661
rect 227717 3621 227729 3655
rect 227763 3652 227775 3655
rect 231210 3652 231216 3664
rect 227763 3624 231216 3652
rect 227763 3621 227775 3624
rect 227717 3615 227775 3621
rect 231210 3612 231216 3624
rect 231268 3612 231274 3664
rect 233436 3652 233464 3692
rect 238018 3680 238024 3692
rect 238076 3680 238082 3732
rect 244090 3680 244096 3732
rect 244148 3720 244154 3732
rect 253198 3720 253204 3732
rect 244148 3692 253204 3720
rect 244148 3680 244154 3692
rect 253198 3680 253204 3692
rect 253256 3680 253262 3732
rect 287882 3680 287888 3732
rect 287940 3720 287946 3732
rect 498194 3720 498200 3732
rect 287940 3692 498200 3720
rect 287940 3680 287946 3692
rect 498194 3680 498200 3692
rect 498252 3680 498258 3732
rect 501598 3680 501604 3732
rect 501656 3720 501662 3732
rect 502076 3720 502104 3828
rect 576118 3748 576124 3800
rect 576176 3788 576182 3800
rect 578602 3788 578608 3800
rect 576176 3760 578608 3788
rect 576176 3748 576182 3760
rect 578602 3748 578608 3760
rect 578660 3748 578666 3800
rect 513558 3720 513564 3732
rect 501656 3692 501920 3720
rect 502076 3692 513564 3720
rect 501656 3680 501662 3692
rect 238110 3652 238116 3664
rect 233436 3624 238116 3652
rect 238110 3612 238116 3624
rect 238168 3612 238174 3664
rect 240502 3612 240508 3664
rect 240560 3652 240566 3664
rect 249978 3652 249984 3664
rect 240560 3624 249984 3652
rect 240560 3612 240566 3624
rect 249978 3612 249984 3624
rect 250036 3612 250042 3664
rect 287790 3612 287796 3664
rect 287848 3652 287854 3664
rect 501782 3652 501788 3664
rect 287848 3624 501788 3652
rect 287848 3612 287854 3624
rect 501782 3612 501788 3624
rect 501840 3612 501846 3664
rect 501892 3652 501920 3692
rect 513558 3680 513564 3692
rect 513616 3680 513622 3732
rect 517146 3652 517152 3664
rect 501892 3624 517152 3652
rect 517146 3612 517152 3624
rect 517204 3612 517210 3664
rect 551278 3612 551284 3664
rect 551336 3652 551342 3664
rect 559742 3652 559748 3664
rect 551336 3624 559748 3652
rect 551336 3612 551342 3624
rect 559742 3612 559748 3624
rect 559800 3612 559806 3664
rect 23014 3544 23020 3596
rect 23072 3584 23078 3596
rect 231118 3584 231124 3596
rect 23072 3556 231124 3584
rect 23072 3544 23078 3556
rect 231118 3544 231124 3556
rect 231176 3544 231182 3596
rect 239306 3544 239312 3596
rect 239364 3584 239370 3596
rect 250530 3584 250536 3596
rect 239364 3556 250536 3584
rect 239364 3544 239370 3556
rect 250530 3544 250536 3556
rect 250588 3544 250594 3596
rect 256418 3544 256424 3596
rect 256476 3584 256482 3596
rect 260650 3584 260656 3596
rect 256476 3556 260656 3584
rect 256476 3544 256482 3556
rect 260650 3544 260656 3556
rect 260708 3544 260714 3596
rect 284294 3544 284300 3596
rect 284352 3584 284358 3596
rect 285398 3584 285404 3596
rect 284352 3556 285404 3584
rect 284352 3544 284358 3556
rect 285398 3544 285404 3556
rect 285456 3544 285462 3596
rect 289354 3544 289360 3596
rect 289412 3584 289418 3596
rect 505370 3584 505376 3596
rect 289412 3556 505376 3584
rect 289412 3544 289418 3556
rect 505370 3544 505376 3556
rect 505428 3544 505434 3596
rect 508498 3544 508504 3596
rect 508556 3584 508562 3596
rect 524230 3584 524236 3596
rect 508556 3556 524236 3584
rect 508556 3544 508562 3556
rect 524230 3544 524236 3556
rect 524288 3544 524294 3596
rect 534902 3544 534908 3596
rect 534960 3584 534966 3596
rect 536926 3584 536932 3596
rect 534960 3556 536932 3584
rect 534960 3544 534966 3556
rect 536926 3544 536932 3556
rect 536984 3544 536990 3596
rect 564434 3544 564440 3596
rect 564492 3584 564498 3596
rect 565630 3584 565636 3596
rect 564492 3556 565636 3584
rect 564492 3544 564498 3556
rect 565630 3544 565636 3556
rect 565688 3544 565694 3596
rect 574830 3544 574836 3596
rect 574888 3584 574894 3596
rect 577406 3584 577412 3596
rect 574888 3556 577412 3584
rect 574888 3544 574894 3556
rect 577406 3544 577412 3556
rect 577464 3544 577470 3596
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 10318 3516 10324 3528
rect 8812 3488 10324 3516
rect 8812 3476 8818 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24762 3516 24768 3528
rect 24268 3488 24768 3516
rect 24268 3476 24274 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 24872 3488 229784 3516
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 11698 3448 11704 3460
rect 4120 3420 11704 3448
rect 4120 3408 4126 3420
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 21818 3408 21824 3460
rect 21876 3448 21882 3460
rect 24872 3448 24900 3488
rect 21876 3420 24900 3448
rect 21876 3408 21882 3420
rect 32398 3408 32404 3460
rect 32456 3448 32462 3460
rect 33042 3448 33048 3460
rect 32456 3420 33048 3448
rect 32456 3408 32462 3420
rect 33042 3408 33048 3420
rect 33100 3408 33106 3460
rect 229756 3448 229784 3488
rect 229830 3476 229836 3528
rect 229888 3516 229894 3528
rect 230382 3516 230388 3528
rect 229888 3488 230388 3516
rect 229888 3476 229894 3488
rect 230382 3476 230388 3488
rect 230440 3476 230446 3528
rect 231026 3476 231032 3528
rect 231084 3516 231090 3528
rect 231762 3516 231768 3528
rect 231084 3488 231768 3516
rect 231084 3476 231090 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232222 3476 232228 3528
rect 232280 3516 232286 3528
rect 233142 3516 233148 3528
rect 232280 3488 233148 3516
rect 232280 3476 232286 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233418 3476 233424 3528
rect 233476 3516 233482 3528
rect 234522 3516 234528 3528
rect 233476 3488 234528 3516
rect 233476 3476 233482 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 237006 3476 237012 3528
rect 237064 3516 237070 3528
rect 249150 3516 249156 3528
rect 237064 3488 249156 3516
rect 237064 3476 237070 3488
rect 249150 3476 249156 3488
rect 249208 3476 249214 3528
rect 249978 3476 249984 3528
rect 250036 3516 250042 3528
rect 254578 3516 254584 3528
rect 250036 3488 254584 3516
rect 250036 3476 250042 3488
rect 254578 3476 254584 3488
rect 254636 3476 254642 3528
rect 254670 3476 254676 3528
rect 254728 3516 254734 3528
rect 255498 3516 255504 3528
rect 254728 3488 255504 3516
rect 254728 3476 254734 3488
rect 255498 3476 255504 3488
rect 255556 3476 255562 3528
rect 256510 3476 256516 3528
rect 256568 3516 256574 3528
rect 258258 3516 258264 3528
rect 256568 3488 258264 3516
rect 256568 3476 256574 3488
rect 258258 3476 258264 3488
rect 258316 3476 258322 3528
rect 258718 3476 258724 3528
rect 258776 3516 258782 3528
rect 259454 3516 259460 3528
rect 258776 3488 259460 3516
rect 258776 3476 258782 3488
rect 259454 3476 259460 3488
rect 259512 3476 259518 3528
rect 264698 3476 264704 3528
rect 264756 3516 264762 3528
rect 265342 3516 265348 3528
rect 264756 3488 265348 3516
rect 264756 3476 264762 3488
rect 265342 3476 265348 3488
rect 265400 3476 265406 3528
rect 289078 3476 289084 3528
rect 289136 3516 289142 3528
rect 508866 3516 508872 3528
rect 289136 3488 508872 3516
rect 289136 3476 289142 3488
rect 508866 3476 508872 3488
rect 508924 3476 508930 3528
rect 519630 3476 519636 3528
rect 519688 3516 519694 3528
rect 519688 3488 528554 3516
rect 519688 3476 519694 3488
rect 231302 3448 231308 3460
rect 33152 3420 229692 3448
rect 229756 3420 231308 3448
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 33152 3380 33180 3420
rect 40586 3380 40592 3392
rect 19484 3352 33180 3380
rect 35866 3352 40592 3380
rect 19484 3340 19490 3352
rect 26510 3272 26516 3324
rect 26568 3312 26574 3324
rect 35866 3312 35894 3352
rect 40586 3340 40592 3352
rect 40644 3340 40650 3392
rect 48958 3340 48964 3392
rect 49016 3380 49022 3392
rect 50338 3380 50344 3392
rect 49016 3352 50344 3380
rect 49016 3340 49022 3352
rect 50338 3340 50344 3352
rect 50396 3340 50402 3392
rect 52546 3340 52552 3392
rect 52604 3380 52610 3392
rect 53742 3380 53748 3392
rect 52604 3352 53748 3380
rect 52604 3340 52610 3352
rect 53742 3340 53748 3352
rect 53800 3340 53806 3392
rect 56042 3340 56048 3392
rect 56100 3380 56106 3392
rect 57146 3380 57152 3392
rect 56100 3352 57152 3380
rect 56100 3340 56106 3352
rect 57146 3340 57152 3352
rect 57204 3340 57210 3392
rect 57238 3340 57244 3392
rect 57296 3380 57302 3392
rect 57882 3380 57888 3392
rect 57296 3352 57888 3380
rect 57296 3340 57302 3352
rect 57882 3340 57888 3352
rect 57940 3340 57946 3392
rect 59630 3340 59636 3392
rect 59688 3380 59694 3392
rect 62758 3380 62764 3392
rect 59688 3352 62764 3380
rect 59688 3340 59694 3352
rect 62758 3340 62764 3352
rect 62816 3340 62822 3392
rect 64322 3340 64328 3392
rect 64380 3380 64386 3392
rect 64782 3380 64788 3392
rect 64380 3352 64788 3380
rect 64380 3340 64386 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 66714 3340 66720 3392
rect 66772 3380 66778 3392
rect 68278 3380 68284 3392
rect 66772 3352 68284 3380
rect 66772 3340 66778 3352
rect 68278 3340 68284 3352
rect 68336 3340 68342 3392
rect 72602 3340 72608 3392
rect 72660 3380 72666 3392
rect 73062 3380 73068 3392
rect 72660 3352 73068 3380
rect 72660 3340 72666 3352
rect 73062 3340 73068 3352
rect 73120 3340 73126 3392
rect 76190 3340 76196 3392
rect 76248 3380 76254 3392
rect 77202 3380 77208 3392
rect 76248 3352 77208 3380
rect 76248 3340 76254 3352
rect 77202 3340 77208 3352
rect 77260 3340 77266 3392
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 81342 3380 81348 3392
rect 80940 3352 81348 3380
rect 80940 3340 80946 3352
rect 81342 3340 81348 3352
rect 81400 3340 81406 3392
rect 83274 3340 83280 3392
rect 83332 3380 83338 3392
rect 84102 3380 84108 3392
rect 83332 3352 84108 3380
rect 83332 3340 83338 3352
rect 84102 3340 84108 3352
rect 84160 3340 84166 3392
rect 84470 3340 84476 3392
rect 84528 3380 84534 3392
rect 86218 3380 86224 3392
rect 84528 3352 86224 3380
rect 84528 3340 84534 3352
rect 86218 3340 86224 3352
rect 86276 3340 86282 3392
rect 89162 3340 89168 3392
rect 89220 3380 89226 3392
rect 89622 3380 89628 3392
rect 89220 3352 89628 3380
rect 89220 3340 89226 3352
rect 89622 3340 89628 3352
rect 89680 3340 89686 3392
rect 90358 3340 90364 3392
rect 90416 3380 90422 3392
rect 91002 3380 91008 3392
rect 90416 3352 91008 3380
rect 90416 3340 90422 3352
rect 91002 3340 91008 3352
rect 91060 3340 91066 3392
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 93118 3380 93124 3392
rect 91612 3352 93124 3380
rect 91612 3340 91618 3352
rect 93118 3340 93124 3352
rect 93176 3340 93182 3392
rect 93946 3340 93952 3392
rect 94004 3380 94010 3392
rect 95050 3380 95056 3392
rect 94004 3352 95056 3380
rect 94004 3340 94010 3352
rect 95050 3340 95056 3352
rect 95108 3340 95114 3392
rect 97442 3340 97448 3392
rect 97500 3380 97506 3392
rect 97902 3380 97908 3392
rect 97500 3352 97908 3380
rect 97500 3340 97506 3352
rect 97902 3340 97908 3352
rect 97960 3340 97966 3392
rect 98638 3340 98644 3392
rect 98696 3380 98702 3392
rect 99282 3380 99288 3392
rect 98696 3352 99288 3380
rect 98696 3340 98702 3352
rect 99282 3340 99288 3352
rect 99340 3340 99346 3392
rect 101030 3340 101036 3392
rect 101088 3380 101094 3392
rect 102042 3380 102048 3392
rect 101088 3352 102048 3380
rect 101088 3340 101094 3352
rect 102042 3340 102048 3352
rect 102100 3340 102106 3392
rect 102226 3340 102232 3392
rect 102284 3380 102290 3392
rect 229557 3383 229615 3389
rect 229557 3380 229569 3383
rect 102284 3352 229569 3380
rect 102284 3340 102290 3352
rect 229557 3349 229569 3352
rect 229603 3349 229615 3383
rect 229664 3380 229692 3420
rect 231302 3408 231308 3420
rect 231360 3408 231366 3460
rect 238110 3408 238116 3460
rect 238168 3448 238174 3460
rect 238168 3420 238754 3448
rect 238168 3408 238174 3420
rect 235258 3380 235264 3392
rect 229664 3352 235264 3380
rect 229557 3343 229615 3349
rect 235258 3340 235264 3352
rect 235316 3340 235322 3392
rect 238726 3380 238754 3420
rect 242894 3408 242900 3460
rect 242952 3448 242958 3460
rect 245102 3448 245108 3460
rect 242952 3420 245108 3448
rect 242952 3408 242958 3420
rect 245102 3408 245108 3420
rect 245160 3408 245166 3460
rect 248782 3408 248788 3460
rect 248840 3448 248846 3460
rect 253382 3448 253388 3460
rect 248840 3420 253388 3448
rect 248840 3408 248846 3420
rect 253382 3408 253388 3420
rect 253440 3408 253446 3460
rect 255866 3408 255872 3460
rect 255924 3448 255930 3460
rect 261754 3448 261760 3460
rect 255924 3420 261760 3448
rect 255924 3408 255930 3420
rect 261754 3408 261760 3420
rect 261812 3408 261818 3460
rect 289262 3408 289268 3460
rect 289320 3448 289326 3460
rect 512454 3448 512460 3460
rect 289320 3420 512460 3448
rect 289320 3408 289326 3420
rect 512454 3408 512460 3420
rect 512512 3408 512518 3460
rect 512638 3408 512644 3460
rect 512696 3448 512702 3460
rect 527818 3448 527824 3460
rect 512696 3420 527824 3448
rect 512696 3408 512702 3420
rect 527818 3408 527824 3420
rect 527876 3408 527882 3460
rect 528526 3448 528554 3488
rect 530578 3476 530584 3528
rect 530636 3516 530642 3528
rect 532510 3516 532516 3528
rect 530636 3488 532516 3516
rect 530636 3476 530642 3488
rect 532510 3476 532516 3488
rect 532568 3476 532574 3528
rect 536098 3476 536104 3528
rect 536156 3516 536162 3528
rect 537018 3516 537024 3528
rect 536156 3488 537024 3516
rect 536156 3476 536162 3488
rect 537018 3476 537024 3488
rect 537076 3476 537082 3528
rect 540330 3476 540336 3528
rect 540388 3516 540394 3528
rect 541986 3516 541992 3528
rect 540388 3488 541992 3516
rect 540388 3476 540394 3488
rect 541986 3476 541992 3488
rect 542044 3476 542050 3528
rect 548518 3476 548524 3528
rect 548576 3516 548582 3528
rect 552658 3516 552664 3528
rect 548576 3488 552664 3516
rect 548576 3476 548582 3488
rect 552658 3476 552664 3488
rect 552716 3476 552722 3528
rect 562318 3476 562324 3528
rect 562376 3516 562382 3528
rect 566826 3516 566832 3528
rect 562376 3488 566832 3516
rect 562376 3476 562382 3488
rect 566826 3476 566832 3488
rect 566884 3476 566890 3528
rect 531314 3448 531320 3460
rect 528526 3420 531320 3448
rect 531314 3408 531320 3420
rect 531372 3408 531378 3460
rect 538950 3408 538956 3460
rect 539008 3448 539014 3460
rect 539594 3448 539600 3460
rect 539008 3420 539600 3448
rect 539008 3408 539014 3420
rect 539594 3408 539600 3420
rect 539652 3408 539658 3460
rect 253290 3380 253296 3392
rect 238726 3352 253296 3380
rect 253290 3340 253296 3352
rect 253348 3340 253354 3392
rect 283558 3340 283564 3392
rect 283616 3380 283622 3392
rect 465721 3383 465779 3389
rect 465721 3380 465733 3383
rect 283616 3352 465733 3380
rect 283616 3340 283622 3352
rect 465721 3349 465733 3352
rect 465767 3349 465779 3383
rect 465721 3343 465779 3349
rect 468478 3340 468484 3392
rect 468536 3380 468542 3392
rect 469858 3380 469864 3392
rect 468536 3352 469864 3380
rect 468536 3340 468542 3352
rect 469858 3340 469864 3352
rect 469916 3340 469922 3392
rect 472618 3340 472624 3392
rect 472676 3380 472682 3392
rect 473446 3380 473452 3392
rect 472676 3352 473452 3380
rect 472676 3340 472682 3352
rect 473446 3340 473452 3352
rect 473504 3340 473510 3392
rect 476758 3340 476764 3392
rect 476816 3380 476822 3392
rect 478138 3380 478144 3392
rect 476816 3352 478144 3380
rect 476816 3340 476822 3352
rect 478138 3340 478144 3352
rect 478196 3340 478202 3392
rect 478233 3383 478291 3389
rect 478233 3349 478245 3383
rect 478279 3380 478291 3383
rect 480530 3380 480536 3392
rect 478279 3352 480536 3380
rect 478279 3349 478291 3352
rect 478233 3343 478291 3349
rect 480530 3340 480536 3352
rect 480588 3340 480594 3392
rect 26568 3284 35894 3312
rect 26568 3272 26574 3284
rect 41874 3272 41880 3324
rect 41932 3312 41938 3324
rect 106826 3312 106832 3324
rect 41932 3284 106832 3312
rect 41932 3272 41938 3284
rect 106826 3272 106832 3284
rect 106884 3272 106890 3324
rect 106918 3272 106924 3324
rect 106976 3312 106982 3324
rect 107562 3312 107568 3324
rect 106976 3284 107568 3312
rect 106976 3272 106982 3284
rect 107562 3272 107568 3284
rect 107620 3272 107626 3324
rect 108114 3272 108120 3324
rect 108172 3312 108178 3324
rect 108942 3312 108948 3324
rect 108172 3284 108948 3312
rect 108172 3272 108178 3284
rect 108942 3272 108948 3284
rect 109000 3272 109006 3324
rect 109310 3272 109316 3324
rect 109368 3312 109374 3324
rect 110322 3312 110328 3324
rect 109368 3284 110328 3312
rect 109368 3272 109374 3284
rect 110322 3272 110328 3284
rect 110380 3272 110386 3324
rect 115198 3272 115204 3324
rect 115256 3312 115262 3324
rect 115842 3312 115848 3324
rect 115256 3284 115848 3312
rect 115256 3272 115262 3284
rect 115842 3272 115848 3284
rect 115900 3272 115906 3324
rect 116394 3272 116400 3324
rect 116452 3312 116458 3324
rect 117222 3312 117228 3324
rect 116452 3284 117228 3312
rect 116452 3272 116458 3284
rect 117222 3272 117228 3284
rect 117280 3272 117286 3324
rect 118786 3272 118792 3324
rect 118844 3312 118850 3324
rect 119798 3312 119804 3324
rect 118844 3284 119804 3312
rect 118844 3272 118850 3284
rect 119798 3272 119804 3284
rect 119856 3272 119862 3324
rect 122282 3272 122288 3324
rect 122340 3312 122346 3324
rect 122742 3312 122748 3324
rect 122340 3284 122748 3312
rect 122340 3272 122346 3284
rect 122742 3272 122748 3284
rect 122800 3272 122806 3324
rect 123478 3272 123484 3324
rect 123536 3312 123542 3324
rect 124122 3312 124128 3324
rect 123536 3284 124128 3312
rect 123536 3272 123542 3284
rect 124122 3272 124128 3284
rect 124180 3272 124186 3324
rect 124674 3272 124680 3324
rect 124732 3312 124738 3324
rect 125502 3312 125508 3324
rect 124732 3284 125508 3312
rect 124732 3272 124738 3284
rect 125502 3272 125508 3284
rect 125560 3272 125566 3324
rect 126974 3272 126980 3324
rect 127032 3312 127038 3324
rect 128262 3312 128268 3324
rect 127032 3284 128268 3312
rect 127032 3272 127038 3284
rect 128262 3272 128268 3284
rect 128320 3272 128326 3324
rect 130562 3272 130568 3324
rect 130620 3312 130626 3324
rect 131022 3312 131028 3324
rect 130620 3284 131028 3312
rect 130620 3272 130626 3284
rect 131022 3272 131028 3284
rect 131080 3272 131086 3324
rect 131758 3272 131764 3324
rect 131816 3312 131822 3324
rect 132402 3312 132408 3324
rect 131816 3284 132408 3312
rect 131816 3272 131822 3284
rect 132402 3272 132408 3284
rect 132460 3272 132466 3324
rect 134150 3272 134156 3324
rect 134208 3312 134214 3324
rect 135162 3312 135168 3324
rect 134208 3284 135168 3312
rect 134208 3272 134214 3284
rect 135162 3272 135168 3284
rect 135220 3272 135226 3324
rect 138842 3272 138848 3324
rect 138900 3312 138906 3324
rect 139302 3312 139308 3324
rect 138900 3284 139308 3312
rect 138900 3272 138906 3284
rect 139302 3272 139308 3284
rect 139360 3272 139366 3324
rect 140038 3272 140044 3324
rect 140096 3312 140102 3324
rect 140682 3312 140688 3324
rect 140096 3284 140688 3312
rect 140096 3272 140102 3284
rect 140682 3272 140688 3284
rect 140740 3272 140746 3324
rect 244642 3312 244648 3324
rect 140792 3284 244648 3312
rect 35986 3204 35992 3256
rect 36044 3244 36050 3256
rect 47578 3244 47584 3256
rect 36044 3216 47584 3244
rect 36044 3204 36050 3216
rect 47578 3204 47584 3216
rect 47636 3204 47642 3256
rect 82078 3204 82084 3256
rect 82136 3244 82142 3256
rect 83458 3244 83464 3256
rect 82136 3216 83464 3244
rect 82136 3204 82142 3216
rect 83458 3204 83464 3216
rect 83516 3204 83522 3256
rect 105722 3204 105728 3256
rect 105780 3244 105786 3256
rect 106182 3244 106188 3256
rect 105780 3216 106188 3244
rect 105780 3204 105786 3216
rect 106182 3204 106188 3216
rect 106240 3204 106246 3256
rect 125870 3204 125876 3256
rect 125928 3244 125934 3256
rect 140792 3244 140820 3284
rect 244642 3272 244648 3284
rect 244700 3272 244706 3324
rect 251174 3272 251180 3324
rect 251232 3312 251238 3324
rect 255682 3312 255688 3324
rect 251232 3284 255688 3312
rect 251232 3272 251238 3284
rect 255682 3272 255688 3284
rect 255740 3272 255746 3324
rect 258350 3272 258356 3324
rect 258408 3312 258414 3324
rect 262950 3312 262956 3324
rect 258408 3284 262956 3312
rect 258408 3272 258414 3284
rect 262950 3272 262956 3284
rect 263008 3272 263014 3324
rect 282178 3272 282184 3324
rect 282236 3312 282242 3324
rect 292574 3312 292580 3324
rect 282236 3284 292580 3312
rect 282236 3272 282242 3284
rect 292574 3272 292580 3284
rect 292632 3272 292638 3324
rect 294598 3272 294604 3324
rect 294656 3312 294662 3324
rect 294656 3284 475332 3312
rect 294656 3272 294662 3284
rect 244918 3244 244924 3256
rect 125928 3216 140820 3244
rect 140884 3216 244924 3244
rect 125928 3204 125934 3216
rect 18230 3136 18236 3188
rect 18288 3176 18294 3188
rect 25498 3176 25504 3188
rect 18288 3148 25504 3176
rect 18288 3136 18294 3148
rect 25498 3136 25504 3148
rect 25556 3136 25562 3188
rect 65518 3136 65524 3188
rect 65576 3176 65582 3188
rect 66162 3176 66168 3188
rect 65576 3148 66168 3176
rect 65576 3136 65582 3148
rect 66162 3136 66168 3148
rect 66220 3136 66226 3188
rect 114002 3136 114008 3188
rect 114060 3176 114066 3188
rect 115106 3176 115112 3188
rect 114060 3148 115112 3176
rect 114060 3136 114066 3148
rect 115106 3136 115112 3148
rect 115164 3136 115170 3188
rect 132954 3136 132960 3188
rect 133012 3176 133018 3188
rect 140884 3176 140912 3216
rect 244918 3204 244924 3216
rect 244976 3204 244982 3256
rect 264422 3204 264428 3256
rect 264480 3244 264486 3256
rect 270034 3244 270040 3256
rect 264480 3216 270040 3244
rect 264480 3204 264486 3216
rect 270034 3204 270040 3216
rect 270092 3204 270098 3256
rect 281074 3204 281080 3256
rect 281132 3244 281138 3256
rect 461578 3244 461584 3256
rect 281132 3216 461584 3244
rect 281132 3204 281138 3216
rect 461578 3204 461584 3216
rect 461636 3204 461642 3256
rect 465721 3247 465779 3253
rect 465721 3213 465733 3247
rect 465767 3244 465779 3247
rect 472250 3244 472256 3256
rect 465767 3216 472256 3244
rect 465767 3213 465779 3216
rect 465721 3207 465779 3213
rect 472250 3204 472256 3216
rect 472308 3204 472314 3256
rect 475304 3244 475332 3284
rect 475378 3272 475384 3324
rect 475436 3312 475442 3324
rect 476942 3312 476948 3324
rect 475436 3284 476948 3312
rect 475436 3272 475442 3284
rect 476942 3272 476948 3284
rect 477000 3272 477006 3324
rect 479518 3272 479524 3324
rect 479576 3312 479582 3324
rect 482830 3312 482836 3324
rect 479576 3284 482836 3312
rect 479576 3272 479582 3284
rect 482830 3272 482836 3284
rect 482888 3272 482894 3324
rect 493318 3272 493324 3324
rect 493376 3312 493382 3324
rect 499390 3312 499396 3324
rect 493376 3284 499396 3312
rect 493376 3272 493382 3284
rect 499390 3272 499396 3284
rect 499448 3272 499454 3324
rect 569218 3272 569224 3324
rect 569276 3312 569282 3324
rect 570322 3312 570328 3324
rect 569276 3284 570328 3312
rect 569276 3272 569282 3284
rect 570322 3272 570328 3284
rect 570380 3272 570386 3324
rect 479334 3244 479340 3256
rect 475304 3216 479340 3244
rect 479334 3204 479340 3216
rect 479392 3204 479398 3256
rect 133012 3148 140912 3176
rect 133012 3136 133018 3148
rect 141234 3136 141240 3188
rect 141292 3176 141298 3188
rect 142062 3176 142068 3188
rect 141292 3148 142068 3176
rect 141292 3136 141298 3148
rect 142062 3136 142068 3148
rect 142120 3136 142126 3188
rect 142430 3136 142436 3188
rect 142488 3176 142494 3188
rect 143442 3176 143448 3188
rect 142488 3148 143448 3176
rect 142488 3136 142494 3148
rect 143442 3136 143448 3148
rect 143500 3136 143506 3188
rect 147122 3136 147128 3188
rect 147180 3176 147186 3188
rect 147582 3176 147588 3188
rect 147180 3148 147588 3176
rect 147180 3136 147186 3148
rect 147582 3136 147588 3148
rect 147640 3136 147646 3188
rect 148318 3136 148324 3188
rect 148376 3176 148382 3188
rect 148962 3176 148968 3188
rect 148376 3148 148968 3176
rect 148376 3136 148382 3148
rect 148962 3136 148968 3148
rect 149020 3136 149026 3188
rect 149514 3136 149520 3188
rect 149572 3176 149578 3188
rect 150342 3176 150348 3188
rect 149572 3148 150348 3176
rect 149572 3136 149578 3148
rect 150342 3136 150348 3148
rect 150400 3136 150406 3188
rect 246114 3176 246120 3188
rect 150452 3148 246120 3176
rect 40678 3068 40684 3120
rect 40736 3108 40742 3120
rect 44818 3108 44824 3120
rect 40736 3080 44824 3108
rect 40736 3068 40742 3080
rect 44818 3068 44824 3080
rect 44876 3068 44882 3120
rect 143534 3068 143540 3120
rect 143592 3108 143598 3120
rect 150452 3108 150480 3148
rect 246114 3136 246120 3148
rect 246172 3136 246178 3188
rect 279786 3136 279792 3188
rect 279844 3176 279850 3188
rect 458082 3176 458088 3188
rect 279844 3148 458088 3176
rect 279844 3136 279850 3148
rect 458082 3136 458088 3148
rect 458140 3136 458146 3188
rect 538858 3136 538864 3188
rect 538916 3176 538922 3188
rect 540790 3176 540796 3188
rect 538916 3148 540796 3176
rect 538916 3136 538922 3148
rect 540790 3136 540796 3148
rect 540848 3136 540854 3188
rect 542998 3136 543004 3188
rect 543056 3176 543062 3188
rect 545482 3176 545488 3188
rect 543056 3148 545488 3176
rect 543056 3136 543062 3148
rect 545482 3136 545488 3148
rect 545540 3136 545546 3188
rect 143592 3080 150480 3108
rect 143592 3068 143598 3080
rect 150618 3068 150624 3120
rect 150676 3108 150682 3120
rect 151722 3108 151728 3120
rect 150676 3080 151728 3108
rect 150676 3068 150682 3080
rect 151722 3068 151728 3080
rect 151780 3068 151786 3120
rect 151814 3068 151820 3120
rect 151872 3108 151878 3120
rect 153102 3108 153108 3120
rect 151872 3080 153108 3108
rect 151872 3068 151878 3080
rect 153102 3068 153108 3080
rect 153160 3068 153166 3120
rect 155402 3068 155408 3120
rect 155460 3108 155466 3120
rect 155862 3108 155868 3120
rect 155460 3080 155868 3108
rect 155460 3068 155466 3080
rect 155862 3068 155868 3080
rect 155920 3068 155926 3120
rect 156598 3068 156604 3120
rect 156656 3108 156662 3120
rect 157242 3108 157248 3120
rect 156656 3080 157248 3108
rect 156656 3068 156662 3080
rect 157242 3068 157248 3080
rect 157300 3068 157306 3120
rect 157794 3068 157800 3120
rect 157852 3108 157858 3120
rect 158622 3108 158628 3120
rect 157852 3080 158628 3108
rect 157852 3068 157858 3080
rect 158622 3068 158628 3080
rect 158680 3068 158686 3120
rect 158898 3068 158904 3120
rect 158956 3108 158962 3120
rect 160002 3108 160008 3120
rect 158956 3080 160008 3108
rect 158956 3068 158962 3080
rect 160002 3068 160008 3080
rect 160060 3068 160066 3120
rect 160094 3068 160100 3120
rect 160152 3108 160158 3120
rect 161382 3108 161388 3120
rect 160152 3080 161388 3108
rect 160152 3068 160158 3080
rect 161382 3068 161388 3080
rect 161440 3068 161446 3120
rect 163682 3068 163688 3120
rect 163740 3108 163746 3120
rect 164142 3108 164148 3120
rect 163740 3080 164148 3108
rect 163740 3068 163746 3080
rect 164142 3068 164148 3080
rect 164200 3068 164206 3120
rect 164878 3068 164884 3120
rect 164936 3108 164942 3120
rect 165522 3108 165528 3120
rect 164936 3080 165528 3108
rect 164936 3068 164942 3080
rect 165522 3068 165528 3080
rect 165580 3068 165586 3120
rect 166074 3068 166080 3120
rect 166132 3108 166138 3120
rect 166902 3108 166908 3120
rect 166132 3080 166908 3108
rect 166132 3068 166138 3080
rect 166902 3068 166908 3080
rect 166960 3068 166966 3120
rect 167178 3068 167184 3120
rect 167236 3108 167242 3120
rect 168282 3108 168288 3120
rect 167236 3080 168288 3108
rect 167236 3068 167242 3080
rect 168282 3068 168288 3080
rect 168340 3068 168346 3120
rect 168374 3068 168380 3120
rect 168432 3108 168438 3120
rect 169662 3108 169668 3120
rect 168432 3080 169668 3108
rect 168432 3068 168438 3080
rect 169662 3068 169668 3080
rect 169720 3068 169726 3120
rect 169757 3111 169815 3117
rect 169757 3077 169769 3111
rect 169803 3108 169815 3111
rect 232498 3108 232504 3120
rect 169803 3080 232504 3108
rect 169803 3077 169815 3080
rect 169757 3071 169815 3077
rect 232498 3068 232504 3080
rect 232556 3068 232562 3120
rect 278038 3068 278044 3120
rect 278096 3108 278102 3120
rect 445018 3108 445024 3120
rect 278096 3080 445024 3108
rect 278096 3068 278102 3080
rect 445018 3068 445024 3080
rect 445076 3068 445082 3120
rect 472710 3068 472716 3120
rect 472768 3108 472774 3120
rect 474550 3108 474556 3120
rect 472768 3080 474556 3108
rect 472768 3068 472774 3080
rect 474550 3068 474556 3080
rect 474608 3068 474614 3120
rect 12342 3000 12348 3052
rect 12400 3040 12406 3052
rect 14458 3040 14464 3052
rect 12400 3012 14464 3040
rect 12400 3000 12406 3012
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 58434 3000 58440 3052
rect 58492 3040 58498 3052
rect 61378 3040 61384 3052
rect 58492 3012 61384 3040
rect 58492 3000 58498 3012
rect 61378 3000 61384 3012
rect 61436 3000 61442 3052
rect 117590 3000 117596 3052
rect 117648 3040 117654 3052
rect 173069 3043 173127 3049
rect 117648 3012 169892 3040
rect 117648 3000 117654 3012
rect 37182 2932 37188 2984
rect 37240 2972 37246 2984
rect 43530 2972 43536 2984
rect 37240 2944 43536 2972
rect 37240 2932 37246 2944
rect 43530 2932 43536 2944
rect 43588 2932 43594 2984
rect 73798 2932 73804 2984
rect 73856 2972 73862 2984
rect 75178 2972 75184 2984
rect 73856 2944 75184 2972
rect 73856 2932 73862 2944
rect 75178 2932 75184 2944
rect 75236 2932 75242 2984
rect 77386 2932 77392 2984
rect 77444 2972 77450 2984
rect 80698 2972 80704 2984
rect 77444 2944 80704 2972
rect 77444 2932 77450 2944
rect 80698 2932 80704 2944
rect 80756 2932 80762 2984
rect 110506 2932 110512 2984
rect 110564 2972 110570 2984
rect 110564 2944 161474 2972
rect 110564 2932 110570 2944
rect 161446 2904 161474 2944
rect 161566 2932 161572 2984
rect 161624 2972 161630 2984
rect 169573 2975 169631 2981
rect 169573 2972 169585 2975
rect 161624 2944 169585 2972
rect 161624 2932 161630 2944
rect 169573 2941 169585 2944
rect 169619 2941 169631 2975
rect 169864 2972 169892 3012
rect 173069 3009 173081 3043
rect 173115 3040 173127 3043
rect 180150 3040 180156 3052
rect 173115 3012 180156 3040
rect 173115 3009 173127 3012
rect 173069 3003 173127 3009
rect 180150 3000 180156 3012
rect 180208 3000 180214 3052
rect 197906 3000 197912 3052
rect 197964 3040 197970 3052
rect 208397 3043 208455 3049
rect 208397 3040 208409 3043
rect 197964 3012 208409 3040
rect 197964 3000 197970 3012
rect 208397 3009 208409 3012
rect 208443 3009 208455 3043
rect 208397 3003 208455 3009
rect 208578 3000 208584 3052
rect 208636 3040 208642 3052
rect 251542 3040 251548 3052
rect 208636 3012 251548 3040
rect 208636 3000 208642 3012
rect 251542 3000 251548 3012
rect 251600 3000 251606 3052
rect 282270 3000 282276 3052
rect 282328 3040 282334 3052
rect 427262 3040 427268 3052
rect 282328 3012 427268 3040
rect 282328 3000 282334 3012
rect 427262 3000 427268 3012
rect 427320 3000 427326 3052
rect 429838 3000 429844 3052
rect 429896 3040 429902 3052
rect 434438 3040 434444 3052
rect 429896 3012 434444 3040
rect 429896 3000 429902 3012
rect 434438 3000 434444 3012
rect 434496 3000 434502 3052
rect 439590 3000 439596 3052
rect 439648 3040 439654 3052
rect 441522 3040 441528 3052
rect 439648 3012 441528 3040
rect 439648 3000 439654 3012
rect 441522 3000 441528 3012
rect 441580 3000 441586 3052
rect 459186 3040 459192 3052
rect 441816 3012 459192 3040
rect 178678 2972 178684 2984
rect 169864 2944 178684 2972
rect 169573 2935 169631 2941
rect 178678 2932 178684 2944
rect 178736 2932 178742 2984
rect 212813 2975 212871 2981
rect 212813 2941 212825 2975
rect 212859 2972 212871 2975
rect 215938 2972 215944 2984
rect 212859 2944 215944 2972
rect 212859 2941 212871 2944
rect 212813 2935 212871 2941
rect 215938 2932 215944 2944
rect 215996 2932 216002 2984
rect 229557 2975 229615 2981
rect 229557 2941 229569 2975
rect 229603 2972 229615 2975
rect 236638 2972 236644 2984
rect 229603 2944 236644 2972
rect 229603 2941 229615 2944
rect 229557 2935 229615 2941
rect 236638 2932 236644 2944
rect 236696 2932 236702 2984
rect 266998 2932 267004 2984
rect 267056 2972 267062 2984
rect 337470 2972 337476 2984
rect 267056 2944 337476 2972
rect 267056 2932 267062 2944
rect 337470 2932 337476 2944
rect 337528 2932 337534 2984
rect 337562 2932 337568 2984
rect 337620 2972 337626 2984
rect 337620 2944 341104 2972
rect 337620 2932 337626 2944
rect 171778 2904 171784 2916
rect 161446 2876 171784 2904
rect 171778 2864 171784 2876
rect 171836 2864 171842 2916
rect 171962 2864 171968 2916
rect 172020 2904 172026 2916
rect 231394 2904 231400 2916
rect 172020 2876 231400 2904
rect 172020 2864 172026 2876
rect 231394 2864 231400 2876
rect 231452 2864 231458 2916
rect 258902 2864 258908 2916
rect 258960 2904 258966 2916
rect 296070 2904 296076 2916
rect 258960 2876 296076 2904
rect 258960 2864 258966 2876
rect 296070 2864 296076 2876
rect 296128 2864 296134 2916
rect 300210 2864 300216 2916
rect 300268 2904 300274 2916
rect 340966 2904 340972 2916
rect 300268 2876 340972 2904
rect 300268 2864 300274 2876
rect 340966 2864 340972 2876
rect 341024 2864 341030 2916
rect 341076 2904 341104 2944
rect 341518 2932 341524 2984
rect 341576 2972 341582 2984
rect 344833 2975 344891 2981
rect 341576 2944 344784 2972
rect 341576 2932 341582 2944
rect 344189 2907 344247 2913
rect 344189 2904 344201 2907
rect 341076 2876 344201 2904
rect 344189 2873 344201 2876
rect 344235 2873 344247 2907
rect 344189 2867 344247 2873
rect 344278 2864 344284 2916
rect 344336 2904 344342 2916
rect 344756 2904 344784 2944
rect 344833 2941 344845 2975
rect 344879 2972 344891 2975
rect 348050 2972 348056 2984
rect 344879 2944 348056 2972
rect 344879 2941 344891 2944
rect 344833 2935 344891 2941
rect 348050 2932 348056 2944
rect 348108 2932 348114 2984
rect 348418 2932 348424 2984
rect 348476 2972 348482 2984
rect 365625 2975 365683 2981
rect 365625 2972 365637 2975
rect 348476 2944 365637 2972
rect 348476 2932 348482 2944
rect 365625 2941 365637 2944
rect 365671 2941 365683 2975
rect 365625 2935 365683 2941
rect 365714 2932 365720 2984
rect 365772 2972 365778 2984
rect 367002 2972 367008 2984
rect 365772 2944 367008 2972
rect 365772 2932 365778 2944
rect 367002 2932 367008 2944
rect 367060 2932 367066 2984
rect 367097 2975 367155 2981
rect 367097 2941 367109 2975
rect 367143 2972 367155 2975
rect 369394 2972 369400 2984
rect 367143 2944 369400 2972
rect 367143 2941 367155 2944
rect 367097 2935 367155 2941
rect 369394 2932 369400 2944
rect 369452 2932 369458 2984
rect 369486 2932 369492 2984
rect 369544 2972 369550 2984
rect 390646 2972 390652 2984
rect 369544 2944 390652 2972
rect 369544 2932 369550 2944
rect 390646 2932 390652 2944
rect 390704 2932 390710 2984
rect 391198 2932 391204 2984
rect 391256 2972 391262 2984
rect 398377 2975 398435 2981
rect 391256 2944 398144 2972
rect 391256 2932 391262 2944
rect 355226 2904 355232 2916
rect 344336 2876 344692 2904
rect 344756 2876 355232 2904
rect 344336 2864 344342 2876
rect 121086 2796 121092 2848
rect 121144 2836 121150 2848
rect 180058 2836 180064 2848
rect 121144 2808 180064 2836
rect 121144 2796 121150 2808
rect 180058 2796 180064 2808
rect 180116 2796 180122 2848
rect 269758 2796 269764 2848
rect 269816 2836 269822 2848
rect 305546 2836 305552 2848
rect 269816 2808 305552 2836
rect 269816 2796 269822 2808
rect 305546 2796 305552 2808
rect 305604 2796 305610 2848
rect 316034 2796 316040 2848
rect 316092 2836 316098 2848
rect 317322 2836 317328 2848
rect 316092 2808 317328 2836
rect 316092 2796 316098 2808
rect 317322 2796 317328 2808
rect 317380 2796 317386 2848
rect 344554 2836 344560 2848
rect 317432 2808 344560 2836
rect 316678 2728 316684 2780
rect 316736 2768 316742 2780
rect 317432 2768 317460 2808
rect 344554 2796 344560 2808
rect 344612 2796 344618 2848
rect 344664 2836 344692 2876
rect 355226 2864 355232 2876
rect 355284 2864 355290 2916
rect 355318 2864 355324 2916
rect 355376 2904 355382 2916
rect 376478 2904 376484 2916
rect 355376 2876 376484 2904
rect 355376 2864 355382 2876
rect 376478 2864 376484 2876
rect 376536 2864 376542 2916
rect 376570 2864 376576 2916
rect 376628 2904 376634 2916
rect 397730 2904 397736 2916
rect 376628 2876 397736 2904
rect 376628 2864 376634 2876
rect 397730 2864 397736 2876
rect 397788 2864 397794 2916
rect 398116 2904 398144 2944
rect 398377 2941 398389 2975
rect 398423 2972 398435 2975
rect 404814 2972 404820 2984
rect 398423 2944 404820 2972
rect 398423 2941 398435 2944
rect 398377 2935 398435 2941
rect 404814 2932 404820 2944
rect 404872 2932 404878 2984
rect 404998 2932 405004 2984
rect 405056 2972 405062 2984
rect 405458 2972 405464 2984
rect 405056 2944 405464 2972
rect 405056 2932 405062 2944
rect 405458 2932 405464 2944
rect 405516 2932 405522 2984
rect 405553 2975 405611 2981
rect 405553 2941 405565 2975
rect 405599 2972 405611 2975
rect 415486 2972 415492 2984
rect 405599 2944 415492 2972
rect 405599 2941 405611 2944
rect 405553 2935 405611 2941
rect 415486 2932 415492 2944
rect 415544 2932 415550 2984
rect 416038 2932 416044 2984
rect 416096 2972 416102 2984
rect 418709 2975 418767 2981
rect 418709 2972 418721 2975
rect 416096 2944 418721 2972
rect 416096 2932 416102 2944
rect 418709 2941 418721 2944
rect 418755 2941 418767 2975
rect 418709 2935 418767 2941
rect 418798 2932 418804 2984
rect 418856 2972 418862 2984
rect 420178 2972 420184 2984
rect 418856 2944 420184 2972
rect 418856 2932 418862 2944
rect 420178 2932 420184 2944
rect 420236 2932 420242 2984
rect 420273 2975 420331 2981
rect 420273 2941 420285 2975
rect 420319 2972 420331 2975
rect 426158 2972 426164 2984
rect 420319 2944 426164 2972
rect 420319 2941 420331 2944
rect 420273 2935 420331 2941
rect 426158 2932 426164 2944
rect 426216 2932 426222 2984
rect 432598 2932 432604 2984
rect 432656 2972 432662 2984
rect 437934 2972 437940 2984
rect 432656 2944 437940 2972
rect 432656 2932 432662 2944
rect 437934 2932 437940 2944
rect 437992 2932 437998 2984
rect 438210 2932 438216 2984
rect 438268 2972 438274 2984
rect 441816 2972 441844 3012
rect 459186 3000 459192 3012
rect 459244 3000 459250 3052
rect 438268 2944 441844 2972
rect 438268 2932 438274 2944
rect 408402 2904 408408 2916
rect 398116 2876 408408 2904
rect 408402 2864 408408 2876
rect 408460 2864 408466 2916
rect 422570 2904 422576 2916
rect 409340 2876 422576 2904
rect 362310 2836 362316 2848
rect 344664 2808 362316 2836
rect 362310 2796 362316 2808
rect 362368 2796 362374 2848
rect 362402 2796 362408 2848
rect 362460 2836 362466 2848
rect 398193 2839 398251 2845
rect 398193 2836 398205 2839
rect 362460 2808 382780 2836
rect 362460 2796 362466 2808
rect 316736 2740 317460 2768
rect 365625 2771 365683 2777
rect 316736 2728 316742 2740
rect 365625 2737 365637 2771
rect 365671 2768 365683 2771
rect 367097 2771 367155 2777
rect 367097 2768 367109 2771
rect 365671 2740 367109 2768
rect 365671 2737 365683 2740
rect 365625 2731 365683 2737
rect 367097 2737 367109 2740
rect 367143 2737 367155 2771
rect 367097 2731 367155 2737
rect 382752 2632 382780 2808
rect 383672 2808 398205 2836
rect 383672 2768 383700 2808
rect 398193 2805 398205 2808
rect 398239 2805 398251 2839
rect 398193 2799 398251 2805
rect 398282 2796 398288 2848
rect 398340 2836 398346 2848
rect 405553 2839 405611 2845
rect 405553 2836 405565 2839
rect 398340 2808 405565 2836
rect 398340 2796 398346 2808
rect 405553 2805 405565 2808
rect 405599 2805 405611 2839
rect 405553 2799 405611 2805
rect 405642 2796 405648 2848
rect 405700 2836 405706 2848
rect 405700 2808 407712 2836
rect 405700 2796 405706 2808
rect 383626 2740 383700 2768
rect 407684 2768 407712 2808
rect 407758 2796 407764 2848
rect 407816 2836 407822 2848
rect 409340 2836 409368 2876
rect 422570 2864 422576 2876
rect 422628 2864 422634 2916
rect 422938 2864 422944 2916
rect 422996 2904 423002 2916
rect 436738 2904 436744 2916
rect 422996 2876 436744 2904
rect 422996 2864 423002 2876
rect 436738 2864 436744 2876
rect 436796 2864 436802 2916
rect 439498 2864 439504 2916
rect 439556 2904 439562 2916
rect 448606 2904 448612 2916
rect 439556 2876 448612 2904
rect 439556 2864 439562 2876
rect 448606 2864 448612 2876
rect 448664 2864 448670 2916
rect 490558 2864 490564 2916
rect 490616 2904 490622 2916
rect 495894 2904 495900 2916
rect 490616 2876 495900 2904
rect 490616 2864 490622 2876
rect 495894 2864 495900 2876
rect 495952 2864 495958 2916
rect 558270 2864 558276 2916
rect 558328 2904 558334 2916
rect 563238 2904 563244 2916
rect 558328 2876 563244 2904
rect 558328 2864 558334 2876
rect 563238 2864 563244 2876
rect 563296 2864 563302 2916
rect 418982 2836 418988 2848
rect 407816 2808 409368 2836
rect 409432 2808 418988 2836
rect 407816 2796 407822 2808
rect 409432 2768 409460 2808
rect 418982 2796 418988 2808
rect 419040 2796 419046 2848
rect 420181 2839 420239 2845
rect 420181 2836 420193 2839
rect 419092 2808 420193 2836
rect 407684 2740 409460 2768
rect 418709 2771 418767 2777
rect 382918 2660 382924 2712
rect 382976 2700 382982 2712
rect 383626 2700 383654 2740
rect 418709 2737 418721 2771
rect 418755 2768 418767 2771
rect 419092 2768 419120 2808
rect 420181 2805 420193 2808
rect 420227 2805 420239 2839
rect 420181 2799 420239 2805
rect 420270 2796 420276 2848
rect 420328 2836 420334 2848
rect 433242 2836 433248 2848
rect 420328 2808 433248 2836
rect 420328 2796 420334 2808
rect 433242 2796 433248 2808
rect 433300 2796 433306 2848
rect 438118 2796 438124 2848
rect 438176 2836 438182 2848
rect 452102 2836 452108 2848
rect 438176 2808 452108 2836
rect 438176 2796 438182 2808
rect 452102 2796 452108 2808
rect 452160 2796 452166 2848
rect 583386 2836 583392 2848
rect 583347 2808 583392 2836
rect 583386 2796 583392 2808
rect 583444 2796 583450 2848
rect 418755 2740 419120 2768
rect 418755 2737 418767 2740
rect 418709 2731 418767 2737
rect 382976 2672 383654 2700
rect 382976 2660 382982 2672
rect 383562 2632 383568 2644
rect 382752 2604 383568 2632
rect 383562 2592 383568 2604
rect 383620 2592 383626 2644
rect 349154 1504 349160 1556
rect 349212 1544 349218 1556
rect 350442 1544 350448 1556
rect 349212 1516 350448 1544
rect 349212 1504 349218 1516
rect 350442 1504 350448 1516
rect 350500 1504 350506 1556
<< via1 >>
rect 254952 700952 255004 701004
rect 397460 700952 397512 701004
rect 255044 700884 255096 700936
rect 413652 700884 413704 700936
rect 89168 700816 89220 700868
rect 259644 700816 259696 700868
rect 273904 700816 273956 700868
rect 300124 700816 300176 700868
rect 72976 700748 73028 700800
rect 259736 700748 259788 700800
rect 271144 700748 271196 700800
rect 364984 700748 365036 700800
rect 253664 700680 253716 700732
rect 462320 700680 462372 700732
rect 40500 700612 40552 700664
rect 260840 700612 260892 700664
rect 269764 700612 269816 700664
rect 429844 700612 429896 700664
rect 255136 700544 255188 700596
rect 478512 700544 478564 700596
rect 24308 700476 24360 700528
rect 261024 700476 261076 700528
rect 282184 700476 282236 700528
rect 494796 700476 494848 700528
rect 170312 700408 170364 700460
rect 240784 700408 240836 700460
rect 252192 700408 252244 700460
rect 527180 700408 527232 700460
rect 8116 700340 8168 700392
rect 260932 700340 260984 700392
rect 280804 700340 280856 700392
rect 559656 700340 559708 700392
rect 105452 700272 105504 700324
rect 242164 700272 242216 700324
rect 253756 700272 253808 700324
rect 543464 700272 543516 700324
rect 137836 700204 137888 700256
rect 258172 700204 258224 700256
rect 154120 700136 154172 700188
rect 259552 700136 259604 700188
rect 256424 700068 256476 700120
rect 348792 700068 348844 700120
rect 256516 700000 256568 700052
rect 332508 700000 332560 700052
rect 202788 699932 202840 699984
rect 258264 699932 258316 699984
rect 218980 699864 219032 699916
rect 258356 699864 258408 699916
rect 257896 699796 257948 699848
rect 283840 699796 283892 699848
rect 257988 699728 258040 699780
rect 267648 699728 267700 699780
rect 235172 699660 235224 699712
rect 238024 699660 238076 699712
rect 252376 696940 252428 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 261116 683204 261168 683256
rect 252284 683136 252336 683188
rect 580172 683136 580224 683188
rect 3424 670760 3476 670812
rect 262220 670760 262272 670812
rect 251088 670692 251140 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 262312 656888 262364 656940
rect 250996 643084 251048 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 262404 632068 262456 632120
rect 250904 630640 250956 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 263600 618264 263652 618316
rect 250812 616836 250864 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 263692 605820 263744 605872
rect 249708 590656 249760 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 263784 579640 263836 579692
rect 249616 576852 249668 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 264980 565836 265032 565888
rect 249524 563048 249576 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 263876 553392 263928 553444
rect 248328 536800 248380 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 265072 527144 265124 527196
rect 248236 524424 248288 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 265164 514768 265216 514820
rect 248144 510620 248196 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 265256 500964 265308 501016
rect 246948 484372 247000 484424
rect 580172 484372 580224 484424
rect 3424 474716 3476 474768
rect 266360 474716 266412 474768
rect 248052 470568 248104 470620
rect 579988 470568 580040 470620
rect 3240 462340 3292 462392
rect 266452 462340 266504 462392
rect 246856 456764 246908 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 266544 448536 266596 448588
rect 246764 430584 246816 430636
rect 580172 430584 580224 430636
rect 3424 422288 3476 422340
rect 267740 422288 267792 422340
rect 246672 418140 246724 418192
rect 580172 418140 580224 418192
rect 3148 409844 3200 409896
rect 267832 409844 267884 409896
rect 245568 404336 245620 404388
rect 580172 404336 580224 404388
rect 3424 397468 3476 397520
rect 268016 397468 268068 397520
rect 242164 391756 242216 391808
rect 259736 391756 259788 391808
rect 269764 391756 269816 391808
rect 255688 391688 255740 391740
rect 271144 391688 271196 391740
rect 256608 391552 256660 391604
rect 273904 391552 273956 391604
rect 254584 391484 254636 391536
rect 240784 391416 240836 391468
rect 258632 391416 258684 391468
rect 238024 391348 238076 391400
rect 257620 391348 257672 391400
rect 252008 391280 252060 391332
rect 280804 391280 280856 391332
rect 253480 391212 253532 391264
rect 282184 391212 282236 391264
rect 242808 390464 242860 390516
rect 245936 390396 245988 390448
rect 246764 390396 246816 390448
rect 247408 390396 247460 390448
rect 248052 390396 248104 390448
rect 248972 390396 249024 390448
rect 249524 390396 249576 390448
rect 250076 390396 250128 390448
rect 250720 390396 250772 390448
rect 251916 390396 251968 390448
rect 252284 390396 252336 390448
rect 253020 390396 253072 390448
rect 253756 390396 253808 390448
rect 244004 390328 244056 390380
rect 249340 390328 249392 390380
rect 249708 390328 249760 390380
rect 250444 390328 250496 390380
rect 250996 390328 251048 390380
rect 251548 390328 251600 390380
rect 252376 390328 252428 390380
rect 257160 390464 257212 390516
rect 257988 390464 258040 390516
rect 258172 390464 258224 390516
rect 259000 390464 259052 390516
rect 259644 390464 259696 390516
rect 260472 390464 260524 390516
rect 262220 390464 262272 390516
rect 262772 390464 262824 390516
rect 265164 390464 265216 390516
rect 266084 390464 266136 390516
rect 266452 390464 266504 390516
rect 267280 390464 267332 390516
rect 267832 390464 267884 390516
rect 268384 390464 268436 390516
rect 280896 390464 280948 390516
rect 291936 390464 291988 390516
rect 254216 390396 254268 390448
rect 255136 390396 255188 390448
rect 256056 390396 256108 390448
rect 256516 390396 256568 390448
rect 540428 390396 540480 390448
rect 544476 390328 544528 390380
rect 547236 390260 547288 390312
rect 245200 390192 245252 390244
rect 241796 390124 241848 390176
rect 241428 390056 241480 390108
rect 285128 390124 285180 390176
rect 286508 390124 286560 390176
rect 289084 390124 289136 390176
rect 152464 389988 152516 390040
rect 277492 389988 277544 390040
rect 285036 390056 285088 390108
rect 292212 390056 292264 390108
rect 282368 389988 282420 390040
rect 292028 389988 292080 390040
rect 248144 389920 248196 389972
rect 248328 389920 248380 389972
rect 395344 389920 395396 389972
rect 40776 389852 40828 389904
rect 273996 389852 274048 389904
rect 281356 389852 281408 389904
rect 291844 389852 291896 389904
rect 39396 389784 39448 389836
rect 272892 389784 272944 389836
rect 281264 389784 281316 389836
rect 296076 389784 296128 389836
rect 36636 389716 36688 389768
rect 271880 389716 271932 389768
rect 279700 389716 279752 389768
rect 288072 389716 288124 389768
rect 35256 389648 35308 389700
rect 270592 389648 270644 389700
rect 282736 389648 282788 389700
rect 292120 389648 292172 389700
rect 33784 389580 33836 389632
rect 275100 389580 275152 389632
rect 278688 389580 278740 389632
rect 294696 389580 294748 389632
rect 35164 389512 35216 389564
rect 276296 389512 276348 389564
rect 280068 389512 280120 389564
rect 418896 389512 418948 389564
rect 15844 389444 15896 389496
rect 269488 389444 269540 389496
rect 284576 389444 284628 389496
rect 439688 389444 439740 389496
rect 21364 389376 21416 389428
rect 277032 389376 277084 389428
rect 282828 389376 282880 389428
rect 438308 389376 438360 389428
rect 242532 389308 242584 389360
rect 279332 389308 279384 389360
rect 288164 389308 288216 389360
rect 240048 389240 240100 389292
rect 284208 389240 284260 389292
rect 297364 389240 297416 389292
rect 283472 389172 283524 389224
rect 293224 389172 293276 389224
rect 32496 389104 32548 389156
rect 272156 389104 272208 389156
rect 236552 389036 236604 389088
rect 295984 389036 296036 389088
rect 235816 388968 235868 389020
rect 300124 388968 300176 389020
rect 236920 388900 236972 388952
rect 302884 388900 302936 388952
rect 237656 388832 237708 388884
rect 313924 388832 313976 388884
rect 235448 388764 235500 388816
rect 318064 388764 318116 388816
rect 243636 388696 243688 388748
rect 443644 388696 443696 388748
rect 33876 388628 33928 388680
rect 270224 388628 270276 388680
rect 29644 388560 29696 388612
rect 273628 388560 273680 388612
rect 21456 388492 21508 388544
rect 272524 388492 272576 388544
rect 18696 388424 18748 388476
rect 271328 388424 271380 388476
rect 17316 388356 17368 388408
rect 270960 388356 271012 388408
rect 14648 388288 14700 388340
rect 269856 388288 269908 388340
rect 18604 388220 18656 388272
rect 276020 388220 276072 388272
rect 14556 388152 14608 388204
rect 273490 388152 273542 388204
rect 7564 388084 7616 388136
rect 268982 388084 269034 388136
rect 277998 388084 278050 388136
rect 447784 388084 447836 388136
rect 11796 388016 11848 388068
rect 274364 388016 274416 388068
rect 278596 388016 278648 388068
rect 449164 388016 449216 388068
rect 4804 387948 4856 388000
rect 275468 387948 275520 388000
rect 280528 387948 280580 388000
rect 481640 387948 481692 388000
rect 3424 387880 3476 387932
rect 276664 387880 276716 387932
rect 282000 387880 282052 387932
rect 485780 387880 485832 387932
rect 243268 387812 243320 387864
rect 537484 387812 537536 387864
rect 263600 387744 263652 387796
rect 263876 387744 263928 387796
rect 237288 387311 237340 387320
rect 237288 387277 237297 387311
rect 237297 387277 237331 387311
rect 237331 387277 237340 387311
rect 237288 387268 237340 387277
rect 238024 387311 238076 387320
rect 238024 387277 238033 387311
rect 238033 387277 238067 387311
rect 238067 387277 238076 387311
rect 238024 387268 238076 387277
rect 238668 387268 238720 387320
rect 239128 387311 239180 387320
rect 239128 387277 239137 387311
rect 239137 387277 239171 387311
rect 239171 387277 239180 387311
rect 239128 387268 239180 387277
rect 239956 387311 240008 387320
rect 239956 387277 239965 387311
rect 239965 387277 239999 387311
rect 239999 387277 240008 387311
rect 239956 387268 240008 387277
rect 241060 387311 241112 387320
rect 241060 387277 241069 387311
rect 241069 387277 241103 387311
rect 241103 387277 241112 387311
rect 241060 387268 241112 387277
rect 242164 387311 242216 387320
rect 242164 387277 242173 387311
rect 242173 387277 242207 387311
rect 242207 387277 242216 387311
rect 242164 387268 242216 387277
rect 244280 387311 244332 387320
rect 244280 387277 244289 387311
rect 244289 387277 244323 387311
rect 244323 387277 244332 387311
rect 244280 387268 244332 387277
rect 244832 387311 244884 387320
rect 244832 387277 244841 387311
rect 244841 387277 244875 387311
rect 244875 387277 244884 387311
rect 244832 387268 244884 387277
rect 269120 387311 269172 387320
rect 269120 387277 269129 387311
rect 269129 387277 269163 387311
rect 269163 387277 269172 387311
rect 269120 387268 269172 387277
rect 274732 387311 274784 387320
rect 274732 387277 274741 387311
rect 274741 387277 274775 387311
rect 274775 387277 274784 387311
rect 274732 387268 274784 387277
rect 283840 387311 283892 387320
rect 283840 387277 283849 387311
rect 283849 387277 283883 387311
rect 283883 387277 283892 387311
rect 283840 387268 283892 387277
rect 580356 387132 580408 387184
rect 17224 387064 17276 387116
rect 3516 386996 3568 387048
rect 288348 386996 288400 387048
rect 471244 386996 471296 387048
rect 555424 386928 555476 386980
rect 580908 386860 580960 386912
rect 580724 386792 580776 386844
rect 580816 386724 580868 386776
rect 580632 386656 580684 386708
rect 580448 386588 580500 386640
rect 580540 386520 580592 386572
rect 580264 386452 580316 386504
rect 293316 386384 293368 386436
rect 288348 385024 288400 385076
rect 298744 385024 298796 385076
rect 288348 383664 288400 383716
rect 468484 383664 468536 383716
rect 287428 381692 287480 381744
rect 294788 381692 294840 381744
rect 288348 379516 288400 379568
rect 465724 379516 465776 379568
rect 288348 378156 288400 378208
rect 297456 378156 297508 378208
rect 287428 376728 287480 376780
rect 293408 376728 293460 376780
rect 287612 375368 287664 375420
rect 293500 375368 293552 375420
rect 288348 374144 288400 374196
rect 293592 374144 293644 374196
rect 287796 371628 287848 371680
rect 292304 371628 292356 371680
rect 3332 371560 3384 371612
rect 7564 371560 7616 371612
rect 287612 370540 287664 370592
rect 290556 370540 290608 370592
rect 288348 368500 288400 368552
rect 446404 368500 446456 368552
rect 287980 367072 288032 367124
rect 297548 367072 297600 367124
rect 287612 365712 287664 365764
rect 296168 365712 296220 365764
rect 289084 365644 289136 365696
rect 580172 365644 580224 365696
rect 288348 364352 288400 364404
rect 296260 364352 296312 364404
rect 287612 362312 287664 362364
rect 296352 362312 296404 362364
rect 287612 360612 287664 360664
rect 296444 360612 296496 360664
rect 287612 358980 287664 359032
rect 289452 358980 289504 359032
rect 3332 358708 3384 358760
rect 15844 358708 15896 358760
rect 288348 357416 288400 357468
rect 474004 357416 474056 357468
rect 287796 356056 287848 356108
rect 298928 356056 298980 356108
rect 288348 354696 288400 354748
rect 298836 354696 298888 354748
rect 287520 351908 287572 351960
rect 472624 351908 472676 351960
rect 287244 351432 287296 351484
rect 294880 351432 294932 351484
rect 232136 349800 232188 349852
rect 232872 349800 232924 349852
rect 288348 349120 288400 349172
rect 467104 349120 467156 349172
rect 287980 347760 288032 347812
rect 299020 347760 299072 347812
rect 287980 346536 288032 346588
rect 294972 346536 295024 346588
rect 288348 345040 288400 345092
rect 295064 345040 295116 345092
rect 288348 342252 288400 342304
rect 464344 342252 464396 342304
rect 288348 340892 288400 340944
rect 297732 340892 297784 340944
rect 287796 339464 287848 339516
rect 292396 339464 292448 339516
rect 446404 338716 446456 338768
rect 488540 338716 488592 338768
rect 234528 338648 234580 338700
rect 467840 338648 467892 338700
rect 232136 338580 232188 338632
rect 297640 338580 297692 338632
rect 232872 338512 232924 338564
rect 289544 338512 289596 338564
rect 234620 338036 234672 338088
rect 233608 337968 233660 338020
rect 242716 337968 242768 338020
rect 234896 337900 234948 337952
rect 235310 337900 235362 337952
rect 235586 337900 235638 337952
rect 236322 337900 236374 337952
rect 237150 337900 237202 337952
rect 237702 337900 237754 337952
rect 237886 337900 237938 337952
rect 238622 337900 238674 337952
rect 238714 337900 238766 337952
rect 238898 337900 238950 337952
rect 239266 337900 239318 337952
rect 239358 337900 239410 337952
rect 239542 337900 239594 337952
rect 239726 337900 239778 337952
rect 241106 337900 241158 337952
rect 241382 337900 241434 337952
rect 242394 337900 242446 337952
rect 243130 337900 243182 337952
rect 245338 337900 245390 337952
rect 245522 337900 245574 337952
rect 248282 337900 248334 337952
rect 248512 337943 248564 337952
rect 248512 337909 248521 337943
rect 248521 337909 248555 337943
rect 248555 337909 248564 337943
rect 248512 337900 248564 337909
rect 235494 337832 235546 337884
rect 235862 337832 235914 337884
rect 237334 337832 237386 337884
rect 238070 337832 238122 337884
rect 238346 337832 238398 337884
rect 238438 337832 238490 337884
rect 235678 337764 235730 337816
rect 236506 337764 236558 337816
rect 236598 337764 236650 337816
rect 237518 337764 237570 337816
rect 239910 337832 239962 337884
rect 240278 337832 240330 337884
rect 240554 337832 240606 337884
rect 241658 337832 241710 337884
rect 242302 337832 242354 337884
rect 243038 337832 243090 337884
rect 243222 337832 243274 337884
rect 243590 337832 243642 337884
rect 243774 337832 243826 337884
rect 244234 337832 244286 337884
rect 244556 337832 244608 337884
rect 245062 337832 245114 337884
rect 245890 337832 245942 337884
rect 246718 337832 246770 337884
rect 246902 337832 246954 337884
rect 247178 337832 247230 337884
rect 248098 337832 248150 337884
rect 249478 337900 249530 337952
rect 249846 337900 249898 337952
rect 250766 337900 250818 337952
rect 251134 337900 251186 337952
rect 251226 337900 251278 337952
rect 251410 337900 251462 337952
rect 251502 337900 251554 337952
rect 251686 337900 251738 337952
rect 252514 337900 252566 337952
rect 253250 337900 253302 337952
rect 253526 337900 253578 337952
rect 253802 337900 253854 337952
rect 254630 337900 254682 337952
rect 254814 337900 254866 337952
rect 248834 337832 248886 337884
rect 248926 337832 248978 337884
rect 249294 337832 249346 337884
rect 249662 337832 249714 337884
rect 250122 337832 250174 337884
rect 238668 337764 238720 337816
rect 238760 337764 238812 337816
rect 239082 337764 239134 337816
rect 239772 337764 239824 337816
rect 242440 337764 242492 337816
rect 244970 337764 245022 337816
rect 245430 337764 245482 337816
rect 252790 337832 252842 337884
rect 253894 337832 253946 337884
rect 254446 337832 254498 337884
rect 250674 337764 250726 337816
rect 250950 337764 251002 337816
rect 251180 337764 251232 337816
rect 251870 337764 251922 337816
rect 253434 337764 253486 337816
rect 253710 337764 253762 337816
rect 255090 337900 255142 337952
rect 255366 337900 255418 337952
rect 255642 337900 255694 337952
rect 255918 337900 255970 337952
rect 256470 337900 256522 337952
rect 257114 337900 257166 337952
rect 257298 337900 257350 337952
rect 257482 337900 257534 337952
rect 257574 337900 257626 337952
rect 257850 337900 257902 337952
rect 258678 337900 258730 337952
rect 258862 337900 258914 337952
rect 259230 337900 259282 337952
rect 259414 337900 259466 337952
rect 259598 337900 259650 337952
rect 260058 337900 260110 337952
rect 260334 337900 260386 337952
rect 261254 337900 261306 337952
rect 262266 337900 262318 337952
rect 262450 337900 262502 337952
rect 262542 337900 262594 337952
rect 264198 337900 264250 337952
rect 264750 337900 264802 337952
rect 264934 337900 264986 337952
rect 265026 337900 265078 337952
rect 265210 337900 265262 337952
rect 265394 337900 265446 337952
rect 266498 337900 266550 337952
rect 266682 337900 266734 337952
rect 266774 337900 266826 337952
rect 267326 337900 267378 337952
rect 268338 337900 268390 337952
rect 268614 337900 268666 337952
rect 269074 337900 269126 337952
rect 269350 337900 269402 337952
rect 270454 337900 270506 337952
rect 270546 337900 270598 337952
rect 272202 337900 272254 337952
rect 272386 337900 272438 337952
rect 272754 337900 272806 337952
rect 274226 337900 274278 337952
rect 274870 337900 274922 337952
rect 275146 337900 275198 337952
rect 275974 337900 276026 337952
rect 276158 337900 276210 337952
rect 276434 337900 276486 337952
rect 277078 337900 277130 337952
rect 278090 337900 278142 337952
rect 278366 337900 278418 337952
rect 278734 337900 278786 337952
rect 287428 338104 287480 338156
rect 296536 338104 296588 338156
rect 279102 337900 279154 337952
rect 281310 337900 281362 337952
rect 281678 337900 281730 337952
rect 281862 337900 281914 337952
rect 282138 337900 282190 337952
rect 282414 337900 282466 337952
rect 282506 337900 282558 337952
rect 254998 337832 255050 337884
rect 255550 337832 255602 337884
rect 256286 337832 256338 337884
rect 256654 337832 256706 337884
rect 257022 337832 257074 337884
rect 258494 337832 258546 337884
rect 258770 337832 258822 337884
rect 260610 337832 260662 337884
rect 261162 337832 261214 337884
rect 261438 337832 261490 337884
rect 262174 337832 262226 337884
rect 262634 337832 262686 337884
rect 262818 337832 262870 337884
rect 263094 337832 263146 337884
rect 263646 337832 263698 337884
rect 264382 337832 264434 337884
rect 266958 337832 267010 337884
rect 267234 337832 267286 337884
rect 267878 337832 267930 337884
rect 268154 337832 268206 337884
rect 255412 337764 255464 337816
rect 255964 337764 256016 337816
rect 257206 337764 257258 337816
rect 258310 337764 258362 337816
rect 260886 337764 260938 337816
rect 268430 337764 268482 337816
rect 268798 337832 268850 337884
rect 268982 337832 269034 337884
rect 269902 337832 269954 337884
rect 270178 337832 270230 337884
rect 271006 337832 271058 337884
rect 271374 337832 271426 337884
rect 271512 337875 271564 337884
rect 271512 337841 271521 337875
rect 271521 337841 271555 337875
rect 271555 337841 271564 337875
rect 271512 337832 271564 337841
rect 271650 337832 271702 337884
rect 272846 337832 272898 337884
rect 273766 337832 273818 337884
rect 273950 337832 274002 337884
rect 274134 337832 274186 337884
rect 275790 337832 275842 337884
rect 276342 337832 276394 337884
rect 277722 337832 277774 337884
rect 277998 337832 278050 337884
rect 279562 337832 279614 337884
rect 280114 337832 280166 337884
rect 280206 337832 280258 337884
rect 280574 337832 280626 337884
rect 280850 337832 280902 337884
rect 285220 337968 285272 338020
rect 283886 337900 283938 337952
rect 284070 337900 284122 337952
rect 288256 337900 288308 337952
rect 284254 337832 284306 337884
rect 278918 337764 278970 337816
rect 436744 337696 436796 337748
rect 232320 337492 232372 337544
rect 479524 337628 479576 337680
rect 235448 337603 235500 337612
rect 235448 337569 235457 337603
rect 235457 337569 235491 337603
rect 235491 337569 235500 337603
rect 235448 337560 235500 337569
rect 235632 337603 235684 337612
rect 235632 337569 235641 337603
rect 235641 337569 235675 337603
rect 235675 337569 235684 337603
rect 235632 337560 235684 337569
rect 237840 337560 237892 337612
rect 238024 337603 238076 337612
rect 238024 337569 238033 337603
rect 238033 337569 238067 337603
rect 238067 337569 238076 337603
rect 238024 337560 238076 337569
rect 238576 337560 238628 337612
rect 239312 337560 239364 337612
rect 483020 337560 483072 337612
rect 234988 337492 235040 337544
rect 241152 337492 241204 337544
rect 243360 337535 243412 337544
rect 243360 337501 243369 337535
rect 243369 337501 243403 337535
rect 243403 337501 243412 337535
rect 243360 337492 243412 337501
rect 244004 337535 244056 337544
rect 244004 337501 244013 337535
rect 244013 337501 244047 337535
rect 244047 337501 244056 337535
rect 244004 337492 244056 337501
rect 246120 337535 246172 337544
rect 246120 337501 246129 337535
rect 246129 337501 246163 337535
rect 246163 337501 246172 337535
rect 246120 337492 246172 337501
rect 246856 337535 246908 337544
rect 246856 337501 246865 337535
rect 246865 337501 246899 337535
rect 246899 337501 246908 337535
rect 246856 337492 246908 337501
rect 247040 337535 247092 337544
rect 247040 337501 247049 337535
rect 247049 337501 247083 337535
rect 247083 337501 247092 337535
rect 247040 337492 247092 337501
rect 249064 337535 249116 337544
rect 249064 337501 249073 337535
rect 249073 337501 249107 337535
rect 249107 337501 249116 337535
rect 249064 337492 249116 337501
rect 253112 337535 253164 337544
rect 253112 337501 253121 337535
rect 253121 337501 253155 337535
rect 253155 337501 253164 337535
rect 253112 337492 253164 337501
rect 253296 337535 253348 337544
rect 253296 337501 253305 337535
rect 253305 337501 253339 337535
rect 253339 337501 253348 337535
rect 253296 337492 253348 337501
rect 253756 337535 253808 337544
rect 253756 337501 253765 337535
rect 253765 337501 253799 337535
rect 253799 337501 253808 337535
rect 253756 337492 253808 337501
rect 254860 337492 254912 337544
rect 256424 337492 256476 337544
rect 257712 337492 257764 337544
rect 258632 337492 258684 337544
rect 260564 337492 260616 337544
rect 262772 337492 262824 337544
rect 262956 337535 263008 337544
rect 262956 337501 262965 337535
rect 262965 337501 262999 337535
rect 262999 337501 263008 337535
rect 262956 337492 263008 337501
rect 265440 337535 265492 337544
rect 265440 337501 265449 337535
rect 265449 337501 265483 337535
rect 265483 337501 265492 337535
rect 265440 337492 265492 337501
rect 268016 337535 268068 337544
rect 268016 337501 268025 337535
rect 268025 337501 268059 337535
rect 268059 337501 268068 337535
rect 268016 337492 268068 337501
rect 269764 337535 269816 337544
rect 269764 337501 269773 337535
rect 269773 337501 269807 337535
rect 269807 337501 269816 337535
rect 269764 337492 269816 337501
rect 270316 337535 270368 337544
rect 270316 337501 270325 337535
rect 270325 337501 270359 337535
rect 270359 337501 270368 337535
rect 270316 337492 270368 337501
rect 271328 337535 271380 337544
rect 271328 337501 271337 337535
rect 271337 337501 271371 337535
rect 271371 337501 271380 337535
rect 271328 337492 271380 337501
rect 271880 337535 271932 337544
rect 271880 337501 271889 337535
rect 271889 337501 271923 337535
rect 271923 337501 271932 337535
rect 271880 337492 271932 337501
rect 275284 337492 275336 337544
rect 275744 337492 275796 337544
rect 276388 337492 276440 337544
rect 277124 337492 277176 337544
rect 278320 337535 278372 337544
rect 278320 337501 278329 337535
rect 278329 337501 278363 337535
rect 278363 337501 278372 337535
rect 278320 337492 278372 337501
rect 282368 337492 282420 337544
rect 282920 337492 282972 337544
rect 284116 337492 284168 337544
rect 285036 337492 285088 337544
rect 580908 337492 580960 337544
rect 234712 337424 234764 337476
rect 530676 337424 530728 337476
rect 233516 337356 233568 337408
rect 538312 337356 538364 337408
rect 232504 337288 232556 337340
rect 250904 337288 250956 337340
rect 251088 337288 251140 337340
rect 254400 337288 254452 337340
rect 254860 337288 254912 337340
rect 254952 337288 255004 337340
rect 255596 337288 255648 337340
rect 275652 337288 275704 337340
rect 278136 337331 278188 337340
rect 278136 337297 278145 337331
rect 278145 337297 278179 337331
rect 278179 337297 278188 337331
rect 278136 337288 278188 337297
rect 278964 337288 279016 337340
rect 236184 337263 236236 337272
rect 236184 337229 236193 337263
rect 236193 337229 236227 337263
rect 236227 337229 236236 337263
rect 236184 337220 236236 337229
rect 237564 337220 237616 337272
rect 420920 337220 420972 337272
rect 254768 337152 254820 337204
rect 266912 337152 266964 337204
rect 269304 337152 269356 337204
rect 273536 337152 273588 337204
rect 278596 337084 278648 337136
rect 536840 337152 536892 337204
rect 279148 337016 279200 337068
rect 279332 337016 279384 337068
rect 279516 337084 279568 337136
rect 538220 337084 538272 337136
rect 282920 337059 282972 337068
rect 282920 337025 282929 337059
rect 282929 337025 282963 337059
rect 282963 337025 282972 337059
rect 282920 337016 282972 337025
rect 283288 337016 283340 337068
rect 283656 337016 283708 337068
rect 242716 336948 242768 337000
rect 265072 336948 265124 337000
rect 276296 336948 276348 337000
rect 276756 336948 276808 337000
rect 276940 336948 276992 337000
rect 538864 337016 538916 337068
rect 287612 336948 287664 337000
rect 538956 336948 539008 337000
rect 33140 336744 33192 336796
rect 237840 336880 237892 336932
rect 243912 336880 243964 336932
rect 264612 336880 264664 336932
rect 275376 336880 275428 336932
rect 283012 336880 283064 336932
rect 543740 336880 543792 336932
rect 237380 336812 237432 336864
rect 269212 336812 269264 336864
rect 240416 336744 240468 336796
rect 240692 336744 240744 336796
rect 241612 336787 241664 336796
rect 241612 336753 241621 336787
rect 241621 336753 241655 336787
rect 241655 336753 241664 336787
rect 241612 336744 241664 336753
rect 267004 336744 267056 336796
rect 103428 336676 103480 336728
rect 240140 336676 240192 336728
rect 247776 336676 247828 336728
rect 263324 336676 263376 336728
rect 266268 336676 266320 336728
rect 275100 336812 275152 336864
rect 277400 336855 277452 336864
rect 277400 336821 277409 336855
rect 277409 336821 277443 336855
rect 277443 336821 277452 336855
rect 277400 336812 277452 336821
rect 279608 336812 279660 336864
rect 557540 336812 557592 336864
rect 274272 336744 274324 336796
rect 274732 336744 274784 336796
rect 279516 336744 279568 336796
rect 561680 336744 561732 336796
rect 341524 336676 341576 336728
rect 96528 336608 96580 336660
rect 242808 336608 242860 336660
rect 249064 336608 249116 336660
rect 254124 336608 254176 336660
rect 259276 336608 259328 336660
rect 263968 336608 264020 336660
rect 268108 336608 268160 336660
rect 95148 336540 95200 336592
rect 259920 336540 259972 336592
rect 344284 336608 344336 336660
rect 46848 336472 46900 336524
rect 78588 336404 78640 336456
rect 243452 336472 243504 336524
rect 267464 336472 267516 336524
rect 348424 336540 348476 336592
rect 45468 336336 45520 336388
rect 238852 336336 238904 336388
rect 240232 336336 240284 336388
rect 240692 336404 240744 336456
rect 244188 336404 244240 336456
rect 263416 336404 263468 336456
rect 355324 336472 355376 336524
rect 362224 336404 362276 336456
rect 243452 336336 243504 336388
rect 261116 336336 261168 336388
rect 89628 336268 89680 336320
rect 64788 336200 64840 336252
rect 261668 336268 261720 336320
rect 264244 336268 264296 336320
rect 267740 336268 267792 336320
rect 268384 336268 268436 336320
rect 369124 336336 369176 336388
rect 376024 336268 376076 336320
rect 237840 336200 237892 336252
rect 240232 336200 240284 336252
rect 248696 336200 248748 336252
rect 260840 336200 260892 336252
rect 262220 336200 262272 336252
rect 263508 336200 263560 336252
rect 265716 336200 265768 336252
rect 39948 336132 40000 336184
rect 238116 336132 238168 336184
rect 238208 336132 238260 336184
rect 243728 336132 243780 336184
rect 261944 336132 261996 336184
rect 267280 336132 267332 336184
rect 24768 336064 24820 336116
rect 236920 336064 236972 336116
rect 238760 336064 238812 336116
rect 260288 336064 260340 336116
rect 233608 335996 233660 336048
rect 242256 335996 242308 336048
rect 242808 335996 242860 336048
rect 256792 335996 256844 336048
rect 117228 335928 117280 335980
rect 244464 335928 244516 335980
rect 250628 335928 250680 335980
rect 262036 335971 262088 335980
rect 262036 335937 262045 335971
rect 262045 335937 262079 335971
rect 262079 335937 262088 335971
rect 262036 335928 262088 335937
rect 119988 335860 120040 335912
rect 239128 335860 239180 335912
rect 251548 335860 251600 335912
rect 255964 335860 256016 335912
rect 259460 335860 259512 335912
rect 262956 336064 263008 336116
rect 269396 336200 269448 336252
rect 270316 336200 270368 336252
rect 382924 336200 382976 336252
rect 391204 336132 391256 336184
rect 267740 335996 267792 336048
rect 269488 335996 269540 336048
rect 279424 336064 279476 336116
rect 405004 336064 405056 336116
rect 171784 335792 171836 335844
rect 248144 335792 248196 335844
rect 256148 335792 256200 335844
rect 258724 335792 258776 335844
rect 262956 335792 263008 335844
rect 263232 335792 263284 335844
rect 264980 335860 265032 335912
rect 268476 335860 268528 335912
rect 269672 335860 269724 335912
rect 270316 335860 270368 335912
rect 271972 335928 272024 335980
rect 272524 335928 272576 335980
rect 407764 335996 407816 336048
rect 337384 335928 337436 335980
rect 274732 335860 274784 335912
rect 275928 335860 275980 335912
rect 277400 335860 277452 335912
rect 278504 335860 278556 335912
rect 280344 335860 280396 335912
rect 283288 335860 283340 335912
rect 264520 335792 264572 335844
rect 178684 335724 178736 335776
rect 239036 335724 239088 335776
rect 245292 335724 245344 335776
rect 257252 335724 257304 335776
rect 257896 335724 257948 335776
rect 269856 335792 269908 335844
rect 273904 335792 273956 335844
rect 274180 335792 274232 335844
rect 180064 335656 180116 335708
rect 244924 335656 244976 335708
rect 251272 335656 251324 335708
rect 259552 335656 259604 335708
rect 261116 335656 261168 335708
rect 283196 335792 283248 335844
rect 283472 335792 283524 335844
rect 344560 335860 344612 335912
rect 344468 335792 344520 335844
rect 280804 335724 280856 335776
rect 282000 335724 282052 335776
rect 282828 335724 282880 335776
rect 344376 335724 344428 335776
rect 316684 335656 316736 335708
rect 231124 335588 231176 335640
rect 236828 335588 236880 335640
rect 243820 335588 243872 335640
rect 240416 335520 240468 335572
rect 257896 335631 257948 335640
rect 257896 335597 257905 335631
rect 257905 335597 257939 335631
rect 257939 335597 257948 335631
rect 257896 335588 257948 335597
rect 260748 335588 260800 335640
rect 232872 335452 232924 335504
rect 231216 335384 231268 335436
rect 234988 335384 235040 335436
rect 237932 335452 237984 335504
rect 242164 335452 242216 335504
rect 243360 335452 243412 335504
rect 242072 335384 242124 335436
rect 242256 335384 242308 335436
rect 247224 335520 247276 335572
rect 244188 335452 244240 335504
rect 260564 335452 260616 335504
rect 260748 335452 260800 335504
rect 244464 335384 244516 335436
rect 6828 335316 6880 335368
rect 238024 335316 238076 335368
rect 241244 335316 241296 335368
rect 255688 335316 255740 335368
rect 256884 335316 256936 335368
rect 257344 335316 257396 335368
rect 260380 335316 260432 335368
rect 260564 335316 260616 335368
rect 261024 335316 261076 335368
rect 261484 335316 261536 335368
rect 261760 335316 261812 335368
rect 261944 335316 261996 335368
rect 262404 335588 262456 335640
rect 263140 335588 263192 335640
rect 300216 335588 300268 335640
rect 271972 335520 272024 335572
rect 274456 335520 274508 335572
rect 274824 335520 274876 335572
rect 275468 335520 275520 335572
rect 277952 335520 278004 335572
rect 278504 335520 278556 335572
rect 281816 335520 281868 335572
rect 282552 335520 282604 335572
rect 283472 335563 283524 335572
rect 283472 335529 283481 335563
rect 283481 335529 283515 335563
rect 283515 335529 283524 335563
rect 283472 335520 283524 335529
rect 283748 335520 283800 335572
rect 268108 335452 268160 335504
rect 269764 335452 269816 335504
rect 272064 335452 272116 335504
rect 272800 335452 272852 335504
rect 273904 335452 273956 335504
rect 274548 335452 274600 335504
rect 281356 335495 281408 335504
rect 281356 335461 281365 335495
rect 281365 335461 281399 335495
rect 281399 335461 281408 335495
rect 281356 335452 281408 335461
rect 282000 335495 282052 335504
rect 282000 335461 282009 335495
rect 282009 335461 282043 335495
rect 282043 335461 282052 335495
rect 282000 335452 282052 335461
rect 282092 335452 282144 335504
rect 282644 335452 282696 335504
rect 262864 335384 262916 335436
rect 263324 335384 263376 335436
rect 263784 335384 263836 335436
rect 270684 335384 270736 335436
rect 271788 335384 271840 335436
rect 201408 335248 201460 335300
rect 244188 335248 244240 335300
rect 245016 335248 245068 335300
rect 254216 335248 254268 335300
rect 263876 335316 263928 335368
rect 264336 335316 264388 335368
rect 267740 335316 267792 335368
rect 267924 335316 267976 335368
rect 269948 335316 270000 335368
rect 270408 335316 270460 335368
rect 274732 335316 274784 335368
rect 274916 335316 274968 335368
rect 275468 335359 275520 335368
rect 275468 335325 275477 335359
rect 275477 335325 275511 335359
rect 275511 335325 275520 335359
rect 275468 335316 275520 335325
rect 275560 335316 275612 335368
rect 275744 335316 275796 335368
rect 277400 335316 277452 335368
rect 277768 335316 277820 335368
rect 277952 335316 278004 335368
rect 278228 335384 278280 335436
rect 278412 335384 278464 335436
rect 283564 335384 283616 335436
rect 284024 335384 284076 335436
rect 262588 335248 262640 335300
rect 268752 335248 268804 335300
rect 208308 335180 208360 335232
rect 282276 335248 282328 335300
rect 282552 335291 282604 335300
rect 282552 335257 282561 335291
rect 282561 335257 282595 335291
rect 282595 335257 282604 335291
rect 282552 335248 282604 335257
rect 197268 335112 197320 335164
rect 250996 335112 251048 335164
rect 282644 335180 282696 335232
rect 194508 335044 194560 335096
rect 251272 335044 251324 335096
rect 255136 335044 255188 335096
rect 261760 335087 261812 335096
rect 261760 335053 261769 335087
rect 261769 335053 261803 335087
rect 261803 335053 261812 335087
rect 261760 335044 261812 335053
rect 190368 334976 190420 335028
rect 250444 334976 250496 335028
rect 183468 334908 183520 334960
rect 243268 334908 243320 334960
rect 244004 334908 244056 334960
rect 245476 334951 245528 334960
rect 245476 334917 245485 334951
rect 245485 334917 245519 334951
rect 245519 334917 245528 334951
rect 245476 334908 245528 334917
rect 186228 334840 186280 334892
rect 252744 334840 252796 334892
rect 253296 334840 253348 334892
rect 284116 335316 284168 335368
rect 284300 335452 284352 335504
rect 285404 335452 285456 335504
rect 284576 335384 284628 335436
rect 285312 335384 285364 335436
rect 284668 335316 284720 335368
rect 284852 335316 284904 335368
rect 285036 335248 285088 335300
rect 285128 335180 285180 335232
rect 288440 335180 288492 335232
rect 286416 335112 286468 335164
rect 179328 334772 179380 334824
rect 249524 334772 249576 334824
rect 258816 334772 258868 334824
rect 283012 335044 283064 335096
rect 289360 335044 289412 335096
rect 273720 335019 273772 335028
rect 273720 334985 273729 335019
rect 273729 334985 273763 335019
rect 273763 334985 273772 335019
rect 273720 334976 273772 334985
rect 316040 334976 316092 335028
rect 369860 334908 369912 334960
rect 277032 334840 277084 334892
rect 401600 334840 401652 334892
rect 271788 334815 271840 334824
rect 271788 334781 271797 334815
rect 271797 334781 271831 334815
rect 271831 334781 271840 334815
rect 271788 334772 271840 334781
rect 271972 334772 272024 334824
rect 415492 334772 415544 334824
rect 169668 334704 169720 334756
rect 240232 334704 240284 334756
rect 248328 334704 248380 334756
rect 272524 334704 272576 334756
rect 438124 334704 438176 334756
rect 176568 334636 176620 334688
rect 248972 334636 249024 334688
rect 260012 334636 260064 334688
rect 265532 334636 265584 334688
rect 374000 334636 374052 334688
rect 395344 334636 395396 334688
rect 580724 334636 580776 334688
rect 165528 334568 165580 334620
rect 238760 334568 238812 334620
rect 240416 334611 240468 334620
rect 240416 334577 240425 334611
rect 240425 334577 240459 334611
rect 240459 334577 240468 334611
rect 240416 334568 240468 334577
rect 240876 334568 240928 334620
rect 241244 334568 241296 334620
rect 243544 334568 243596 334620
rect 243728 334568 243780 334620
rect 244648 334568 244700 334620
rect 245200 334568 245252 334620
rect 251824 334568 251876 334620
rect 252100 334568 252152 334620
rect 254308 334611 254360 334620
rect 254308 334577 254317 334611
rect 254317 334577 254351 334611
rect 254351 334577 254360 334611
rect 254308 334568 254360 334577
rect 274640 334568 274692 334620
rect 280988 334568 281040 334620
rect 554780 334568 554832 334620
rect 204168 334500 204220 334552
rect 244464 334500 244516 334552
rect 265900 334500 265952 334552
rect 276296 334500 276348 334552
rect 283196 334500 283248 334552
rect 286600 334500 286652 334552
rect 210976 334432 211028 334484
rect 252192 334432 252244 334484
rect 215208 334364 215260 334416
rect 272156 334364 272208 334416
rect 272892 334364 272944 334416
rect 276940 334364 276992 334416
rect 222108 334296 222160 334348
rect 253020 334296 253072 334348
rect 287888 334432 287940 334484
rect 289268 334364 289320 334416
rect 226248 334228 226300 334280
rect 253388 334228 253440 334280
rect 269672 334228 269724 334280
rect 229008 334160 229060 334212
rect 253572 334160 253624 334212
rect 275376 334228 275428 334280
rect 289084 334296 289136 334348
rect 289176 334228 289228 334280
rect 282276 334160 282328 334212
rect 282368 334160 282420 334212
rect 219348 334092 219400 334144
rect 239128 334092 239180 334144
rect 240048 334092 240100 334144
rect 240692 334092 240744 334144
rect 240968 334092 241020 334144
rect 242072 334092 242124 334144
rect 242532 334092 242584 334144
rect 243820 334092 243872 334144
rect 245200 334135 245252 334144
rect 245200 334101 245209 334135
rect 245209 334101 245243 334135
rect 245243 334101 245252 334135
rect 245200 334092 245252 334101
rect 272708 334092 272760 334144
rect 276020 334092 276072 334144
rect 278596 334092 278648 334144
rect 285588 334160 285640 334212
rect 287980 334160 288032 334212
rect 287796 334092 287848 334144
rect 231400 334024 231452 334076
rect 248880 334024 248932 334076
rect 250352 334024 250404 334076
rect 254676 334024 254728 334076
rect 268752 334024 268804 334076
rect 282368 334024 282420 334076
rect 287704 334024 287756 334076
rect 232504 333956 232556 334008
rect 250536 333956 250588 334008
rect 254492 333956 254544 334008
rect 271420 333956 271472 334008
rect 278044 333956 278096 334008
rect 282920 333956 282972 334008
rect 284392 333956 284444 334008
rect 290648 333956 290700 334008
rect 180708 333888 180760 333940
rect 258816 333888 258868 333940
rect 264796 333888 264848 333940
rect 362960 333888 363012 333940
rect 177948 333820 178000 333872
rect 249432 333820 249484 333872
rect 365720 333820 365772 333872
rect 173808 333752 173860 333804
rect 249156 333752 249208 333804
rect 265716 333752 265768 333804
rect 376760 333752 376812 333804
rect 169576 333684 169628 333736
rect 266084 333684 266136 333736
rect 380900 333684 380952 333736
rect 166908 333616 166960 333668
rect 387800 333616 387852 333668
rect 162768 333548 162820 333600
rect 244924 333548 244976 333600
rect 245752 333548 245804 333600
rect 266452 333548 266504 333600
rect 383660 333548 383712 333600
rect 151728 333480 151780 333532
rect 242256 333480 242308 333532
rect 247132 333480 247184 333532
rect 390652 333480 390704 333532
rect 154488 333412 154540 333464
rect 247500 333412 247552 333464
rect 394700 333412 394752 333464
rect 148968 333344 149020 333396
rect 147588 333276 147640 333328
rect 245936 333344 245988 333396
rect 253388 333344 253440 333396
rect 255320 333344 255372 333396
rect 267556 333344 267608 333396
rect 398840 333344 398892 333396
rect 253940 333276 253992 333328
rect 256976 333276 257028 333328
rect 257988 333276 258040 333328
rect 264428 333276 264480 333328
rect 405740 333276 405792 333328
rect 131028 333208 131080 333260
rect 245568 333208 245620 333260
rect 252928 333208 252980 333260
rect 255228 333251 255280 333260
rect 255228 333217 255237 333251
rect 255237 333217 255271 333251
rect 255271 333217 255280 333251
rect 255228 333208 255280 333217
rect 256056 333208 256108 333260
rect 256608 333208 256660 333260
rect 264704 333208 264756 333260
rect 408500 333208 408552 333260
rect 184848 333140 184900 333192
rect 249892 333140 249944 333192
rect 251916 333140 251968 333192
rect 254952 333140 255004 333192
rect 257068 333140 257120 333192
rect 259552 333140 259604 333192
rect 261208 333140 261260 333192
rect 262864 333140 262916 333192
rect 263692 333140 263744 333192
rect 358820 333140 358872 333192
rect 187608 333072 187660 333124
rect 250168 333072 250220 333124
rect 356060 333072 356112 333124
rect 191748 333004 191800 333056
rect 250444 333004 250496 333056
rect 320180 333004 320232 333056
rect 194416 332936 194468 332988
rect 250812 332936 250864 332988
rect 263232 332936 263284 332988
rect 264152 332936 264204 332988
rect 351920 332936 351972 332988
rect 202788 332868 202840 332920
rect 309140 332868 309192 332920
rect 205548 332800 205600 332852
rect 260748 332800 260800 332852
rect 306380 332800 306432 332852
rect 216588 332732 216640 332784
rect 252560 332732 252612 332784
rect 259736 332732 259788 332784
rect 302240 332732 302292 332784
rect 219256 332664 219308 332716
rect 249156 332664 249208 332716
rect 254216 332664 254268 332716
rect 299480 332664 299532 332716
rect 234528 332596 234580 332648
rect 249984 332596 250036 332648
rect 254860 332596 254912 332648
rect 271052 332596 271104 332648
rect 272340 332596 272392 332648
rect 272892 332596 272944 332648
rect 276480 332596 276532 332648
rect 277216 332596 277268 332648
rect 279608 332596 279660 332648
rect 283564 332596 283616 332648
rect 283748 332596 283800 332648
rect 283932 332596 283984 332648
rect 284116 332596 284168 332648
rect 286692 332596 286744 332648
rect 160008 332528 160060 332580
rect 247960 332528 248012 332580
rect 252468 332528 252520 332580
rect 255412 332528 255464 332580
rect 269488 332528 269540 332580
rect 429844 332528 429896 332580
rect 155868 332460 155920 332512
rect 247684 332460 247736 332512
rect 269396 332460 269448 332512
rect 430580 332460 430632 332512
rect 153108 332392 153160 332444
rect 247408 332392 247460 332444
rect 272984 332392 273036 332444
rect 276388 332392 276440 332444
rect 276572 332392 276624 332444
rect 434720 332392 434772 332444
rect 144828 332324 144880 332376
rect 246764 332324 246816 332376
rect 439596 332324 439648 332376
rect 142068 332256 142120 332308
rect 246488 332256 246540 332308
rect 256792 332256 256844 332308
rect 137928 332188 137980 332240
rect 246212 332188 246264 332240
rect 436836 332256 436888 332308
rect 276940 332188 276992 332240
rect 536932 332188 536984 332240
rect 135168 332120 135220 332172
rect 274180 332120 274232 332172
rect 279608 332120 279660 332172
rect 282368 332120 282420 332172
rect 128176 332052 128228 332104
rect 276848 332052 276900 332104
rect 279240 332052 279292 332104
rect 540336 332120 540388 332172
rect 543004 332052 543056 332104
rect 230388 331984 230440 332036
rect 274180 331984 274232 332036
rect 279332 331984 279384 332036
rect 547144 331984 547196 332036
rect 88248 331916 88300 331968
rect 232872 331916 232924 331968
rect 234712 331916 234764 331968
rect 235816 331916 235868 331968
rect 236460 331916 236512 331968
rect 238116 331916 238168 331968
rect 239404 331916 239456 331968
rect 279240 331959 279292 331968
rect 279240 331925 279249 331959
rect 279249 331925 279283 331959
rect 279283 331925 279292 331959
rect 279240 331916 279292 331925
rect 548524 331916 548576 331968
rect 43536 331848 43588 331900
rect 237840 331848 237892 331900
rect 164148 331780 164200 331832
rect 260840 331848 260892 331900
rect 280160 331848 280212 331900
rect 286876 331848 286928 331900
rect 556160 331848 556212 331900
rect 239496 331823 239548 331832
rect 239496 331789 239505 331823
rect 239505 331789 239539 331823
rect 239539 331789 239548 331823
rect 239496 331780 239548 331789
rect 246304 331780 246356 331832
rect 265348 331780 265400 331832
rect 371240 331780 371292 331832
rect 168288 331712 168340 331764
rect 248512 331712 248564 331764
rect 367100 331712 367152 331764
rect 186136 331644 186188 331696
rect 249892 331644 249944 331696
rect 259644 331644 259696 331696
rect 299572 331644 299624 331696
rect 200028 331576 200080 331628
rect 251180 331576 251232 331628
rect 261116 331576 261168 331628
rect 298100 331576 298152 331628
rect 212448 331508 212500 331560
rect 252284 331508 252336 331560
rect 217968 331440 218020 331492
rect 252652 331440 252704 331492
rect 263508 331440 263560 331492
rect 289820 331440 289872 331492
rect 223488 331372 223540 331424
rect 253204 331372 253256 331424
rect 258448 331372 258500 331424
rect 285680 331372 285732 331424
rect 291200 331372 291252 331424
rect 227628 331304 227680 331356
rect 110328 331236 110380 331288
rect 233608 331236 233660 331288
rect 237288 331304 237340 331356
rect 238944 331304 238996 331356
rect 239864 331304 239916 331356
rect 240692 331304 240744 331356
rect 294604 331304 294656 331356
rect 252744 331236 252796 331288
rect 253204 331236 253256 331288
rect 258264 331236 258316 331288
rect 278780 331236 278832 331288
rect 175188 331168 175240 331220
rect 249340 331168 249392 331220
rect 265624 331168 265676 331220
rect 374092 331168 374144 331220
rect 171048 331100 171100 331152
rect 378140 331100 378192 331152
rect 157248 331032 157300 331084
rect 247592 331032 247644 331084
rect 266176 331032 266228 331084
rect 382372 331032 382424 331084
rect 153016 330964 153068 331016
rect 247316 330964 247368 331016
rect 385040 330964 385092 331016
rect 150348 330896 150400 330948
rect 247040 330896 247092 330948
rect 256700 330896 256752 330948
rect 266360 330896 266412 330948
rect 389180 330896 389232 330948
rect 143448 330828 143500 330880
rect 246672 330828 246724 330880
rect 267096 330828 267148 330880
rect 391940 330828 391992 330880
rect 139308 330760 139360 330812
rect 243176 330760 243228 330812
rect 396080 330760 396132 330812
rect 132408 330692 132460 330744
rect 245660 330692 245712 330744
rect 267648 330692 267700 330744
rect 398932 330692 398984 330744
rect 102048 330624 102100 330676
rect 84108 330556 84160 330608
rect 241704 330556 241756 330608
rect 268660 330556 268712 330608
rect 402980 330624 403032 330676
rect 73068 330488 73120 330540
rect 241244 330488 241296 330540
rect 177856 330420 177908 330472
rect 268292 330488 268344 330540
rect 407212 330556 407264 330608
rect 409880 330488 409932 330540
rect 364340 330420 364392 330472
rect 188988 330352 189040 330404
rect 250260 330352 250312 330404
rect 264612 330352 264664 330404
rect 360200 330352 360252 330404
rect 193128 330284 193180 330336
rect 357440 330284 357492 330336
rect 202696 330216 202748 330268
rect 264336 330216 264388 330268
rect 353300 330216 353352 330268
rect 206928 330148 206980 330200
rect 252100 330148 252152 330200
rect 253296 330148 253348 330200
rect 254400 330148 254452 330200
rect 262588 330148 262640 330200
rect 316132 330148 316184 330200
rect 213828 330080 213880 330132
rect 252376 330080 252428 330132
rect 260564 330080 260616 330132
rect 310520 330080 310572 330132
rect 220728 330012 220780 330064
rect 252836 330012 252888 330064
rect 259828 330012 259880 330064
rect 303620 330012 303672 330064
rect 224868 329944 224920 329996
rect 259000 329944 259052 329996
rect 292672 329944 292724 329996
rect 227536 329876 227588 329928
rect 273352 329876 273404 329928
rect 273720 329876 273772 329928
rect 277676 329876 277728 329928
rect 278320 329876 278372 329928
rect 284300 329876 284352 329928
rect 284944 329876 284996 329928
rect 285496 329876 285548 329928
rect 288348 329876 288400 329928
rect 235264 329808 235316 329860
rect 267740 329808 267792 329860
rect 97908 329740 97960 329792
rect 242900 329740 242952 329792
rect 273904 329740 273956 329792
rect 95056 329672 95108 329724
rect 242624 329672 242676 329724
rect 276296 329740 276348 329792
rect 277308 329740 277360 329792
rect 279148 329740 279200 329792
rect 542360 329740 542412 329792
rect 277584 329672 277636 329724
rect 277952 329672 278004 329724
rect 279976 329672 280028 329724
rect 544384 329672 544436 329724
rect 91008 329604 91060 329656
rect 279700 329604 279752 329656
rect 279792 329604 279844 329656
rect 546500 329604 546552 329656
rect 86868 329536 86920 329588
rect 241888 329536 241940 329588
rect 284484 329536 284536 329588
rect 289636 329536 289688 329588
rect 553400 329536 553452 329588
rect 79968 329468 80020 329520
rect 241428 329468 241480 329520
rect 560300 329468 560352 329520
rect 77208 329400 77260 329452
rect 233240 329400 233292 329452
rect 280528 329400 280580 329452
rect 556252 329400 556304 329452
rect 50344 329332 50396 329384
rect 239036 329332 239088 329384
rect 281080 329332 281132 329384
rect 564532 329332 564584 329384
rect 46204 329264 46256 329316
rect 258172 329264 258224 329316
rect 258448 329264 258500 329316
rect 281264 329264 281316 329316
rect 566464 329264 566516 329316
rect 44824 329196 44876 329248
rect 237472 329196 237524 329248
rect 571340 329196 571392 329248
rect 22744 329128 22796 329180
rect 236000 329128 236052 329180
rect 282828 329128 282880 329180
rect 574100 329128 574152 329180
rect 14464 329060 14516 329112
rect 235908 329060 235960 329112
rect 281080 329060 281132 329112
rect 282460 329060 282512 329112
rect 576124 329060 576176 329112
rect 104808 328992 104860 329044
rect 243728 328992 243780 329044
rect 269212 328992 269264 329044
rect 416780 328992 416832 329044
rect 108948 328924 109000 328976
rect 261392 328924 261444 328976
rect 414020 328924 414072 328976
rect 111708 328856 111760 328908
rect 244096 328856 244148 328908
rect 322940 328856 322992 328908
rect 115848 328788 115900 328840
rect 244372 328788 244424 328840
rect 293960 328788 294012 328840
rect 119896 328720 119948 328772
rect 244740 328720 244792 328772
rect 280620 328720 280672 328772
rect 122748 328652 122800 328704
rect 161388 328584 161440 328636
rect 248052 328584 248104 328636
rect 86224 328380 86276 328432
rect 241796 328380 241848 328432
rect 80704 328312 80756 328364
rect 240876 328312 240928 328364
rect 266636 328312 266688 328364
rect 386420 328312 386472 328364
rect 75184 328244 75236 328296
rect 241060 328244 241112 328296
rect 267188 328244 267240 328296
rect 393320 328244 393372 328296
rect 70216 328176 70268 328228
rect 240600 328176 240652 328228
rect 267832 328176 267884 328228
rect 400220 328176 400272 328228
rect 68284 328108 68336 328160
rect 240324 328108 240376 328160
rect 283472 328108 283524 328160
rect 447048 328108 447100 328160
rect 62764 328040 62816 328092
rect 238944 328040 238996 328092
rect 283840 328040 283892 328092
rect 476028 328040 476080 328092
rect 57244 327972 57296 328024
rect 238852 327972 238904 328024
rect 282552 327972 282604 328024
rect 476580 327972 476632 328024
rect 51724 327904 51776 327956
rect 237196 327904 237248 327956
rect 283380 327904 283432 327956
rect 481732 327904 481784 327956
rect 53748 327836 53800 327888
rect 239312 327836 239364 327888
rect 283656 327836 283708 327888
rect 484860 327836 484912 327888
rect 11704 327768 11756 327820
rect 234896 327768 234948 327820
rect 283932 327768 283984 327820
rect 490564 327768 490616 327820
rect 10324 327700 10376 327752
rect 235632 327700 235684 327752
rect 283748 327700 283800 327752
rect 492680 327700 492732 327752
rect 93124 327632 93176 327684
rect 242440 327632 242492 327684
rect 99288 327564 99340 327616
rect 243820 327564 243872 327616
rect 195888 327496 195940 327548
rect 250904 327496 250956 327548
rect 231768 327428 231820 327480
rect 253756 327428 253808 327480
rect 215944 327360 215996 327412
rect 236460 327360 236512 327412
rect 125508 327020 125560 327072
rect 245108 327020 245160 327072
rect 124128 326952 124180 327004
rect 243452 326952 243504 327004
rect 115204 326884 115256 326936
rect 243268 326884 243320 326936
rect 106924 326816 106976 326868
rect 238668 326816 238720 326868
rect 107568 326748 107620 326800
rect 243636 326748 243688 326800
rect 106188 326680 106240 326732
rect 242164 326680 242216 326732
rect 83464 326612 83516 326664
rect 242716 326612 242768 326664
rect 63408 326544 63460 326596
rect 239128 326544 239180 326596
rect 58624 326476 58676 326528
rect 237748 326476 237800 326528
rect 255688 326476 255740 326528
rect 47584 326408 47636 326460
rect 237564 326408 237616 326460
rect 255412 326408 255464 326460
rect 255596 326408 255648 326460
rect 255964 326408 256016 326460
rect 257436 326408 257488 326460
rect 257620 326408 257672 326460
rect 257896 326408 257948 326460
rect 260012 326408 260064 326460
rect 260196 326408 260248 326460
rect 26884 326340 26936 326392
rect 234712 326340 234764 326392
rect 234988 326340 235040 326392
rect 235356 326340 235408 326392
rect 236736 326340 236788 326392
rect 237288 326340 237340 326392
rect 246028 326340 246080 326392
rect 246212 326340 246264 326392
rect 248788 326340 248840 326392
rect 249708 326340 249760 326392
rect 250168 326340 250220 326392
rect 251088 326340 251140 326392
rect 254584 326204 254636 326256
rect 255228 326204 255280 326256
rect 255872 326204 255924 326256
rect 256332 326340 256384 326392
rect 256516 326340 256568 326392
rect 262312 326340 262364 326392
rect 263140 326340 263192 326392
rect 267280 326476 267332 326528
rect 269488 326408 269540 326460
rect 269856 326408 269908 326460
rect 271420 326408 271472 326460
rect 271696 326408 271748 326460
rect 272708 326451 272760 326460
rect 272708 326417 272717 326451
rect 272717 326417 272751 326451
rect 272751 326417 272760 326451
rect 272708 326408 272760 326417
rect 329840 326408 329892 326460
rect 436928 326340 436980 326392
rect 257712 326204 257764 326256
rect 257804 326204 257856 326256
rect 257988 326204 258040 326256
rect 260012 326204 260064 326256
rect 260472 326204 260524 326256
rect 180156 325728 180208 325780
rect 236736 325728 236788 325780
rect 50436 325660 50488 325712
rect 235356 325660 235408 325712
rect 443644 325592 443696 325644
rect 580172 325592 580224 325644
rect 5448 324912 5500 324964
rect 235080 324912 235132 324964
rect 269672 324912 269724 324964
rect 270040 324912 270092 324964
rect 113088 323552 113140 323604
rect 240968 323552 241020 323604
rect 254492 323144 254544 323196
rect 254768 323144 254820 323196
rect 255504 322940 255556 322992
rect 255780 322940 255832 322992
rect 467104 322872 467156 322924
rect 471244 322872 471296 322924
rect 479524 322872 479576 322924
rect 480628 322872 480680 322924
rect 472256 322804 472308 322856
rect 474004 322804 474056 322856
rect 479156 322804 479208 322856
rect 232688 322736 232740 322788
rect 496820 322736 496872 322788
rect 232596 322668 232648 322720
rect 494244 322668 494296 322720
rect 464344 322600 464396 322652
rect 469404 322600 469456 322652
rect 472624 322600 472676 322652
rect 474556 322600 474608 322652
rect 506940 322600 506992 322652
rect 468484 322532 468536 322584
rect 504180 322532 504232 322584
rect 272708 322507 272760 322516
rect 272708 322473 272717 322507
rect 272717 322473 272751 322507
rect 272751 322473 272760 322507
rect 272708 322464 272760 322473
rect 284760 322464 284812 322516
rect 505468 322464 505520 322516
rect 285312 322396 285364 322448
rect 498660 322396 498712 322448
rect 285404 322328 285456 322380
rect 498200 322328 498252 322380
rect 287612 322260 287664 322312
rect 484400 322260 484452 322312
rect 233148 322192 233200 322244
rect 253020 322192 253072 322244
rect 447048 322192 447100 322244
rect 495532 322192 495584 322244
rect 519544 322192 519596 322244
rect 537116 322192 537168 322244
rect 465724 322124 465776 322176
rect 501052 322124 501104 322176
rect 447784 322056 447836 322108
rect 470692 322056 470744 322108
rect 476028 322056 476080 322108
rect 492220 322056 492272 322108
rect 449164 321988 449216 322040
rect 471980 321988 472032 322040
rect 233240 321920 233292 321972
rect 503260 321920 503312 321972
rect 232780 321852 232832 321904
rect 500684 321852 500736 321904
rect 232228 321784 232280 321836
rect 475476 321784 475528 321836
rect 232412 321716 232464 321768
rect 478236 321716 478288 321768
rect 481732 321580 481784 321632
rect 488172 321580 488224 321632
rect 530032 321580 530084 321632
rect 530676 321580 530728 321632
rect 537208 321580 537260 321632
rect 286784 320832 286836 320884
rect 581000 320832 581052 320884
rect 251640 320152 251692 320204
rect 252008 320152 252060 320204
rect 3516 320084 3568 320136
rect 14648 320084 14700 320136
rect 547236 313216 547288 313268
rect 580172 313216 580224 313268
rect 3516 306280 3568 306332
rect 35256 306280 35308 306332
rect 537484 299412 537536 299464
rect 580172 299412 580224 299464
rect 3056 293904 3108 293956
rect 33876 293904 33928 293956
rect 246304 274592 246356 274644
rect 437480 274592 437532 274644
rect 540428 273164 540480 273216
rect 579988 273164 580040 273216
rect 245200 272484 245252 272536
rect 436652 272484 436704 272536
rect 248604 271804 248656 271856
rect 436836 271804 436888 271856
rect 250720 270444 250772 270496
rect 436836 270444 436888 270496
rect 268568 269764 268620 269816
rect 357532 269764 357584 269816
rect 436928 269016 436980 269068
rect 437296 269016 437348 269068
rect 3516 267656 3568 267708
rect 17316 267656 17368 267708
rect 245108 266976 245160 267028
rect 436100 266976 436152 267028
rect 544476 259360 544528 259412
rect 580172 259360 580224 259412
rect 3148 255212 3200 255264
rect 36636 255212 36688 255264
rect 232044 248344 232096 248396
rect 436100 248344 436152 248396
rect 3516 241408 3568 241460
rect 18696 241408 18748 241460
rect 282644 240728 282696 240780
rect 439136 240728 439188 240780
rect 297732 239980 297784 240032
rect 439872 239980 439924 240032
rect 445668 239912 445720 239964
rect 538496 239912 538548 239964
rect 438676 239844 438728 239896
rect 445760 239844 445812 239896
rect 522672 239844 522724 239896
rect 438768 239776 438820 239828
rect 523132 239776 523184 239828
rect 438584 239708 438636 239760
rect 523040 239708 523092 239760
rect 284852 239640 284904 239692
rect 436008 239640 436060 239692
rect 445760 239640 445812 239692
rect 445852 239640 445904 239692
rect 451096 239640 451148 239692
rect 451188 239640 451240 239692
rect 456064 239640 456116 239692
rect 537208 239640 537260 239692
rect 437388 239572 437440 239624
rect 505008 239572 505060 239624
rect 299020 239504 299072 239556
rect 298928 239436 298980 239488
rect 452568 239436 452620 239488
rect 452752 239504 452804 239556
rect 456064 239504 456116 239556
rect 460940 239504 460992 239556
rect 461032 239504 461084 239556
rect 473176 239504 473228 239556
rect 288164 239368 288216 239420
rect 479340 239436 479392 239488
rect 471980 239368 472032 239420
rect 288072 239300 288124 239352
rect 475660 239300 475712 239352
rect 297548 239232 297600 239284
rect 487896 239232 487948 239284
rect 297456 239164 297508 239216
rect 501880 239164 501932 239216
rect 297364 239096 297416 239148
rect 503076 239096 503128 239148
rect 298744 239028 298796 239080
rect 505560 239028 505612 239080
rect 292212 238960 292264 239012
rect 506756 238960 506808 239012
rect 232964 238892 233016 238944
rect 495624 238892 495676 238944
rect 233056 238824 233108 238876
rect 496820 238824 496872 238876
rect 234436 238756 234488 238808
rect 500500 238756 500552 238808
rect 296260 238688 296312 238740
rect 485412 238688 485464 238740
rect 291844 238620 291896 238672
rect 477684 238620 477736 238672
rect 296076 238552 296128 238604
rect 484400 238552 484452 238604
rect 292028 238484 292080 238536
rect 483388 238484 483440 238536
rect 290556 238416 290608 238468
rect 482284 238416 482336 238468
rect 292304 238348 292356 238400
rect 484860 238348 484912 238400
rect 293592 238280 293644 238332
rect 488172 238280 488224 238332
rect 292120 238212 292172 238264
rect 485964 238212 486016 238264
rect 293500 238144 293552 238196
rect 491668 238144 491720 238196
rect 259092 238076 259144 238128
rect 284392 238076 284444 238128
rect 294788 238076 294840 238128
rect 495164 238076 495216 238128
rect 258816 238008 258868 238060
rect 287060 238008 287112 238060
rect 293408 238008 293460 238060
rect 492772 238008 492824 238060
rect 296352 237940 296404 237992
rect 481732 237940 481784 237992
rect 291936 237872 291988 237924
rect 476580 237872 476632 237924
rect 296444 237804 296496 237856
rect 480628 237804 480680 237856
rect 294880 237736 294932 237788
rect 467196 237736 467248 237788
rect 296536 237668 296588 237720
rect 467840 237668 467892 237720
rect 294696 237600 294748 237652
rect 465080 237600 465132 237652
rect 292396 237532 292448 237584
rect 462320 237532 462372 237584
rect 295064 237464 295116 237516
rect 463700 237464 463752 237516
rect 438308 237396 438360 237448
rect 485780 237396 485832 237448
rect 233792 237328 233844 237380
rect 470600 237328 470652 237380
rect 505008 237328 505060 237380
rect 521660 237328 521712 237380
rect 233700 237260 233752 237312
rect 467840 237260 467892 237312
rect 288348 237192 288400 237244
rect 503720 237192 503772 237244
rect 289636 237124 289688 237176
rect 498200 237124 498252 237176
rect 285220 237056 285272 237108
rect 492680 237056 492732 237108
rect 288256 236988 288308 237040
rect 494060 236988 494112 237040
rect 286692 236920 286744 236972
rect 491300 236920 491352 236972
rect 286600 236852 286652 236904
rect 490288 236852 490340 236904
rect 282092 236784 282144 236836
rect 473360 236784 473412 236836
rect 258448 236716 258500 236768
rect 282920 236716 282972 236768
rect 296168 236716 296220 236768
rect 485780 236716 485832 236768
rect 281816 236648 281868 236700
rect 469220 236648 469272 236700
rect 289452 236580 289504 236632
rect 471980 236580 472032 236632
rect 298836 236512 298888 236564
rect 476120 236512 476172 236564
rect 289544 236444 289596 236496
rect 461124 236444 461176 236496
rect 294972 236376 295024 236428
rect 465080 236376 465132 236428
rect 344560 236308 344612 236360
rect 488540 236308 488592 236360
rect 344468 236240 344520 236292
rect 474740 236240 474792 236292
rect 344376 236172 344428 236224
rect 470876 236172 470928 236224
rect 440240 236104 440292 236156
rect 495440 236104 495492 236156
rect 439136 236036 439188 236088
rect 469220 236036 469272 236088
rect 275376 235900 275428 235952
rect 488540 235900 488592 235952
rect 274824 235832 274876 235884
rect 490564 235832 490616 235884
rect 275560 235764 275612 235816
rect 493324 235764 493376 235816
rect 276664 235696 276716 235748
rect 497464 235696 497516 235748
rect 276572 235628 276624 235680
rect 500224 235628 500276 235680
rect 276480 235560 276532 235612
rect 501604 235560 501656 235612
rect 276756 235492 276808 235544
rect 502340 235492 502392 235544
rect 276848 235424 276900 235476
rect 506480 235424 506532 235476
rect 277400 235356 277452 235408
rect 508504 235356 508556 235408
rect 278136 235288 278188 235340
rect 512644 235288 512696 235340
rect 277952 235220 278004 235272
rect 520280 235220 520332 235272
rect 273996 235152 274048 235204
rect 484400 235152 484452 235204
rect 275468 235084 275520 235136
rect 483664 235084 483716 235136
rect 274088 235016 274140 235068
rect 481732 235016 481784 235068
rect 274180 234948 274232 235000
rect 475384 234948 475436 235000
rect 273260 234880 273312 234932
rect 472624 234880 472676 234932
rect 272800 234812 272852 234864
rect 459560 234812 459612 234864
rect 272892 234744 272944 234796
rect 456892 234744 456944 234796
rect 271236 234676 271288 234728
rect 441620 234676 441672 234728
rect 418896 234608 418948 234660
rect 477500 234608 477552 234660
rect 272984 234540 273036 234592
rect 466460 234540 466512 234592
rect 274364 234472 274416 234524
rect 470600 234472 470652 234524
rect 274272 234404 274324 234456
rect 472716 234404 472768 234456
rect 273628 234336 273680 234388
rect 476764 234336 476816 234388
rect 273352 234268 273404 234320
rect 479524 234268 479576 234320
rect 275744 234200 275796 234252
rect 490012 234200 490064 234252
rect 275008 234132 275060 234184
rect 492680 234132 492732 234184
rect 275652 234064 275704 234116
rect 496820 234064 496872 234116
rect 276940 233996 276992 234048
rect 503720 233996 503772 234048
rect 277032 233928 277084 233980
rect 506572 233928 506624 233980
rect 278228 233860 278280 233912
rect 519544 233860 519596 233912
rect 271880 233792 271932 233844
rect 463700 233792 463752 233844
rect 271420 233724 271472 233776
rect 448612 233724 448664 233776
rect 271328 233656 271380 233708
rect 445760 233656 445812 233708
rect 270868 232908 270920 232960
rect 440332 232908 440384 232960
rect 271512 232840 271564 232892
rect 443000 232840 443052 232892
rect 272064 232772 272116 232824
rect 465172 232772 465224 232824
rect 277124 232704 277176 232756
rect 510620 232704 510672 232756
rect 278320 232636 278372 232688
rect 521660 232636 521712 232688
rect 278504 232568 278556 232620
rect 524420 232568 524472 232620
rect 260104 232500 260156 232552
rect 276020 232500 276072 232552
rect 278412 232500 278464 232552
rect 528560 232500 528612 232552
rect 274916 231140 274968 231192
rect 499580 231140 499632 231192
rect 276112 231072 276164 231124
rect 514760 231072 514812 231124
rect 286508 219376 286560 219428
rect 580172 219376 580224 219428
rect 3332 215228 3384 215280
rect 32496 215228 32548 215280
rect 3056 202784 3108 202836
rect 39396 202784 39448 202836
rect 3516 188980 3568 189032
rect 21456 188980 21508 189032
rect 543096 179324 543148 179376
rect 579620 179324 579672 179376
rect 271052 177352 271104 177404
rect 447140 177352 447192 177404
rect 276296 177284 276348 177336
rect 517520 177284 517572 177336
rect 277676 175924 277728 175976
rect 530584 175924 530636 175976
rect 3240 164160 3292 164212
rect 14556 164160 14608 164212
rect 3516 150356 3568 150408
rect 40776 150356 40828 150408
rect 573364 139340 573416 139392
rect 580172 139340 580224 139392
rect 3516 137912 3568 137964
rect 29644 137912 29696 137964
rect 3148 111732 3200 111784
rect 11796 111732 11848 111784
rect 569316 100648 569368 100700
rect 580172 100648 580224 100700
rect 3516 97928 3568 97980
rect 33784 97928 33836 97980
rect 264520 93100 264572 93152
rect 273260 93100 273312 93152
rect 313924 86912 313976 86964
rect 580172 86912 580224 86964
rect 3516 85484 3568 85536
rect 17224 85484 17276 85536
rect 302884 73108 302936 73160
rect 580172 73108 580224 73160
rect 2780 71612 2832 71664
rect 4804 71612 4856 71664
rect 555424 60664 555476 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 35164 59304 35216 59356
rect 295984 46860 296036 46912
rect 580172 46860 580224 46912
rect 3516 45500 3568 45552
rect 18604 45500 18656 45552
rect 300124 33056 300176 33108
rect 580172 33056 580224 33108
rect 3424 20612 3476 20664
rect 152464 20612 152516 20664
rect 540244 20612 540296 20664
rect 579988 20612 580040 20664
rect 265716 18572 265768 18624
rect 372620 18572 372672 18624
rect 51816 13064 51868 13116
rect 238576 13064 238628 13116
rect 357532 11704 357584 11756
rect 358728 11704 358780 11756
rect 374092 11704 374144 11756
rect 375288 11704 375340 11756
rect 398932 11704 398984 11756
rect 400128 11704 400180 11756
rect 448612 11704 448664 11756
rect 449808 11704 449860 11756
rect 260472 10956 260524 11008
rect 314660 10956 314712 11008
rect 261576 10888 261628 10940
rect 317972 10888 318024 10940
rect 261760 10820 261812 10872
rect 322112 10820 322164 10872
rect 261668 10752 261720 10804
rect 324320 10752 324372 10804
rect 261852 10684 261904 10736
rect 328736 10684 328788 10736
rect 261484 10616 261536 10668
rect 332692 10616 332744 10668
rect 262772 10548 262824 10600
rect 336280 10548 336332 10600
rect 262680 10480 262732 10532
rect 339500 10480 339552 10532
rect 263048 10412 263100 10464
rect 342904 10412 342956 10464
rect 262956 10344 263008 10396
rect 346952 10344 347004 10396
rect 245108 10276 245160 10328
rect 254492 10276 254544 10328
rect 262864 10276 262916 10328
rect 349160 10276 349212 10328
rect 252652 9528 252704 9580
rect 254308 9528 254360 9580
rect 253480 8440 253532 8492
rect 255596 8440 255648 8492
rect 3424 6808 3476 6860
rect 21364 6808 21416 6860
rect 318064 6808 318116 6860
rect 580172 6808 580224 6860
rect 259552 6672 259604 6724
rect 313832 6672 313884 6724
rect 262036 6604 262088 6656
rect 324412 6604 324464 6656
rect 261944 6536 261996 6588
rect 328000 6536 328052 6588
rect 262128 6468 262180 6520
rect 331588 6468 331640 6520
rect 263140 6400 263192 6452
rect 335084 6400 335136 6452
rect 263232 6332 263284 6384
rect 338672 6332 338724 6384
rect 263324 6264 263376 6316
rect 342168 6264 342220 6316
rect 262404 6196 262456 6248
rect 345756 6196 345808 6248
rect 75000 6128 75052 6180
rect 240692 6128 240744 6180
rect 262220 6128 262272 6180
rect 349252 6128 349304 6180
rect 257068 5448 257120 5500
rect 278320 5448 278372 5500
rect 286416 5448 286468 5500
rect 411904 5448 411956 5500
rect 269304 5380 269356 5432
rect 424968 5380 425020 5432
rect 256332 5312 256384 5364
rect 264152 5312 264204 5364
rect 269672 5312 269724 5364
rect 429660 5312 429712 5364
rect 257804 5244 257856 5296
rect 268844 5244 268896 5296
rect 270224 5244 270276 5296
rect 432052 5244 432104 5296
rect 257436 5176 257488 5228
rect 284944 5176 284996 5228
rect 454500 5176 454552 5228
rect 234620 5108 234672 5160
rect 249064 5108 249116 5160
rect 257620 5108 257672 5160
rect 270592 5108 270644 5160
rect 270684 5108 270736 5160
rect 450912 5108 450964 5160
rect 209780 5040 209832 5092
rect 251640 5040 251692 5092
rect 257252 5040 257304 5092
rect 281908 5040 281960 5092
rect 286324 5040 286376 5092
rect 468668 5040 468720 5092
rect 181444 4972 181496 5024
rect 248788 4972 248840 5024
rect 257712 4972 257764 5024
rect 272432 4972 272484 5024
rect 273904 4972 273956 5024
rect 455696 4972 455748 5024
rect 145932 4904 145984 4956
rect 246672 4904 246724 4956
rect 257896 4904 257948 4956
rect 279516 4904 279568 4956
rect 279608 4904 279660 4956
rect 486424 4904 486476 4956
rect 135260 4836 135312 4888
rect 246212 4836 246264 4888
rect 257344 4836 257396 4888
rect 267740 4836 267792 4888
rect 276020 4836 276072 4888
rect 301964 4836 302016 4888
rect 304264 4836 304316 4888
rect 582196 4836 582248 4888
rect 67916 4768 67968 4820
rect 240600 4768 240652 4820
rect 258632 4768 258684 4820
rect 297272 4768 297324 4820
rect 299572 4768 299624 4820
rect 300768 4768 300820 4820
rect 304448 4768 304500 4820
rect 265808 4700 265860 4752
rect 379980 4700 380032 4752
rect 268384 4632 268436 4684
rect 269856 4564 269908 4616
rect 351644 4564 351696 4616
rect 365812 4564 365864 4616
rect 264244 4496 264296 4548
rect 260012 4428 260064 4480
rect 312636 4428 312688 4480
rect 326804 4428 326856 4480
rect 257528 4360 257580 4412
rect 274824 4360 274876 4412
rect 285036 4360 285088 4412
rect 333888 4360 333940 4412
rect 259920 4292 259972 4344
rect 307944 4292 307996 4344
rect 269948 4224 270000 4276
rect 309048 4224 309100 4276
rect 268476 4156 268528 4208
rect 13544 4088 13596 4140
rect 22744 4088 22796 4140
rect 27712 4088 27764 4140
rect 51724 4088 51776 4140
rect 99840 4088 99892 4140
rect 247592 4088 247644 4140
rect 251180 4088 251232 4140
rect 270592 4156 270644 4208
rect 271236 4156 271288 4208
rect 285128 4156 285180 4208
rect 319720 4156 319772 4208
rect 324320 4156 324372 4208
rect 325608 4156 325660 4208
rect 279700 4088 279752 4140
rect 475752 4088 475804 4140
rect 483664 4088 483716 4140
rect 492312 4088 492364 4140
rect 547144 4088 547196 4140
rect 549076 4088 549128 4140
rect 566464 4088 566516 4140
rect 568028 4088 568080 4140
rect 572 4020 624 4072
rect 32312 4020 32364 4072
rect 34796 4020 34848 4072
rect 58624 4020 58676 4072
rect 92756 4020 92808 4072
rect 242072 4020 242124 4072
rect 257068 4020 257120 4072
rect 259460 4020 259512 4072
rect 280804 4020 280856 4072
rect 544384 4020 544436 4072
rect 550272 4020 550324 4072
rect 1676 3952 1728 4004
rect 36544 3952 36596 4004
rect 44272 3952 44324 4004
rect 46204 3952 46256 4004
rect 85672 3952 85724 4004
rect 241980 3952 242032 4004
rect 245200 3952 245252 4004
rect 251916 3952 251968 4004
rect 287980 3952 288032 4004
rect 491116 3952 491168 4004
rect 20628 3884 20680 3936
rect 173164 3884 173216 3936
rect 173716 3884 173768 3936
rect 174268 3884 174320 3936
rect 175188 3884 175240 3936
rect 175464 3884 175516 3936
rect 176568 3884 176620 3936
rect 176660 3884 176712 3936
rect 177948 3884 178000 3936
rect 180248 3884 180300 3936
rect 180708 3884 180760 3936
rect 182548 3884 182600 3936
rect 183468 3884 183520 3936
rect 183744 3884 183796 3936
rect 184848 3884 184900 3936
rect 184940 3884 184992 3936
rect 186044 3884 186096 3936
rect 188528 3884 188580 3936
rect 188988 3884 189040 3936
rect 189724 3884 189776 3936
rect 190368 3884 190420 3936
rect 190828 3884 190880 3936
rect 191748 3884 191800 3936
rect 192024 3884 192076 3936
rect 193128 3884 193180 3936
rect 193220 3884 193272 3936
rect 194508 3884 194560 3936
rect 196808 3884 196860 3936
rect 197268 3884 197320 3936
rect 199108 3884 199160 3936
rect 200028 3884 200080 3936
rect 200304 3884 200356 3936
rect 201408 3884 201460 3936
rect 201500 3884 201552 3936
rect 202788 3884 202840 3936
rect 205088 3884 205140 3936
rect 205548 3884 205600 3936
rect 206192 3884 206244 3936
rect 206928 3884 206980 3936
rect 207388 3884 207440 3936
rect 208308 3884 208360 3936
rect 250168 3884 250220 3936
rect 280988 3884 281040 3936
rect 484032 3884 484084 3936
rect 497464 3884 497516 3936
rect 510068 3884 510120 3936
rect 2872 3816 2924 3868
rect 39304 3816 39356 3868
rect 7656 3748 7708 3800
rect 43444 3816 43496 3868
rect 43076 3748 43128 3800
rect 51816 3816 51868 3868
rect 69112 3816 69164 3868
rect 70216 3816 70268 3868
rect 71504 3816 71556 3868
rect 235816 3816 235868 3868
rect 245016 3816 245068 3868
rect 246396 3816 246448 3868
rect 252652 3816 252704 3868
rect 280896 3816 280948 3868
rect 487620 3816 487672 3868
rect 500316 3816 500368 3868
rect 11152 3680 11204 3732
rect 50436 3748 50488 3800
rect 60832 3748 60884 3800
rect 50160 3680 50212 3732
rect 50988 3680 51040 3732
rect 51356 3680 51408 3732
rect 53104 3680 53156 3732
rect 53656 3680 53708 3732
rect 239404 3748 239456 3800
rect 241704 3748 241756 3800
rect 250444 3748 250496 3800
rect 287704 3748 287756 3800
rect 494704 3748 494756 3800
rect 9956 3612 10008 3664
rect 26884 3612 26936 3664
rect 28908 3612 28960 3664
rect 213368 3612 213420 3664
rect 213828 3612 213880 3664
rect 214472 3612 214524 3664
rect 215208 3612 215260 3664
rect 215668 3612 215720 3664
rect 216588 3612 216640 3664
rect 216864 3612 216916 3664
rect 217968 3612 218020 3664
rect 218060 3612 218112 3664
rect 219348 3612 219400 3664
rect 221556 3612 221608 3664
rect 222108 3612 222160 3664
rect 222752 3612 222804 3664
rect 223488 3612 223540 3664
rect 223948 3612 224000 3664
rect 224868 3612 224920 3664
rect 225144 3612 225196 3664
rect 226248 3612 226300 3664
rect 226340 3612 226392 3664
rect 227628 3612 227680 3664
rect 231216 3612 231268 3664
rect 238024 3680 238076 3732
rect 244096 3680 244148 3732
rect 253204 3680 253256 3732
rect 287888 3680 287940 3732
rect 498200 3680 498252 3732
rect 501604 3680 501656 3732
rect 576124 3748 576176 3800
rect 578608 3748 578660 3800
rect 238116 3612 238168 3664
rect 240508 3612 240560 3664
rect 249984 3612 250036 3664
rect 287796 3612 287848 3664
rect 501788 3612 501840 3664
rect 513564 3680 513616 3732
rect 517152 3612 517204 3664
rect 551284 3612 551336 3664
rect 559748 3612 559800 3664
rect 23020 3544 23072 3596
rect 231124 3544 231176 3596
rect 239312 3544 239364 3596
rect 250536 3544 250588 3596
rect 256424 3544 256476 3596
rect 260656 3544 260708 3596
rect 284300 3544 284352 3596
rect 285404 3544 285456 3596
rect 289360 3544 289412 3596
rect 505376 3544 505428 3596
rect 508504 3544 508556 3596
rect 524236 3544 524288 3596
rect 534908 3544 534960 3596
rect 536932 3544 536984 3596
rect 564440 3544 564492 3596
rect 565636 3544 565688 3596
rect 574836 3544 574888 3596
rect 577412 3544 577464 3596
rect 8760 3476 8812 3528
rect 10324 3476 10376 3528
rect 24216 3476 24268 3528
rect 24768 3476 24820 3528
rect 4068 3408 4120 3460
rect 11704 3408 11756 3460
rect 21824 3408 21876 3460
rect 32404 3408 32456 3460
rect 33048 3408 33100 3460
rect 229836 3476 229888 3528
rect 230388 3476 230440 3528
rect 231032 3476 231084 3528
rect 231768 3476 231820 3528
rect 232228 3476 232280 3528
rect 233148 3476 233200 3528
rect 233424 3476 233476 3528
rect 234528 3476 234580 3528
rect 237012 3476 237064 3528
rect 249156 3476 249208 3528
rect 249984 3476 250036 3528
rect 254584 3476 254636 3528
rect 254676 3476 254728 3528
rect 255504 3476 255556 3528
rect 256516 3476 256568 3528
rect 258264 3476 258316 3528
rect 258724 3476 258776 3528
rect 259460 3476 259512 3528
rect 264704 3476 264756 3528
rect 265348 3476 265400 3528
rect 289084 3476 289136 3528
rect 508872 3476 508924 3528
rect 519636 3476 519688 3528
rect 19432 3340 19484 3392
rect 26516 3272 26568 3324
rect 40592 3340 40644 3392
rect 48964 3340 49016 3392
rect 50344 3340 50396 3392
rect 52552 3340 52604 3392
rect 53748 3340 53800 3392
rect 56048 3340 56100 3392
rect 57152 3340 57204 3392
rect 57244 3340 57296 3392
rect 57888 3340 57940 3392
rect 59636 3340 59688 3392
rect 62764 3340 62816 3392
rect 64328 3340 64380 3392
rect 64788 3340 64840 3392
rect 66720 3340 66772 3392
rect 68284 3340 68336 3392
rect 72608 3340 72660 3392
rect 73068 3340 73120 3392
rect 76196 3340 76248 3392
rect 77208 3340 77260 3392
rect 80888 3340 80940 3392
rect 81348 3340 81400 3392
rect 83280 3340 83332 3392
rect 84108 3340 84160 3392
rect 84476 3340 84528 3392
rect 86224 3340 86276 3392
rect 89168 3340 89220 3392
rect 89628 3340 89680 3392
rect 90364 3340 90416 3392
rect 91008 3340 91060 3392
rect 91560 3340 91612 3392
rect 93124 3340 93176 3392
rect 93952 3340 94004 3392
rect 95056 3340 95108 3392
rect 97448 3340 97500 3392
rect 97908 3340 97960 3392
rect 98644 3340 98696 3392
rect 99288 3340 99340 3392
rect 101036 3340 101088 3392
rect 102048 3340 102100 3392
rect 102232 3340 102284 3392
rect 231308 3408 231360 3460
rect 238116 3408 238168 3460
rect 235264 3340 235316 3392
rect 242900 3408 242952 3460
rect 245108 3408 245160 3460
rect 248788 3408 248840 3460
rect 253388 3408 253440 3460
rect 255872 3408 255924 3460
rect 261760 3408 261812 3460
rect 289268 3408 289320 3460
rect 512460 3408 512512 3460
rect 512644 3408 512696 3460
rect 527824 3408 527876 3460
rect 530584 3476 530636 3528
rect 532516 3476 532568 3528
rect 536104 3476 536156 3528
rect 537024 3476 537076 3528
rect 540336 3476 540388 3528
rect 541992 3476 542044 3528
rect 548524 3476 548576 3528
rect 552664 3476 552716 3528
rect 562324 3476 562376 3528
rect 566832 3476 566884 3528
rect 531320 3408 531372 3460
rect 538956 3408 539008 3460
rect 539600 3408 539652 3460
rect 253296 3340 253348 3392
rect 283564 3340 283616 3392
rect 468484 3340 468536 3392
rect 469864 3340 469916 3392
rect 472624 3340 472676 3392
rect 473452 3340 473504 3392
rect 476764 3340 476816 3392
rect 478144 3340 478196 3392
rect 480536 3340 480588 3392
rect 41880 3272 41932 3324
rect 106832 3272 106884 3324
rect 106924 3272 106976 3324
rect 107568 3272 107620 3324
rect 108120 3272 108172 3324
rect 108948 3272 109000 3324
rect 109316 3272 109368 3324
rect 110328 3272 110380 3324
rect 115204 3272 115256 3324
rect 115848 3272 115900 3324
rect 116400 3272 116452 3324
rect 117228 3272 117280 3324
rect 118792 3272 118844 3324
rect 119804 3272 119856 3324
rect 122288 3272 122340 3324
rect 122748 3272 122800 3324
rect 123484 3272 123536 3324
rect 124128 3272 124180 3324
rect 124680 3272 124732 3324
rect 125508 3272 125560 3324
rect 126980 3272 127032 3324
rect 128268 3272 128320 3324
rect 130568 3272 130620 3324
rect 131028 3272 131080 3324
rect 131764 3272 131816 3324
rect 132408 3272 132460 3324
rect 134156 3272 134208 3324
rect 135168 3272 135220 3324
rect 138848 3272 138900 3324
rect 139308 3272 139360 3324
rect 140044 3272 140096 3324
rect 140688 3272 140740 3324
rect 35992 3204 36044 3256
rect 47584 3204 47636 3256
rect 82084 3204 82136 3256
rect 83464 3204 83516 3256
rect 105728 3204 105780 3256
rect 106188 3204 106240 3256
rect 125876 3204 125928 3256
rect 244648 3272 244700 3324
rect 251180 3272 251232 3324
rect 255688 3272 255740 3324
rect 258356 3272 258408 3324
rect 262956 3272 263008 3324
rect 282184 3272 282236 3324
rect 292580 3272 292632 3324
rect 294604 3272 294656 3324
rect 18236 3136 18288 3188
rect 25504 3136 25556 3188
rect 65524 3136 65576 3188
rect 66168 3136 66220 3188
rect 114008 3136 114060 3188
rect 115112 3136 115164 3188
rect 132960 3136 133012 3188
rect 244924 3204 244976 3256
rect 264428 3204 264480 3256
rect 270040 3204 270092 3256
rect 281080 3204 281132 3256
rect 461584 3204 461636 3256
rect 472256 3204 472308 3256
rect 475384 3272 475436 3324
rect 476948 3272 477000 3324
rect 479524 3272 479576 3324
rect 482836 3272 482888 3324
rect 493324 3272 493376 3324
rect 499396 3272 499448 3324
rect 569224 3272 569276 3324
rect 570328 3272 570380 3324
rect 479340 3204 479392 3256
rect 141240 3136 141292 3188
rect 142068 3136 142120 3188
rect 142436 3136 142488 3188
rect 143448 3136 143500 3188
rect 147128 3136 147180 3188
rect 147588 3136 147640 3188
rect 148324 3136 148376 3188
rect 148968 3136 149020 3188
rect 149520 3136 149572 3188
rect 150348 3136 150400 3188
rect 40684 3068 40736 3120
rect 44824 3068 44876 3120
rect 143540 3068 143592 3120
rect 246120 3136 246172 3188
rect 279792 3136 279844 3188
rect 458088 3136 458140 3188
rect 538864 3136 538916 3188
rect 540796 3136 540848 3188
rect 543004 3136 543056 3188
rect 545488 3136 545540 3188
rect 150624 3068 150676 3120
rect 151728 3068 151780 3120
rect 151820 3068 151872 3120
rect 153108 3068 153160 3120
rect 155408 3068 155460 3120
rect 155868 3068 155920 3120
rect 156604 3068 156656 3120
rect 157248 3068 157300 3120
rect 157800 3068 157852 3120
rect 158628 3068 158680 3120
rect 158904 3068 158956 3120
rect 160008 3068 160060 3120
rect 160100 3068 160152 3120
rect 161388 3068 161440 3120
rect 163688 3068 163740 3120
rect 164148 3068 164200 3120
rect 164884 3068 164936 3120
rect 165528 3068 165580 3120
rect 166080 3068 166132 3120
rect 166908 3068 166960 3120
rect 167184 3068 167236 3120
rect 168288 3068 168340 3120
rect 168380 3068 168432 3120
rect 169668 3068 169720 3120
rect 232504 3068 232556 3120
rect 278044 3068 278096 3120
rect 445024 3068 445076 3120
rect 472716 3068 472768 3120
rect 474556 3068 474608 3120
rect 12348 3000 12400 3052
rect 14464 3000 14516 3052
rect 58440 3000 58492 3052
rect 61384 3000 61436 3052
rect 117596 3000 117648 3052
rect 37188 2932 37240 2984
rect 43536 2932 43588 2984
rect 73804 2932 73856 2984
rect 75184 2932 75236 2984
rect 77392 2932 77444 2984
rect 80704 2932 80756 2984
rect 110512 2932 110564 2984
rect 161572 2932 161624 2984
rect 180156 3000 180208 3052
rect 197912 3000 197964 3052
rect 208584 3000 208636 3052
rect 251548 3000 251600 3052
rect 282276 3000 282328 3052
rect 427268 3000 427320 3052
rect 429844 3000 429896 3052
rect 434444 3000 434496 3052
rect 439596 3000 439648 3052
rect 441528 3000 441580 3052
rect 178684 2932 178736 2984
rect 215944 2932 215996 2984
rect 236644 2932 236696 2984
rect 267004 2932 267056 2984
rect 337476 2932 337528 2984
rect 337568 2932 337620 2984
rect 171784 2864 171836 2916
rect 171968 2864 172020 2916
rect 231400 2864 231452 2916
rect 258908 2864 258960 2916
rect 296076 2864 296128 2916
rect 300216 2864 300268 2916
rect 340972 2864 341024 2916
rect 341524 2932 341576 2984
rect 344284 2864 344336 2916
rect 348056 2932 348108 2984
rect 348424 2932 348476 2984
rect 365720 2932 365772 2984
rect 367008 2932 367060 2984
rect 369400 2932 369452 2984
rect 369492 2932 369544 2984
rect 390652 2932 390704 2984
rect 391204 2932 391256 2984
rect 121092 2796 121144 2848
rect 180064 2796 180116 2848
rect 269764 2796 269816 2848
rect 305552 2796 305604 2848
rect 316040 2796 316092 2848
rect 317328 2796 317380 2848
rect 316684 2728 316736 2780
rect 344560 2796 344612 2848
rect 355232 2864 355284 2916
rect 355324 2864 355376 2916
rect 376484 2864 376536 2916
rect 376576 2864 376628 2916
rect 397736 2864 397788 2916
rect 404820 2932 404872 2984
rect 405004 2932 405056 2984
rect 405464 2932 405516 2984
rect 415492 2932 415544 2984
rect 416044 2932 416096 2984
rect 418804 2932 418856 2984
rect 420184 2932 420236 2984
rect 426164 2932 426216 2984
rect 432604 2932 432656 2984
rect 437940 2932 437992 2984
rect 438216 2932 438268 2984
rect 459192 3000 459244 3052
rect 408408 2864 408460 2916
rect 362316 2796 362368 2848
rect 362408 2796 362460 2848
rect 398288 2796 398340 2848
rect 405648 2796 405700 2848
rect 407764 2796 407816 2848
rect 422576 2864 422628 2916
rect 422944 2864 422996 2916
rect 436744 2864 436796 2916
rect 439504 2864 439556 2916
rect 448612 2864 448664 2916
rect 490564 2864 490616 2916
rect 495900 2864 495952 2916
rect 558276 2864 558328 2916
rect 563244 2864 563296 2916
rect 418988 2796 419040 2848
rect 382924 2660 382976 2712
rect 420276 2796 420328 2848
rect 433248 2796 433300 2848
rect 438124 2796 438176 2848
rect 452108 2796 452160 2848
rect 583392 2839 583444 2848
rect 583392 2805 583401 2839
rect 583401 2805 583435 2839
rect 583435 2805 583444 2839
rect 583392 2796 583444 2805
rect 383568 2592 383620 2644
rect 349160 1504 349212 1556
rect 350448 1504 350500 1556
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700398 8156 703520
rect 24320 700534 24348 703520
rect 40512 700670 40540 703520
rect 72988 700806 73016 703520
rect 89180 700874 89208 703520
rect 89168 700868 89220 700874
rect 89168 700810 89220 700816
rect 72976 700800 73028 700806
rect 72976 700742 73028 700748
rect 40500 700664 40552 700670
rect 40500 700606 40552 700612
rect 24308 700528 24360 700534
rect 24308 700470 24360 700476
rect 8116 700392 8168 700398
rect 8116 700334 8168 700340
rect 105464 700330 105492 703520
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 137848 700262 137876 703520
rect 137836 700256 137888 700262
rect 137836 700198 137888 700204
rect 154132 700194 154160 703520
rect 170324 700466 170352 703520
rect 170312 700460 170364 700466
rect 170312 700402 170364 700408
rect 154120 700188 154172 700194
rect 154120 700130 154172 700136
rect 202800 699990 202828 703520
rect 202788 699984 202840 699990
rect 202788 699926 202840 699932
rect 218992 699922 219020 703520
rect 218980 699916 219032 699922
rect 218980 699858 219032 699864
rect 235184 699718 235212 703520
rect 254952 701004 255004 701010
rect 254952 700946 255004 700952
rect 253664 700732 253716 700738
rect 253664 700674 253716 700680
rect 240784 700460 240836 700466
rect 240784 700402 240836 700408
rect 252192 700460 252244 700466
rect 252192 700402 252244 700408
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 238024 699712 238076 699718
rect 238024 699654 238076 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 670818 3464 671191
rect 3424 670812 3476 670818
rect 3424 670754 3476 670760
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 238036 391406 238064 699654
rect 240796 391474 240824 700402
rect 242164 700324 242216 700330
rect 242164 700266 242216 700272
rect 242176 391814 242204 700266
rect 251088 670744 251140 670750
rect 251088 670686 251140 670692
rect 250996 643136 251048 643142
rect 250996 643078 251048 643084
rect 250904 630692 250956 630698
rect 250904 630634 250956 630640
rect 250812 616888 250864 616894
rect 250812 616830 250864 616836
rect 249708 590708 249760 590714
rect 249708 590650 249760 590656
rect 249616 576904 249668 576910
rect 249616 576846 249668 576852
rect 249524 563100 249576 563106
rect 249524 563042 249576 563048
rect 248328 536852 248380 536858
rect 248328 536794 248380 536800
rect 248236 524476 248288 524482
rect 248236 524418 248288 524424
rect 248144 510672 248196 510678
rect 248144 510614 248196 510620
rect 246948 484424 247000 484430
rect 246948 484366 247000 484372
rect 246856 456816 246908 456822
rect 246856 456758 246908 456764
rect 246764 430636 246816 430642
rect 246764 430578 246816 430584
rect 246672 418192 246724 418198
rect 246672 418134 246724 418140
rect 245568 404388 245620 404394
rect 245568 404330 245620 404336
rect 242164 391808 242216 391814
rect 242164 391750 242216 391756
rect 240784 391468 240836 391474
rect 240784 391410 240836 391416
rect 238024 391400 238076 391406
rect 238024 391342 238076 391348
rect 242808 390516 242860 390522
rect 242808 390458 242860 390464
rect 241796 390176 241848 390182
rect 241796 390118 241848 390124
rect 241428 390108 241480 390114
rect 241428 390050 241480 390056
rect 152464 390040 152516 390046
rect 152464 389982 152516 389988
rect 40776 389904 40828 389910
rect 40776 389846 40828 389852
rect 39396 389836 39448 389842
rect 39396 389778 39448 389784
rect 36636 389768 36688 389774
rect 36636 389710 36688 389716
rect 35256 389700 35308 389706
rect 35256 389642 35308 389648
rect 33784 389632 33836 389638
rect 33784 389574 33836 389580
rect 15844 389496 15896 389502
rect 15844 389438 15896 389444
rect 14648 388340 14700 388346
rect 14648 388282 14700 388288
rect 14556 388204 14608 388210
rect 14556 388146 14608 388152
rect 7564 388136 7616 388142
rect 7564 388078 7616 388084
rect 4804 388000 4856 388006
rect 4804 387942 4856 387948
rect 3424 387932 3476 387938
rect 3424 387874 3476 387880
rect 3332 371612 3384 371618
rect 3332 371554 3384 371560
rect 3344 371385 3372 371554
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3056 293956 3108 293962
rect 3056 293898 3108 293904
rect 3068 293185 3096 293898
rect 3054 293176 3110 293185
rect 3054 293111 3110 293120
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 2780 71664 2832 71670
rect 2778 71632 2780 71641
rect 2832 71632 2834 71641
rect 2778 71567 2834 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3436 32473 3464 387874
rect 3516 387048 3568 387054
rect 3516 386990 3568 386996
rect 3528 345409 3556 386990
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 3516 320136 3568 320142
rect 3516 320078 3568 320084
rect 3528 319297 3556 320078
rect 3514 319288 3570 319297
rect 3514 319223 3570 319232
rect 3516 306332 3568 306338
rect 3516 306274 3568 306280
rect 3528 306241 3556 306274
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 4816 71670 4844 387942
rect 7576 371618 7604 388078
rect 11796 388068 11848 388074
rect 11796 388010 11848 388016
rect 7564 371612 7616 371618
rect 7564 371554 7616 371560
rect 6828 335368 6880 335374
rect 6828 335310 6880 335316
rect 5448 324964 5500 324970
rect 5448 324906 5500 324912
rect 4804 71664 4856 71670
rect 4804 71606 4856 71612
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 5460 6914 5488 324906
rect 6840 6914 6868 335310
rect 11704 327820 11756 327826
rect 11704 327762 11756 327768
rect 10324 327752 10376 327758
rect 10324 327694 10376 327700
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 572 4072 624 4078
rect 572 4014 624 4020
rect 584 480 612 4014
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1688 480 1716 3946
rect 2872 3868 2924 3874
rect 2872 3810 2924 3816
rect 2884 480 2912 3810
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 480 4108 3402
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 7656 3800 7708 3806
rect 7656 3742 7708 3748
rect 7668 480 7696 3742
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8772 480 8800 3470
rect 9968 480 9996 3606
rect 10336 3534 10364 327694
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 11164 480 11192 3674
rect 11716 3466 11744 327762
rect 11808 111790 11836 388010
rect 14464 329112 14516 329118
rect 14464 329054 14516 329060
rect 11796 111784 11848 111790
rect 11796 111726 11848 111732
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12360 480 12388 2994
rect 13556 480 13584 4082
rect 14476 3058 14504 329054
rect 14568 164218 14596 388146
rect 14660 320142 14688 388282
rect 15856 358766 15884 389438
rect 21364 389428 21416 389434
rect 21364 389370 21416 389376
rect 18696 388476 18748 388482
rect 18696 388418 18748 388424
rect 17316 388408 17368 388414
rect 17316 388350 17368 388356
rect 17224 387116 17276 387122
rect 17224 387058 17276 387064
rect 15844 358760 15896 358766
rect 15844 358702 15896 358708
rect 15106 336016 15162 336025
rect 15106 335951 15162 335960
rect 14648 320136 14700 320142
rect 14648 320078 14700 320084
rect 14556 164212 14608 164218
rect 14556 164154 14608 164160
rect 15120 6914 15148 335951
rect 15198 335608 15254 335617
rect 15198 335543 15254 335552
rect 15212 16574 15240 335543
rect 16578 334656 16634 334665
rect 16578 334591 16634 334600
rect 16592 16574 16620 334591
rect 17236 85542 17264 387058
rect 17328 267714 17356 388350
rect 18604 388272 18656 388278
rect 18604 388214 18656 388220
rect 17316 267708 17368 267714
rect 17316 267650 17368 267656
rect 17224 85536 17276 85542
rect 17224 85478 17276 85484
rect 18616 45558 18644 388214
rect 18708 241466 18736 388418
rect 18696 241460 18748 241466
rect 18696 241402 18748 241408
rect 18604 45552 18656 45558
rect 18604 45494 18656 45500
rect 15212 16546 15976 16574
rect 16592 16546 17080 16574
rect 14752 6886 15148 6914
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14752 480 14780 6886
rect 15948 480 15976 16546
rect 17052 480 17080 16546
rect 21376 6866 21404 389370
rect 32496 389156 32548 389162
rect 32496 389098 32548 389104
rect 29644 388612 29696 388618
rect 29644 388554 29696 388560
rect 21456 388544 21508 388550
rect 21456 388486 21508 388492
rect 21468 189038 21496 388486
rect 24768 336116 24820 336122
rect 24768 336058 24820 336064
rect 22744 329180 22796 329186
rect 22744 329122 22796 329128
rect 21456 189032 21508 189038
rect 21456 188974 21508 188980
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 22756 4146 22784 329122
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18248 480 18276 3130
rect 19444 480 19472 3334
rect 20640 480 20668 3878
rect 23020 3596 23072 3602
rect 23020 3538 23072 3544
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 21836 480 21864 3402
rect 23032 480 23060 3538
rect 24780 3534 24808 336058
rect 24858 335472 24914 335481
rect 24858 335407 24914 335416
rect 24872 16574 24900 335407
rect 28998 333296 29054 333305
rect 28998 333231 29054 333240
rect 25502 330440 25558 330449
rect 25502 330375 25558 330384
rect 24872 16546 25360 16574
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 24228 480 24256 3470
rect 25332 480 25360 16546
rect 25516 3194 25544 330375
rect 26884 326392 26936 326398
rect 26884 326334 26936 326340
rect 26896 3670 26924 326334
rect 29012 16574 29040 333231
rect 29656 137970 29684 388554
rect 31666 336288 31722 336297
rect 31666 336223 31722 336232
rect 29644 137964 29696 137970
rect 29644 137906 29696 137912
rect 29012 16546 30144 16574
rect 27712 4140 27764 4146
rect 27712 4082 27764 4088
rect 26884 3664 26936 3670
rect 26884 3606 26936 3612
rect 26516 3324 26568 3330
rect 26516 3266 26568 3272
rect 25504 3188 25556 3194
rect 25504 3130 25556 3136
rect 26528 480 26556 3266
rect 27724 480 27752 4082
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 28920 480 28948 3606
rect 30116 480 30144 16546
rect 31680 6914 31708 336223
rect 32402 333432 32458 333441
rect 32402 333367 32458 333376
rect 32416 6914 32444 333367
rect 32508 215286 32536 389098
rect 33140 336796 33192 336802
rect 33140 336738 33192 336744
rect 33046 336424 33102 336433
rect 33046 336359 33102 336368
rect 32496 215280 32548 215286
rect 32496 215222 32548 215228
rect 31312 6886 31708 6914
rect 32324 6886 32444 6914
rect 31312 480 31340 6886
rect 32324 4078 32352 6886
rect 32312 4072 32364 4078
rect 32312 4014 32364 4020
rect 33060 3466 33088 336359
rect 33152 16574 33180 336738
rect 33796 97986 33824 389574
rect 35164 389564 35216 389570
rect 35164 389506 35216 389512
rect 33876 388680 33928 388686
rect 33876 388622 33928 388628
rect 33888 293962 33916 388622
rect 33876 293956 33928 293962
rect 33876 293898 33928 293904
rect 33784 97980 33836 97986
rect 33784 97922 33836 97928
rect 35176 59362 35204 389506
rect 35268 306338 35296 389642
rect 36542 331800 36598 331809
rect 36542 331735 36598 331744
rect 35256 306332 35308 306338
rect 35256 306274 35308 306280
rect 35164 59356 35216 59362
rect 35164 59298 35216 59304
rect 33152 16546 33640 16574
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 33048 3460 33100 3466
rect 33048 3402 33100 3408
rect 32416 480 32444 3402
rect 33612 480 33640 16546
rect 34796 4072 34848 4078
rect 34796 4014 34848 4020
rect 34808 480 34836 4014
rect 36556 4010 36584 331735
rect 36648 255270 36676 389710
rect 38566 336560 38622 336569
rect 38566 336495 38622 336504
rect 36636 255264 36688 255270
rect 36636 255206 36688 255212
rect 38580 6914 38608 336495
rect 39302 331936 39358 331945
rect 39302 331871 39358 331880
rect 38396 6886 38608 6914
rect 36544 4004 36596 4010
rect 36544 3946 36596 3952
rect 35992 3256 36044 3262
rect 35992 3198 36044 3204
rect 36004 480 36032 3198
rect 37188 2984 37240 2990
rect 37188 2926 37240 2932
rect 37200 480 37228 2926
rect 38396 480 38424 6886
rect 39316 3874 39344 331871
rect 39408 202842 39436 389778
rect 39948 336184 40000 336190
rect 39948 336126 40000 336132
rect 39396 202836 39448 202842
rect 39396 202778 39448 202784
rect 39960 6914 39988 336126
rect 40682 333568 40738 333577
rect 40682 333503 40738 333512
rect 40696 6914 40724 333503
rect 40788 150414 40816 389846
rect 103428 336728 103480 336734
rect 50986 336696 51042 336705
rect 103428 336670 103480 336676
rect 50986 336631 51042 336640
rect 96528 336660 96580 336666
rect 46848 336524 46900 336530
rect 46848 336466 46900 336472
rect 45468 336388 45520 336394
rect 45468 336330 45520 336336
rect 43442 332072 43498 332081
rect 43442 332007 43498 332016
rect 40776 150408 40828 150414
rect 40776 150350 40828 150356
rect 39592 6886 39988 6914
rect 40604 6886 40724 6914
rect 39304 3868 39356 3874
rect 39304 3810 39356 3816
rect 39592 480 39620 6886
rect 40604 3398 40632 6886
rect 43456 3874 43484 332007
rect 43536 331900 43588 331906
rect 43536 331842 43588 331848
rect 43444 3868 43496 3874
rect 43444 3810 43496 3816
rect 43076 3800 43128 3806
rect 43076 3742 43128 3748
rect 40592 3392 40644 3398
rect 40592 3334 40644 3340
rect 41880 3324 41932 3330
rect 41880 3266 41932 3272
rect 40684 3120 40736 3126
rect 40684 3062 40736 3068
rect 40696 480 40724 3062
rect 41892 480 41920 3266
rect 43088 480 43116 3742
rect 43548 2990 43576 331842
rect 44824 329248 44876 329254
rect 44824 329190 44876 329196
rect 44272 4004 44324 4010
rect 44272 3946 44324 3952
rect 43536 2984 43588 2990
rect 43536 2926 43588 2932
rect 44284 480 44312 3946
rect 44836 3126 44864 329190
rect 44824 3120 44876 3126
rect 44824 3062 44876 3068
rect 45480 480 45508 336330
rect 46204 329316 46256 329322
rect 46204 329258 46256 329264
rect 46216 4010 46244 329258
rect 46860 6914 46888 336466
rect 48226 333704 48282 333713
rect 48226 333639 48282 333648
rect 47584 326460 47636 326466
rect 47584 326402 47636 326408
rect 46676 6886 46888 6914
rect 46204 4004 46256 4010
rect 46204 3946 46256 3952
rect 46676 480 46704 6886
rect 47596 3262 47624 326402
rect 48240 6914 48268 333639
rect 50344 329384 50396 329390
rect 50344 329326 50396 329332
rect 47872 6886 48268 6914
rect 47584 3256 47636 3262
rect 47584 3198 47636 3204
rect 47872 480 47900 6886
rect 50160 3732 50212 3738
rect 50160 3674 50212 3680
rect 48964 3392 49016 3398
rect 48964 3334 49016 3340
rect 48976 480 49004 3334
rect 50172 480 50200 3674
rect 50356 3398 50384 329326
rect 50436 325712 50488 325718
rect 50436 325654 50488 325660
rect 50448 3806 50476 325654
rect 50436 3800 50488 3806
rect 50436 3742 50488 3748
rect 51000 3738 51028 336631
rect 96528 336602 96580 336608
rect 95148 336592 95200 336598
rect 95148 336534 95200 336540
rect 78588 336456 78640 336462
rect 78588 336398 78640 336404
rect 64788 336252 64840 336258
rect 64788 336194 64840 336200
rect 57886 335880 57942 335889
rect 57886 335815 57942 335824
rect 55126 334792 55182 334801
rect 55126 334727 55182 334736
rect 53102 332208 53158 332217
rect 53102 332143 53158 332152
rect 51724 327956 51776 327962
rect 51724 327898 51776 327904
rect 51736 4146 51764 327898
rect 51816 13116 51868 13122
rect 51816 13058 51868 13064
rect 51724 4140 51776 4146
rect 51724 4082 51776 4088
rect 51828 3874 51856 13058
rect 51816 3868 51868 3874
rect 51816 3810 51868 3816
rect 53116 3738 53144 332143
rect 53748 327888 53800 327894
rect 53748 327830 53800 327836
rect 50988 3732 51040 3738
rect 50988 3674 51040 3680
rect 51356 3732 51408 3738
rect 51356 3674 51408 3680
rect 53104 3732 53156 3738
rect 53104 3674 53156 3680
rect 53656 3732 53708 3738
rect 53656 3674 53708 3680
rect 50344 3392 50396 3398
rect 50344 3334 50396 3340
rect 51368 480 51396 3674
rect 52552 3392 52604 3398
rect 52552 3334 52604 3340
rect 52564 480 52592 3334
rect 53668 1850 53696 3674
rect 53760 3398 53788 327830
rect 55140 6914 55168 334727
rect 57244 328024 57296 328030
rect 57244 327966 57296 327972
rect 57256 6914 57284 327966
rect 54956 6886 55168 6914
rect 57164 6886 57284 6914
rect 53748 3392 53800 3398
rect 53748 3334 53800 3340
rect 53668 1822 53788 1850
rect 53760 480 53788 1822
rect 54956 480 54984 6886
rect 57164 3398 57192 6886
rect 57900 3398 57928 335815
rect 62026 330712 62082 330721
rect 62026 330647 62082 330656
rect 61382 330576 61438 330585
rect 61382 330511 61438 330520
rect 58624 326528 58676 326534
rect 58624 326470 58676 326476
rect 58636 4078 58664 326470
rect 58624 4072 58676 4078
rect 58624 4014 58676 4020
rect 60832 3800 60884 3806
rect 60832 3742 60884 3748
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 57152 3392 57204 3398
rect 57152 3334 57204 3340
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 57888 3392 57940 3398
rect 57888 3334 57940 3340
rect 59636 3392 59688 3398
rect 59636 3334 59688 3340
rect 56060 480 56088 3334
rect 57256 480 57284 3334
rect 58440 3052 58492 3058
rect 58440 2994 58492 3000
rect 58452 480 58480 2994
rect 59648 480 59676 3334
rect 60844 480 60872 3742
rect 61396 3058 61424 330511
rect 61384 3052 61436 3058
rect 61384 2994 61436 3000
rect 62040 480 62068 330647
rect 62764 328092 62816 328098
rect 62764 328034 62816 328040
rect 62776 3398 62804 328034
rect 63408 326596 63460 326602
rect 63408 326538 63460 326544
rect 63420 6914 63448 326538
rect 63236 6886 63448 6914
rect 62764 3392 62816 3398
rect 62764 3334 62816 3340
rect 63236 480 63264 6886
rect 64800 3398 64828 336194
rect 66166 332344 66222 332353
rect 66166 332279 66222 332288
rect 64328 3392 64380 3398
rect 64328 3334 64380 3340
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 64340 480 64368 3334
rect 66180 3194 66208 332279
rect 70306 330848 70362 330857
rect 70306 330783 70362 330792
rect 70216 328228 70268 328234
rect 70216 328170 70268 328176
rect 68284 328160 68336 328166
rect 68284 328102 68336 328108
rect 67916 4820 67968 4826
rect 67916 4762 67968 4768
rect 66720 3392 66772 3398
rect 66720 3334 66772 3340
rect 65524 3188 65576 3194
rect 65524 3130 65576 3136
rect 66168 3188 66220 3194
rect 66168 3130 66220 3136
rect 65536 480 65564 3130
rect 66732 480 66760 3334
rect 67928 480 67956 4762
rect 68296 3398 68324 328102
rect 70228 16574 70256 328170
rect 70136 16546 70256 16574
rect 69112 3868 69164 3874
rect 69112 3810 69164 3816
rect 68284 3392 68336 3398
rect 68284 3334 68336 3340
rect 69124 480 69152 3810
rect 70136 3482 70164 16546
rect 70320 6914 70348 330783
rect 73068 330540 73120 330546
rect 73068 330482 73120 330488
rect 70228 6886 70348 6914
rect 70228 3874 70256 6886
rect 70216 3868 70268 3874
rect 70216 3810 70268 3816
rect 71504 3868 71556 3874
rect 71504 3810 71556 3816
rect 70136 3454 70348 3482
rect 70320 480 70348 3454
rect 71516 480 71544 3810
rect 73080 3398 73108 330482
rect 77208 329452 77260 329458
rect 77208 329394 77260 329400
rect 75184 328296 75236 328302
rect 75184 328238 75236 328244
rect 75000 6180 75052 6186
rect 75000 6122 75052 6128
rect 72608 3392 72660 3398
rect 72608 3334 72660 3340
rect 73068 3392 73120 3398
rect 73068 3334 73120 3340
rect 72620 480 72648 3334
rect 73804 2984 73856 2990
rect 73804 2926 73856 2932
rect 73816 480 73844 2926
rect 75012 480 75040 6122
rect 75196 2990 75224 328238
rect 77220 3398 77248 329394
rect 76196 3392 76248 3398
rect 76196 3334 76248 3340
rect 77208 3392 77260 3398
rect 77208 3334 77260 3340
rect 75184 2984 75236 2990
rect 75184 2926 75236 2932
rect 76208 480 76236 3334
rect 77392 2984 77444 2990
rect 77392 2926 77444 2932
rect 77404 480 77432 2926
rect 78600 480 78628 336398
rect 89628 336320 89680 336326
rect 89628 336262 89680 336268
rect 81346 333840 81402 333849
rect 81346 333775 81402 333784
rect 79968 329520 80020 329526
rect 79968 329462 80020 329468
rect 79980 6914 80008 329462
rect 80704 328364 80756 328370
rect 80704 328306 80756 328312
rect 79704 6886 80008 6914
rect 79704 480 79732 6886
rect 80716 2990 80744 328306
rect 81360 3398 81388 333775
rect 88248 331968 88300 331974
rect 88248 331910 88300 331916
rect 84108 330608 84160 330614
rect 84108 330550 84160 330556
rect 83464 326664 83516 326670
rect 83464 326606 83516 326612
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 81348 3392 81400 3398
rect 81348 3334 81400 3340
rect 83280 3392 83332 3398
rect 83280 3334 83332 3340
rect 80704 2984 80756 2990
rect 80704 2926 80756 2932
rect 80900 480 80928 3334
rect 82084 3256 82136 3262
rect 82084 3198 82136 3204
rect 82096 480 82124 3198
rect 83292 480 83320 3334
rect 83476 3262 83504 326606
rect 84120 3398 84148 330550
rect 86868 329588 86920 329594
rect 86868 329530 86920 329536
rect 86224 328432 86276 328438
rect 86224 328374 86276 328380
rect 85672 4004 85724 4010
rect 85672 3946 85724 3952
rect 84108 3392 84160 3398
rect 84108 3334 84160 3340
rect 84476 3392 84528 3398
rect 84476 3334 84528 3340
rect 83464 3256 83516 3262
rect 83464 3198 83516 3204
rect 84488 480 84516 3334
rect 85684 480 85712 3946
rect 86236 3398 86264 328374
rect 86224 3392 86276 3398
rect 86224 3334 86276 3340
rect 86880 480 86908 329530
rect 88260 6914 88288 331910
rect 87984 6886 88288 6914
rect 87984 480 88012 6886
rect 89640 3398 89668 336262
rect 95056 329724 95108 329730
rect 95056 329666 95108 329672
rect 91008 329656 91060 329662
rect 91008 329598 91060 329604
rect 91020 3398 91048 329598
rect 93124 327684 93176 327690
rect 93124 327626 93176 327632
rect 92756 4072 92808 4078
rect 92756 4014 92808 4020
rect 89168 3392 89220 3398
rect 89168 3334 89220 3340
rect 89628 3392 89680 3398
rect 89628 3334 89680 3340
rect 90364 3392 90416 3398
rect 90364 3334 90416 3340
rect 91008 3392 91060 3398
rect 91008 3334 91060 3340
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 89180 480 89208 3334
rect 90376 480 90404 3334
rect 91572 480 91600 3334
rect 92768 480 92796 4014
rect 93136 3398 93164 327626
rect 95068 3398 95096 329666
rect 93124 3392 93176 3398
rect 93124 3334 93176 3340
rect 93952 3392 94004 3398
rect 93952 3334 94004 3340
rect 95056 3392 95108 3398
rect 95056 3334 95108 3340
rect 93964 480 93992 3334
rect 95160 480 95188 336534
rect 96540 6914 96568 336602
rect 102048 330676 102100 330682
rect 102048 330618 102100 330624
rect 97908 329792 97960 329798
rect 97908 329734 97960 329740
rect 96264 6886 96568 6914
rect 96264 480 96292 6886
rect 97920 3398 97948 329734
rect 99288 327616 99340 327622
rect 99288 327558 99340 327564
rect 99300 3398 99328 327558
rect 99840 4140 99892 4146
rect 99840 4082 99892 4088
rect 97448 3392 97500 3398
rect 97448 3334 97500 3340
rect 97908 3392 97960 3398
rect 97908 3334 97960 3340
rect 98644 3392 98696 3398
rect 98644 3334 98696 3340
rect 99288 3392 99340 3398
rect 99288 3334 99340 3340
rect 97460 480 97488 3334
rect 98656 480 98684 3334
rect 99852 480 99880 4082
rect 102060 3398 102088 330618
rect 103440 6914 103468 336670
rect 117228 335980 117280 335986
rect 117228 335922 117280 335928
rect 110328 331288 110380 331294
rect 110328 331230 110380 331236
rect 104808 329044 104860 329050
rect 104808 328986 104860 328992
rect 104820 6914 104848 328986
rect 108948 328976 109000 328982
rect 108948 328918 109000 328924
rect 106924 326868 106976 326874
rect 106924 326810 106976 326816
rect 106188 326732 106240 326738
rect 106188 326674 106240 326680
rect 103348 6886 103468 6914
rect 104544 6886 104848 6914
rect 101036 3392 101088 3398
rect 101036 3334 101088 3340
rect 102048 3392 102100 3398
rect 102048 3334 102100 3340
rect 102232 3392 102284 3398
rect 102232 3334 102284 3340
rect 101048 480 101076 3334
rect 102244 480 102272 3334
rect 103348 480 103376 6886
rect 104544 480 104572 6886
rect 106200 3262 106228 326674
rect 106936 6914 106964 326810
rect 107568 326800 107620 326806
rect 107568 326742 107620 326748
rect 106844 6886 106964 6914
rect 106844 3330 106872 6886
rect 107580 3330 107608 326742
rect 108960 3330 108988 328918
rect 110340 3330 110368 331230
rect 111708 328908 111760 328914
rect 111708 328850 111760 328856
rect 111720 6914 111748 328850
rect 115848 328840 115900 328846
rect 115848 328782 115900 328788
rect 115204 326936 115256 326942
rect 115204 326878 115256 326884
rect 113088 323604 113140 323610
rect 113088 323546 113140 323552
rect 113100 6914 113128 323546
rect 115216 6914 115244 326878
rect 111628 6886 111748 6914
rect 112824 6886 113128 6914
rect 115124 6886 115244 6914
rect 106832 3324 106884 3330
rect 106832 3266 106884 3272
rect 106924 3324 106976 3330
rect 106924 3266 106976 3272
rect 107568 3324 107620 3330
rect 107568 3266 107620 3272
rect 108120 3324 108172 3330
rect 108120 3266 108172 3272
rect 108948 3324 109000 3330
rect 108948 3266 109000 3272
rect 109316 3324 109368 3330
rect 109316 3266 109368 3272
rect 110328 3324 110380 3330
rect 110328 3266 110380 3272
rect 105728 3256 105780 3262
rect 105728 3198 105780 3204
rect 106188 3256 106240 3262
rect 106188 3198 106240 3204
rect 105740 480 105768 3198
rect 106936 480 106964 3266
rect 108132 480 108160 3266
rect 109328 480 109356 3266
rect 110512 2984 110564 2990
rect 110512 2926 110564 2932
rect 110524 480 110552 2926
rect 111628 480 111656 6886
rect 112824 480 112852 6886
rect 115124 3194 115152 6886
rect 115860 3330 115888 328782
rect 117240 3330 117268 335922
rect 119988 335912 120040 335918
rect 119988 335854 120040 335860
rect 119896 328772 119948 328778
rect 119896 328714 119948 328720
rect 119908 16574 119936 328714
rect 119816 16546 119936 16574
rect 119816 3330 119844 16546
rect 120000 6914 120028 335854
rect 140686 335200 140742 335209
rect 140686 335135 140742 335144
rect 136454 335064 136510 335073
rect 136454 334999 136510 335008
rect 129646 334928 129702 334937
rect 129646 334863 129702 334872
rect 128266 333976 128322 333985
rect 128266 333911 128322 333920
rect 128176 332104 128228 332110
rect 128176 332046 128228 332052
rect 122748 328704 122800 328710
rect 122748 328646 122800 328652
rect 119908 6886 120028 6914
rect 115204 3324 115256 3330
rect 115204 3266 115256 3272
rect 115848 3324 115900 3330
rect 115848 3266 115900 3272
rect 116400 3324 116452 3330
rect 116400 3266 116452 3272
rect 117228 3324 117280 3330
rect 117228 3266 117280 3272
rect 118792 3324 118844 3330
rect 118792 3266 118844 3272
rect 119804 3324 119856 3330
rect 119804 3266 119856 3272
rect 114008 3188 114060 3194
rect 114008 3130 114060 3136
rect 115112 3188 115164 3194
rect 115112 3130 115164 3136
rect 114020 480 114048 3130
rect 115216 480 115244 3266
rect 116412 480 116440 3266
rect 117596 3052 117648 3058
rect 117596 2994 117648 3000
rect 117608 480 117636 2994
rect 118804 480 118832 3266
rect 119908 480 119936 6886
rect 122760 3330 122788 328646
rect 125508 327072 125560 327078
rect 125508 327014 125560 327020
rect 124128 327004 124180 327010
rect 124128 326946 124180 326952
rect 124140 3330 124168 326946
rect 125520 3330 125548 327014
rect 122288 3324 122340 3330
rect 122288 3266 122340 3272
rect 122748 3324 122800 3330
rect 122748 3266 122800 3272
rect 123484 3324 123536 3330
rect 123484 3266 123536 3272
rect 124128 3324 124180 3330
rect 124128 3266 124180 3272
rect 124680 3324 124732 3330
rect 124680 3266 124732 3272
rect 125508 3324 125560 3330
rect 125508 3266 125560 3272
rect 126980 3324 127032 3330
rect 126980 3266 127032 3272
rect 121092 2848 121144 2854
rect 121092 2790 121144 2796
rect 121104 480 121132 2790
rect 122300 480 122328 3266
rect 123496 480 123524 3266
rect 124692 480 124720 3266
rect 125876 3256 125928 3262
rect 125876 3198 125928 3204
rect 125888 480 125916 3198
rect 126992 480 127020 3266
rect 128188 480 128216 332046
rect 128280 3330 128308 333911
rect 129660 6914 129688 334863
rect 131028 333260 131080 333266
rect 131028 333202 131080 333208
rect 129384 6886 129688 6914
rect 128268 3324 128320 3330
rect 128268 3266 128320 3272
rect 129384 480 129412 6886
rect 131040 3330 131068 333202
rect 135168 332172 135220 332178
rect 135168 332114 135220 332120
rect 132408 330744 132460 330750
rect 132408 330686 132460 330692
rect 132420 3330 132448 330686
rect 135180 3330 135208 332114
rect 135260 4888 135312 4894
rect 135260 4830 135312 4836
rect 130568 3324 130620 3330
rect 130568 3266 130620 3272
rect 131028 3324 131080 3330
rect 131028 3266 131080 3272
rect 131764 3324 131816 3330
rect 131764 3266 131816 3272
rect 132408 3324 132460 3330
rect 132408 3266 132460 3272
rect 134156 3324 134208 3330
rect 134156 3266 134208 3272
rect 135168 3324 135220 3330
rect 135168 3266 135220 3272
rect 130580 480 130608 3266
rect 131776 480 131804 3266
rect 132960 3188 133012 3194
rect 132960 3130 133012 3136
rect 132972 480 133000 3130
rect 134168 480 134196 3266
rect 135272 480 135300 4830
rect 136468 480 136496 334999
rect 137928 332240 137980 332246
rect 137928 332182 137980 332188
rect 137940 6914 137968 332182
rect 139308 330812 139360 330818
rect 139308 330754 139360 330760
rect 137664 6886 137968 6914
rect 137664 480 137692 6886
rect 139320 3330 139348 330754
rect 140700 3330 140728 335135
rect 151728 333532 151780 333538
rect 151728 333474 151780 333480
rect 148968 333396 149020 333402
rect 148968 333338 149020 333344
rect 147588 333328 147640 333334
rect 147588 333270 147640 333276
rect 144828 332376 144880 332382
rect 144828 332318 144880 332324
rect 142068 332308 142120 332314
rect 142068 332250 142120 332256
rect 138848 3324 138900 3330
rect 138848 3266 138900 3272
rect 139308 3324 139360 3330
rect 139308 3266 139360 3272
rect 140044 3324 140096 3330
rect 140044 3266 140096 3272
rect 140688 3324 140740 3330
rect 140688 3266 140740 3272
rect 138860 480 138888 3266
rect 140056 480 140084 3266
rect 142080 3194 142108 332250
rect 143448 330880 143500 330886
rect 143448 330822 143500 330828
rect 143460 3194 143488 330822
rect 144840 6914 144868 332318
rect 144748 6886 144868 6914
rect 141240 3188 141292 3194
rect 141240 3130 141292 3136
rect 142068 3188 142120 3194
rect 142068 3130 142120 3136
rect 142436 3188 142488 3194
rect 142436 3130 142488 3136
rect 143448 3188 143500 3194
rect 143448 3130 143500 3136
rect 141252 480 141280 3130
rect 142448 480 142476 3130
rect 143540 3120 143592 3126
rect 143540 3062 143592 3068
rect 143552 480 143580 3062
rect 144748 480 144776 6886
rect 145932 4956 145984 4962
rect 145932 4898 145984 4904
rect 145944 480 145972 4898
rect 147600 3194 147628 333270
rect 148980 3194 149008 333338
rect 150348 330948 150400 330954
rect 150348 330890 150400 330896
rect 150360 3194 150388 330890
rect 147128 3188 147180 3194
rect 147128 3130 147180 3136
rect 147588 3188 147640 3194
rect 147588 3130 147640 3136
rect 148324 3188 148376 3194
rect 148324 3130 148376 3136
rect 148968 3188 149020 3194
rect 148968 3130 149020 3136
rect 149520 3188 149572 3194
rect 149520 3130 149572 3136
rect 150348 3188 150400 3194
rect 150348 3130 150400 3136
rect 147140 480 147168 3130
rect 148336 480 148364 3130
rect 149532 480 149560 3130
rect 151740 3126 151768 333474
rect 152476 20670 152504 389982
rect 240690 389600 240746 389609
rect 240690 389535 240746 389544
rect 235906 389464 235962 389473
rect 235906 389399 235962 389408
rect 235816 389020 235868 389026
rect 235816 388962 235868 388968
rect 235448 388816 235500 388822
rect 235448 388758 235500 388764
rect 235460 387954 235488 388758
rect 235828 387954 235856 388962
rect 235244 387926 235488 387954
rect 235612 387926 235856 387954
rect 235920 387954 235948 389399
rect 238390 389328 238446 389337
rect 238390 389263 238446 389272
rect 240048 389292 240100 389298
rect 236552 389088 236604 389094
rect 236552 389030 236604 389036
rect 236564 387954 236592 389030
rect 236920 388952 236972 388958
rect 236920 388894 236972 388900
rect 236932 387954 236960 388894
rect 237656 388884 237708 388890
rect 237656 388826 237708 388832
rect 237668 387954 237696 388826
rect 238404 387954 238432 389263
rect 240048 389234 240100 389240
rect 239494 389192 239550 389201
rect 239494 389127 239550 389136
rect 239508 387954 239536 389127
rect 235920 387926 235980 387954
rect 236348 387926 236592 387954
rect 236716 387926 236960 387954
rect 237452 387926 237696 387954
rect 238188 387926 238432 387954
rect 239292 387926 239536 387954
rect 240060 387954 240088 389234
rect 240704 387954 240732 389535
rect 241440 387954 241468 390050
rect 241808 387954 241836 390118
rect 242532 389360 242584 389366
rect 242532 389302 242584 389308
rect 242544 387954 242572 389302
rect 242820 387954 242848 390458
rect 244004 390380 244056 390386
rect 244004 390322 244056 390328
rect 243636 388748 243688 388754
rect 243636 388690 243688 388696
rect 243648 387954 243676 388690
rect 244016 387954 244044 390322
rect 245200 390244 245252 390250
rect 245200 390186 245252 390192
rect 245212 387954 245240 390186
rect 245580 387954 245608 404330
rect 245936 390448 245988 390454
rect 245936 390390 245988 390396
rect 245948 387954 245976 390390
rect 246684 389174 246712 418134
rect 246776 390454 246804 430578
rect 246764 390448 246816 390454
rect 246764 390390 246816 390396
rect 246316 389146 246712 389174
rect 246316 387954 246344 389146
rect 246868 388090 246896 456758
rect 246684 388062 246896 388090
rect 246684 387954 246712 388062
rect 246960 387954 246988 484366
rect 248052 470620 248104 470626
rect 248052 470562 248104 470568
rect 248064 390454 248092 470562
rect 247408 390448 247460 390454
rect 247408 390390 247460 390396
rect 248052 390448 248104 390454
rect 248052 390390 248104 390396
rect 247420 387954 247448 390390
rect 248156 390266 248184 510614
rect 247788 390238 248184 390266
rect 247788 387954 247816 390238
rect 248144 389972 248196 389978
rect 248144 389914 248196 389920
rect 248156 387954 248184 389914
rect 240060 387926 240120 387954
rect 240488 387926 240732 387954
rect 241224 387926 241468 387954
rect 241592 387926 241836 387954
rect 242328 387926 242572 387954
rect 242696 387926 242848 387954
rect 243432 387926 243676 387954
rect 243800 387926 244044 387954
rect 244996 387926 245240 387954
rect 245364 387926 245608 387954
rect 245732 387926 245976 387954
rect 246100 387926 246344 387954
rect 246468 387926 246712 387954
rect 246836 387926 246988 387954
rect 247204 387926 247448 387954
rect 247572 387926 247816 387954
rect 247940 387926 248184 387954
rect 248248 387954 248276 524418
rect 248340 389978 248368 536794
rect 249536 390454 249564 563042
rect 248972 390448 249024 390454
rect 248972 390390 249024 390396
rect 249524 390448 249576 390454
rect 249524 390390 249576 390396
rect 248328 389972 248380 389978
rect 248328 389914 248380 389920
rect 248984 387954 249012 390390
rect 249340 390380 249392 390386
rect 249340 390322 249392 390328
rect 249352 387954 249380 390322
rect 249628 387954 249656 576846
rect 249720 390386 249748 590650
rect 250824 402974 250852 616830
rect 250732 402946 250852 402974
rect 250732 390454 250760 402946
rect 250076 390448 250128 390454
rect 250076 390390 250128 390396
rect 250720 390448 250772 390454
rect 250720 390390 250772 390396
rect 249708 390380 249760 390386
rect 249708 390322 249760 390328
rect 250088 387954 250116 390390
rect 250444 390380 250496 390386
rect 250444 390322 250496 390328
rect 250456 387954 250484 390322
rect 250916 389174 250944 630634
rect 251008 390386 251036 643078
rect 250996 390380 251048 390386
rect 250996 390322 251048 390328
rect 250824 389146 250944 389174
rect 250824 387954 250852 389146
rect 251100 387954 251128 670686
rect 252008 391332 252060 391338
rect 252008 391274 252060 391280
rect 251916 390448 251968 390454
rect 251916 390390 251968 390396
rect 251548 390380 251600 390386
rect 251548 390322 251600 390328
rect 251560 387954 251588 390322
rect 251928 387954 251956 390390
rect 248248 387926 248308 387954
rect 248676 387926 249012 387954
rect 249136 387926 249380 387954
rect 249504 387926 249656 387954
rect 249872 387926 250116 387954
rect 250240 387926 250484 387954
rect 250608 387926 250852 387954
rect 250976 387926 251128 387954
rect 251344 387926 251588 387954
rect 251712 387926 251956 387954
rect 243268 387864 243320 387870
rect 243064 387812 243268 387818
rect 243064 387806 243320 387812
rect 252020 387818 252048 391274
rect 252204 387954 252232 700402
rect 252376 696992 252428 696998
rect 252376 696934 252428 696940
rect 252284 683188 252336 683194
rect 252284 683130 252336 683136
rect 252296 390454 252324 683130
rect 252284 390448 252336 390454
rect 252284 390390 252336 390396
rect 252388 390386 252416 696934
rect 253480 391264 253532 391270
rect 253480 391206 253532 391212
rect 253020 390448 253072 390454
rect 253020 390390 253072 390396
rect 252376 390380 252428 390386
rect 252376 390322 252428 390328
rect 253032 387954 253060 390390
rect 253492 387954 253520 391206
rect 253676 388226 253704 700674
rect 253756 700324 253808 700330
rect 253756 700266 253808 700272
rect 253768 390454 253796 700266
rect 254584 391536 254636 391542
rect 254584 391478 254636 391484
rect 253756 390448 253808 390454
rect 253756 390390 253808 390396
rect 254216 390448 254268 390454
rect 254216 390390 254268 390396
rect 252204 387926 252448 387954
rect 252816 387926 253060 387954
rect 253184 387926 253520 387954
rect 253630 388198 253704 388226
rect 253630 387940 253658 388198
rect 254228 387954 254256 390390
rect 254596 387954 254624 391478
rect 254964 387954 254992 700946
rect 255044 700936 255096 700942
rect 255044 700878 255096 700884
rect 254012 387926 254256 387954
rect 254380 387926 254624 387954
rect 254748 387926 254992 387954
rect 255056 387954 255084 700878
rect 259644 700868 259696 700874
rect 259644 700810 259696 700816
rect 255136 700596 255188 700602
rect 255136 700538 255188 700544
rect 255148 390454 255176 700538
rect 258172 700256 258224 700262
rect 258172 700198 258224 700204
rect 256424 700120 256476 700126
rect 256424 700062 256476 700068
rect 255688 391740 255740 391746
rect 255688 391682 255740 391688
rect 255136 390448 255188 390454
rect 255136 390390 255188 390396
rect 255700 387954 255728 391682
rect 256056 390448 256108 390454
rect 256056 390390 256108 390396
rect 256068 387954 256096 390390
rect 256436 387954 256464 700062
rect 256516 700052 256568 700058
rect 256516 699994 256568 700000
rect 256528 390454 256556 699994
rect 257896 699848 257948 699854
rect 257896 699790 257948 699796
rect 257908 393314 257936 699790
rect 257988 699780 258040 699786
rect 257988 699722 258040 699728
rect 257540 393286 257936 393314
rect 256608 391604 256660 391610
rect 256608 391546 256660 391552
rect 256516 390448 256568 390454
rect 256516 390390 256568 390396
rect 256620 388090 256648 391546
rect 257160 390516 257212 390522
rect 257160 390458 257212 390464
rect 255056 387926 255116 387954
rect 255484 387926 255728 387954
rect 255852 387926 256096 387954
rect 256220 387926 256464 387954
rect 256528 388062 256648 388090
rect 256528 387818 256556 388062
rect 257172 387954 257200 390458
rect 257540 387954 257568 393286
rect 257620 391400 257672 391406
rect 257620 391342 257672 391348
rect 256956 387926 257200 387954
rect 257324 387926 257568 387954
rect 257632 387954 257660 391342
rect 258000 390522 258028 699722
rect 258184 390522 258212 700198
rect 259552 700188 259604 700194
rect 259552 700130 259604 700136
rect 258264 699984 258316 699990
rect 258264 699926 258316 699932
rect 257988 390516 258040 390522
rect 257988 390458 258040 390464
rect 258172 390516 258224 390522
rect 258172 390458 258224 390464
rect 258276 387954 258304 699926
rect 258356 699916 258408 699922
rect 258356 699858 258408 699864
rect 257632 387926 257692 387954
rect 258152 387926 258304 387954
rect 258368 387954 258396 699858
rect 258632 391468 258684 391474
rect 258632 391410 258684 391416
rect 258644 387954 258672 391410
rect 259000 390516 259052 390522
rect 259000 390458 259052 390464
rect 259012 387954 259040 390458
rect 259564 387954 259592 700130
rect 259656 390522 259684 700810
rect 259736 700800 259788 700806
rect 259736 700742 259788 700748
rect 259748 402974 259776 700742
rect 260840 700664 260892 700670
rect 260840 700606 260892 700612
rect 259748 402946 260144 402974
rect 259736 391808 259788 391814
rect 259736 391750 259788 391756
rect 259644 390516 259696 390522
rect 259644 390458 259696 390464
rect 259748 387954 259776 391750
rect 260116 387954 260144 402946
rect 260472 390516 260524 390522
rect 260472 390458 260524 390464
rect 260484 387954 260512 390458
rect 260852 387954 260880 700606
rect 261024 700528 261076 700534
rect 261024 700470 261076 700476
rect 260932 700392 260984 700398
rect 260932 700334 260984 700340
rect 260944 388090 260972 700334
rect 261036 393314 261064 700470
rect 267660 699786 267688 703520
rect 273904 700868 273956 700874
rect 273904 700810 273956 700816
rect 271144 700800 271196 700806
rect 271144 700742 271196 700748
rect 269764 700664 269816 700670
rect 269764 700606 269816 700612
rect 267648 699780 267700 699786
rect 267648 699722 267700 699728
rect 261116 683256 261168 683262
rect 261116 683198 261168 683204
rect 261128 402974 261156 683198
rect 262220 670812 262272 670818
rect 262220 670754 262272 670760
rect 261128 402946 261984 402974
rect 261036 393286 261616 393314
rect 260944 388062 261248 388090
rect 261220 387954 261248 388062
rect 261588 387954 261616 393286
rect 261956 387954 261984 402946
rect 262232 390522 262260 670754
rect 262312 656940 262364 656946
rect 262312 656882 262364 656888
rect 262220 390516 262272 390522
rect 262220 390458 262272 390464
rect 262324 387954 262352 656882
rect 262404 632120 262456 632126
rect 262404 632062 262456 632068
rect 262416 402974 262444 632062
rect 263600 618316 263652 618322
rect 263600 618258 263652 618264
rect 262416 402946 263180 402974
rect 262772 390516 262824 390522
rect 262772 390458 262824 390464
rect 262784 387954 262812 390458
rect 263152 387954 263180 402946
rect 258368 387926 258520 387954
rect 258644 387926 258888 387954
rect 259012 387926 259256 387954
rect 259564 387926 259624 387954
rect 259748 387926 259992 387954
rect 260116 387926 260360 387954
rect 260484 387926 260728 387954
rect 260852 387926 261096 387954
rect 261220 387926 261464 387954
rect 261588 387926 261832 387954
rect 261956 387926 262200 387954
rect 262324 387926 262660 387954
rect 262784 387926 263028 387954
rect 263152 387926 263396 387954
rect 243064 387790 243308 387806
rect 252020 387790 252080 387818
rect 256528 387790 256588 387818
rect 263612 387802 263640 618258
rect 263692 605872 263744 605878
rect 263692 605814 263744 605820
rect 263704 387954 263732 605814
rect 263784 579692 263836 579698
rect 263784 579634 263836 579640
rect 263796 388090 263824 579634
rect 264980 565888 265032 565894
rect 264980 565830 265032 565836
rect 263876 553444 263928 553450
rect 263876 553386 263928 553392
rect 263888 402974 263916 553386
rect 263888 402946 264652 402974
rect 263796 388062 264284 388090
rect 264256 387954 264284 388062
rect 264624 387954 264652 402946
rect 264992 387954 265020 565830
rect 265072 527196 265124 527202
rect 265072 527138 265124 527144
rect 265084 388090 265112 527138
rect 265164 514820 265216 514826
rect 265164 514762 265216 514768
rect 265176 390522 265204 514762
rect 265256 501016 265308 501022
rect 265256 500958 265308 500964
rect 265268 402974 265296 500958
rect 266360 474768 266412 474774
rect 266360 474710 266412 474716
rect 265268 402946 265756 402974
rect 265164 390516 265216 390522
rect 265164 390458 265216 390464
rect 265084 388062 265388 388090
rect 265360 387954 265388 388062
rect 265728 387954 265756 402946
rect 266084 390516 266136 390522
rect 266084 390458 266136 390464
rect 266096 387954 266124 390458
rect 266372 388090 266400 474710
rect 266452 462392 266504 462398
rect 266452 462334 266504 462340
rect 266464 390522 266492 462334
rect 266544 448588 266596 448594
rect 266544 448530 266596 448536
rect 266556 402974 266584 448530
rect 267740 422340 267792 422346
rect 267740 422282 267792 422288
rect 266556 402946 266860 402974
rect 266452 390516 266504 390522
rect 266452 390458 266504 390464
rect 266372 388062 266492 388090
rect 266464 387954 266492 388062
rect 266832 387954 266860 402946
rect 267280 390516 267332 390522
rect 267280 390458 267332 390464
rect 267292 387954 267320 390458
rect 267752 387954 267780 422282
rect 267832 409896 267884 409902
rect 267832 409838 267884 409844
rect 267844 390522 267872 409838
rect 268016 397520 268068 397526
rect 268016 397462 268068 397468
rect 267832 390516 267884 390522
rect 267832 390458 267884 390464
rect 268028 387954 268056 397462
rect 269776 391814 269804 700606
rect 269764 391808 269816 391814
rect 269764 391750 269816 391756
rect 271156 391746 271184 700742
rect 271144 391740 271196 391746
rect 271144 391682 271196 391688
rect 273916 391610 273944 700810
rect 282184 700528 282236 700534
rect 282184 700470 282236 700476
rect 280804 700392 280856 700398
rect 280804 700334 280856 700340
rect 273904 391604 273956 391610
rect 273904 391546 273956 391552
rect 280816 391338 280844 700334
rect 280804 391332 280856 391338
rect 280804 391274 280856 391280
rect 282196 391270 282224 700470
rect 283852 699854 283880 703520
rect 300136 700874 300164 703520
rect 300124 700868 300176 700874
rect 300124 700810 300176 700816
rect 332520 700058 332548 703520
rect 348804 700126 348832 703520
rect 364996 700806 365024 703520
rect 397472 701010 397500 703520
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 413664 700942 413692 703520
rect 413652 700936 413704 700942
rect 413652 700878 413704 700884
rect 364984 700800 365036 700806
rect 364984 700742 365036 700748
rect 429856 700670 429884 703520
rect 462332 700738 462360 703520
rect 462320 700732 462372 700738
rect 462320 700674 462372 700680
rect 429844 700664 429896 700670
rect 429844 700606 429896 700612
rect 478524 700602 478552 703520
rect 478512 700596 478564 700602
rect 478512 700538 478564 700544
rect 494808 700534 494836 703520
rect 494796 700528 494848 700534
rect 494796 700470 494848 700476
rect 527192 700466 527220 703520
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 543476 700330 543504 703520
rect 559668 700398 559696 703520
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 348792 700120 348844 700126
rect 348792 700062 348844 700068
rect 332508 700052 332560 700058
rect 332508 699994 332560 700000
rect 283840 699848 283892 699854
rect 283840 699790 283892 699796
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 282184 391264 282236 391270
rect 282184 391206 282236 391212
rect 268384 390516 268436 390522
rect 268384 390458 268436 390464
rect 280896 390516 280948 390522
rect 280896 390458 280948 390464
rect 291936 390516 291988 390522
rect 291936 390458 291988 390464
rect 268396 387954 268424 390458
rect 277492 390040 277544 390046
rect 277492 389982 277544 389988
rect 273996 389904 274048 389910
rect 273996 389846 274048 389852
rect 272892 389836 272944 389842
rect 272892 389778 272944 389784
rect 271880 389768 271932 389774
rect 271880 389710 271932 389716
rect 270592 389700 270644 389706
rect 270592 389642 270644 389648
rect 269488 389496 269540 389502
rect 269488 389438 269540 389444
rect 268982 388136 269034 388142
rect 268982 388078 269034 388084
rect 263704 387926 263764 387954
rect 264256 387926 264500 387954
rect 264624 387926 264868 387954
rect 264992 387926 265236 387954
rect 265360 387926 265604 387954
rect 265728 387926 265972 387954
rect 266096 387926 266340 387954
rect 266464 387926 266708 387954
rect 266832 387926 267168 387954
rect 267292 387926 267536 387954
rect 267752 387926 267904 387954
rect 268028 387926 268272 387954
rect 268396 387926 268640 387954
rect 268994 387940 269022 388078
rect 269500 387954 269528 389438
rect 270224 388680 270276 388686
rect 270224 388622 270276 388628
rect 269856 388340 269908 388346
rect 269856 388282 269908 388288
rect 269868 387954 269896 388282
rect 270236 387954 270264 388622
rect 270604 387954 270632 389642
rect 271328 388476 271380 388482
rect 271328 388418 271380 388424
rect 270960 388408 271012 388414
rect 270960 388350 271012 388356
rect 270972 387954 271000 388350
rect 271340 387954 271368 388418
rect 271892 387954 271920 389710
rect 272156 389156 272208 389162
rect 272156 389098 272208 389104
rect 272168 387954 272196 389098
rect 272524 388544 272576 388550
rect 272524 388486 272576 388492
rect 272536 387954 272564 388486
rect 272904 387954 272932 389778
rect 273628 388612 273680 388618
rect 273628 388554 273680 388560
rect 273490 388204 273542 388210
rect 273490 388146 273542 388152
rect 269500 387926 269744 387954
rect 269868 387926 270112 387954
rect 270236 387926 270480 387954
rect 270604 387926 270848 387954
rect 270972 387926 271216 387954
rect 271340 387926 271676 387954
rect 271892 387926 272044 387954
rect 272168 387926 272412 387954
rect 272536 387926 272780 387954
rect 272904 387926 273148 387954
rect 273502 387940 273530 388146
rect 273640 387954 273668 388554
rect 274008 387954 274036 389846
rect 275100 389632 275152 389638
rect 275100 389574 275152 389580
rect 274364 388068 274416 388074
rect 274364 388010 274416 388016
rect 274376 387954 274404 388010
rect 275112 387954 275140 389574
rect 276296 389564 276348 389570
rect 276296 389506 276348 389512
rect 276020 388272 276072 388278
rect 276020 388214 276072 388220
rect 275468 388000 275520 388006
rect 273640 387926 273884 387954
rect 274008 387926 274252 387954
rect 274376 387926 274620 387954
rect 275112 387926 275356 387954
rect 276032 387954 276060 388214
rect 276308 387954 276336 389506
rect 277032 389428 277084 389434
rect 277032 389370 277084 389376
rect 277044 387954 277072 389370
rect 277504 387954 277532 389982
rect 279700 389768 279752 389774
rect 279700 389710 279752 389716
rect 278688 389632 278740 389638
rect 278688 389574 278740 389580
rect 277998 388136 278050 388142
rect 277998 388078 278050 388084
rect 275520 387948 275724 387954
rect 275468 387942 275724 387948
rect 275480 387926 275724 387942
rect 276032 387926 276184 387954
rect 276308 387926 276552 387954
rect 276676 387938 276920 387954
rect 276664 387932 276920 387938
rect 276716 387926 276920 387932
rect 277044 387926 277288 387954
rect 277504 387926 277656 387954
rect 278010 387940 278038 388078
rect 278596 388068 278648 388074
rect 278596 388010 278648 388016
rect 278608 387954 278636 388010
rect 278392 387926 278636 387954
rect 278700 387954 278728 389574
rect 279332 389360 279384 389366
rect 279332 389302 279384 389308
rect 279344 387954 279372 389302
rect 279712 387954 279740 389710
rect 280068 389564 280120 389570
rect 280068 389506 280120 389512
rect 280080 387954 280108 389506
rect 280528 388000 280580 388006
rect 278700 387926 278760 387954
rect 279128 387926 279372 387954
rect 279496 387926 279740 387954
rect 279864 387926 280108 387954
rect 280232 387948 280528 387954
rect 280908 387954 280936 390458
rect 285128 390176 285180 390182
rect 285128 390118 285180 390124
rect 286508 390176 286560 390182
rect 286508 390118 286560 390124
rect 289084 390176 289136 390182
rect 289084 390118 289136 390124
rect 285036 390108 285088 390114
rect 285036 390050 285088 390056
rect 282368 390040 282420 390046
rect 282368 389982 282420 389988
rect 281356 389904 281408 389910
rect 281356 389846 281408 389852
rect 281264 389836 281316 389842
rect 281264 389778 281316 389784
rect 281276 387954 281304 389778
rect 280232 387942 280580 387948
rect 280232 387926 280568 387942
rect 280692 387926 280936 387954
rect 281060 387926 281304 387954
rect 276664 387874 276716 387880
rect 281368 387818 281396 389846
rect 282380 387954 282408 389982
rect 282736 389700 282788 389706
rect 282736 389642 282788 389648
rect 282748 387954 282776 389642
rect 284576 389496 284628 389502
rect 284576 389438 284628 389444
rect 282828 389428 282880 389434
rect 282828 389370 282880 389376
rect 281796 387938 282040 387954
rect 281796 387932 282052 387938
rect 281796 387926 282000 387932
rect 282164 387926 282408 387954
rect 282532 387926 282776 387954
rect 282840 387954 282868 389370
rect 284208 389292 284260 389298
rect 284208 389234 284260 389240
rect 283472 389224 283524 389230
rect 283472 389166 283524 389172
rect 283484 387954 283512 389166
rect 284220 387954 284248 389234
rect 284588 387954 284616 389438
rect 285048 387954 285076 390050
rect 282840 387926 282900 387954
rect 283268 387926 283512 387954
rect 284004 387926 284248 387954
rect 284372 387926 284616 387954
rect 284740 387926 285076 387954
rect 282000 387874 282052 387880
rect 263888 387802 264132 387818
rect 263600 387796 263652 387802
rect 263600 387738 263652 387744
rect 263876 387796 264132 387802
rect 263928 387790 264132 387796
rect 281368 387790 281428 387818
rect 263876 387738 263928 387744
rect 237288 387320 237340 387326
rect 237084 387268 237288 387274
rect 238024 387320 238076 387326
rect 237084 387262 237340 387268
rect 237820 387268 238024 387274
rect 238668 387320 238720 387326
rect 237820 387262 238076 387268
rect 238556 387268 238668 387274
rect 239128 387320 239180 387326
rect 238556 387262 238720 387268
rect 238924 387268 239128 387274
rect 239956 387320 240008 387326
rect 238924 387262 239180 387268
rect 239660 387268 239956 387274
rect 241060 387320 241112 387326
rect 239660 387262 240008 387268
rect 240856 387268 241060 387274
rect 242164 387320 242216 387326
rect 240856 387262 241112 387268
rect 241960 387268 242164 387274
rect 244280 387320 244332 387326
rect 241960 387262 242216 387268
rect 244168 387268 244280 387274
rect 244832 387320 244884 387326
rect 244168 387262 244332 387268
rect 244628 387268 244832 387274
rect 244628 387262 244884 387268
rect 269120 387320 269172 387326
rect 274732 387320 274784 387326
rect 269172 387268 269376 387274
rect 269120 387262 269376 387268
rect 283840 387320 283892 387326
rect 274784 387268 274988 387274
rect 274732 387262 274988 387268
rect 237084 387246 237328 387262
rect 237820 387246 238064 387262
rect 238556 387246 238708 387262
rect 238924 387246 239168 387262
rect 239660 387246 239996 387262
rect 240856 387246 241100 387262
rect 241960 387246 242204 387262
rect 244168 387246 244320 387262
rect 244628 387246 244872 387262
rect 269132 387246 269376 387262
rect 274744 387246 274988 387262
rect 283636 387268 283840 387274
rect 283636 387262 283892 387268
rect 283636 387246 283880 387262
rect 233146 387016 233202 387025
rect 233146 386951 233202 386960
rect 232778 385112 232834 385121
rect 232778 385047 232834 385056
rect 232686 379400 232742 379409
rect 232686 379335 232742 379344
rect 232594 373552 232650 373561
rect 232594 373487 232650 373496
rect 232502 364032 232558 364041
rect 232502 363967 232558 363976
rect 232318 358184 232374 358193
rect 232318 358119 232374 358128
rect 232226 352472 232282 352481
rect 232226 352407 232282 352416
rect 232136 349852 232188 349858
rect 232136 349794 232188 349800
rect 232042 342816 232098 342825
rect 232042 342751 232098 342760
rect 171784 335844 171836 335850
rect 171784 335786 171836 335792
rect 158626 335336 158682 335345
rect 158626 335271 158682 335280
rect 154488 333464 154540 333470
rect 154488 333406 154540 333412
rect 153108 332444 153160 332450
rect 153108 332386 153160 332392
rect 153016 331016 153068 331022
rect 153016 330958 153068 330964
rect 152464 20664 152516 20670
rect 152464 20606 152516 20612
rect 150624 3120 150676 3126
rect 150624 3062 150676 3068
rect 151728 3120 151780 3126
rect 151728 3062 151780 3068
rect 151820 3120 151872 3126
rect 151820 3062 151872 3068
rect 150636 480 150664 3062
rect 151832 480 151860 3062
rect 153028 480 153056 330958
rect 153120 3126 153148 332386
rect 154500 6914 154528 333406
rect 155868 332512 155920 332518
rect 155868 332454 155920 332460
rect 154224 6886 154528 6914
rect 153108 3120 153160 3126
rect 153108 3062 153160 3068
rect 154224 480 154252 6886
rect 155880 3126 155908 332454
rect 157248 331084 157300 331090
rect 157248 331026 157300 331032
rect 157260 3126 157288 331026
rect 158640 3126 158668 335271
rect 169668 334756 169720 334762
rect 169668 334698 169720 334704
rect 165528 334620 165580 334626
rect 165528 334562 165580 334568
rect 162768 333600 162820 333606
rect 162768 333542 162820 333548
rect 160008 332580 160060 332586
rect 160008 332522 160060 332528
rect 160020 3126 160048 332522
rect 161388 328636 161440 328642
rect 161388 328578 161440 328584
rect 161400 3126 161428 328578
rect 162780 6914 162808 333542
rect 164148 331832 164200 331838
rect 164148 331774 164200 331780
rect 162504 6886 162808 6914
rect 155408 3120 155460 3126
rect 155408 3062 155460 3068
rect 155868 3120 155920 3126
rect 155868 3062 155920 3068
rect 156604 3120 156656 3126
rect 156604 3062 156656 3068
rect 157248 3120 157300 3126
rect 157248 3062 157300 3068
rect 157800 3120 157852 3126
rect 157800 3062 157852 3068
rect 158628 3120 158680 3126
rect 158628 3062 158680 3068
rect 158904 3120 158956 3126
rect 158904 3062 158956 3068
rect 160008 3120 160060 3126
rect 160008 3062 160060 3068
rect 160100 3120 160152 3126
rect 160100 3062 160152 3068
rect 161388 3120 161440 3126
rect 161388 3062 161440 3068
rect 155420 480 155448 3062
rect 156616 480 156644 3062
rect 157812 480 157840 3062
rect 158916 480 158944 3062
rect 160112 480 160140 3062
rect 161572 2984 161624 2990
rect 161308 2932 161572 2938
rect 161308 2926 161624 2932
rect 161308 2910 161612 2926
rect 161308 480 161336 2910
rect 162504 480 162532 6886
rect 164160 3126 164188 331774
rect 165540 3126 165568 334562
rect 169576 333736 169628 333742
rect 169576 333678 169628 333684
rect 166908 333668 166960 333674
rect 166908 333610 166960 333616
rect 166920 3126 166948 333610
rect 168288 331764 168340 331770
rect 168288 331706 168340 331712
rect 168300 3126 168328 331706
rect 163688 3120 163740 3126
rect 163688 3062 163740 3068
rect 164148 3120 164200 3126
rect 164148 3062 164200 3068
rect 164884 3120 164936 3126
rect 164884 3062 164936 3068
rect 165528 3120 165580 3126
rect 165528 3062 165580 3068
rect 166080 3120 166132 3126
rect 166080 3062 166132 3068
rect 166908 3120 166960 3126
rect 166908 3062 166960 3068
rect 167184 3120 167236 3126
rect 167184 3062 167236 3068
rect 168288 3120 168340 3126
rect 168288 3062 168340 3068
rect 168380 3120 168432 3126
rect 168380 3062 168432 3068
rect 163700 480 163728 3062
rect 164896 480 164924 3062
rect 166092 480 166120 3062
rect 167196 480 167224 3062
rect 168392 480 168420 3062
rect 169588 480 169616 333678
rect 169680 3126 169708 334698
rect 171048 331152 171100 331158
rect 171048 331094 171100 331100
rect 171060 6914 171088 331094
rect 170784 6886 171088 6914
rect 169668 3120 169720 3126
rect 169668 3062 169720 3068
rect 170784 480 170812 6886
rect 171796 2922 171824 335786
rect 178684 335776 178736 335782
rect 178684 335718 178736 335724
rect 176568 334688 176620 334694
rect 176568 334630 176620 334636
rect 173808 333804 173860 333810
rect 173808 333746 173860 333752
rect 173820 6914 173848 333746
rect 175188 331220 175240 331226
rect 175188 331162 175240 331168
rect 173728 6886 173848 6914
rect 173728 3942 173756 6886
rect 175200 3942 175228 331162
rect 176580 3942 176608 334630
rect 177948 333872 178000 333878
rect 177948 333814 178000 333820
rect 177856 330472 177908 330478
rect 177856 330414 177908 330420
rect 173164 3936 173216 3942
rect 173164 3878 173216 3884
rect 173716 3936 173768 3942
rect 173716 3878 173768 3884
rect 174268 3936 174320 3942
rect 174268 3878 174320 3884
rect 175188 3936 175240 3942
rect 175188 3878 175240 3884
rect 175464 3936 175516 3942
rect 175464 3878 175516 3884
rect 176568 3936 176620 3942
rect 176568 3878 176620 3884
rect 176660 3936 176712 3942
rect 176660 3878 176712 3884
rect 171784 2916 171836 2922
rect 171784 2858 171836 2864
rect 171968 2916 172020 2922
rect 171968 2858 172020 2864
rect 171980 480 172008 2858
rect 173176 480 173204 3878
rect 174280 480 174308 3878
rect 175476 480 175504 3878
rect 176672 480 176700 3878
rect 177868 480 177896 330414
rect 177960 3942 177988 333814
rect 177948 3936 178000 3942
rect 177948 3878 178000 3884
rect 178696 2990 178724 335718
rect 180064 335708 180116 335714
rect 180064 335650 180116 335656
rect 179328 334824 179380 334830
rect 179328 334766 179380 334772
rect 179340 6914 179368 334766
rect 179064 6886 179368 6914
rect 178684 2984 178736 2990
rect 178684 2926 178736 2932
rect 179064 480 179092 6886
rect 180076 2854 180104 335650
rect 231124 335640 231176 335646
rect 231124 335582 231176 335588
rect 201408 335300 201460 335306
rect 201408 335242 201460 335248
rect 197268 335164 197320 335170
rect 197268 335106 197320 335112
rect 194508 335096 194560 335102
rect 194508 335038 194560 335044
rect 190368 335028 190420 335034
rect 190368 334970 190420 334976
rect 183468 334960 183520 334966
rect 183468 334902 183520 334908
rect 180708 333940 180760 333946
rect 180708 333882 180760 333888
rect 180156 325780 180208 325786
rect 180156 325722 180208 325728
rect 180168 3058 180196 325722
rect 180720 3942 180748 333882
rect 181444 5024 181496 5030
rect 181444 4966 181496 4972
rect 180248 3936 180300 3942
rect 180248 3878 180300 3884
rect 180708 3936 180760 3942
rect 180708 3878 180760 3884
rect 180156 3052 180208 3058
rect 180156 2994 180208 3000
rect 180064 2848 180116 2854
rect 180064 2790 180116 2796
rect 180260 480 180288 3878
rect 181456 480 181484 4966
rect 183480 3942 183508 334902
rect 186228 334892 186280 334898
rect 186228 334834 186280 334840
rect 184848 333192 184900 333198
rect 184848 333134 184900 333140
rect 184860 3942 184888 333134
rect 186136 331696 186188 331702
rect 186136 331638 186188 331644
rect 186148 16574 186176 331638
rect 186056 16546 186176 16574
rect 186056 3942 186084 16546
rect 186240 6914 186268 334834
rect 187608 333124 187660 333130
rect 187608 333066 187660 333072
rect 187620 6914 187648 333066
rect 188988 330404 189040 330410
rect 188988 330346 189040 330352
rect 186148 6886 186268 6914
rect 187344 6886 187648 6914
rect 182548 3936 182600 3942
rect 182548 3878 182600 3884
rect 183468 3936 183520 3942
rect 183468 3878 183520 3884
rect 183744 3936 183796 3942
rect 183744 3878 183796 3884
rect 184848 3936 184900 3942
rect 184848 3878 184900 3884
rect 184940 3936 184992 3942
rect 184940 3878 184992 3884
rect 186044 3936 186096 3942
rect 186044 3878 186096 3884
rect 182560 480 182588 3878
rect 183756 480 183784 3878
rect 184952 480 184980 3878
rect 186148 480 186176 6886
rect 187344 480 187372 6886
rect 189000 3942 189028 330346
rect 190380 3942 190408 334970
rect 191748 333056 191800 333062
rect 191748 332998 191800 333004
rect 191760 3942 191788 332998
rect 194416 332988 194468 332994
rect 194416 332930 194468 332936
rect 193128 330336 193180 330342
rect 193128 330278 193180 330284
rect 193140 3942 193168 330278
rect 188528 3936 188580 3942
rect 188528 3878 188580 3884
rect 188988 3936 189040 3942
rect 188988 3878 189040 3884
rect 189724 3936 189776 3942
rect 189724 3878 189776 3884
rect 190368 3936 190420 3942
rect 190368 3878 190420 3884
rect 190828 3936 190880 3942
rect 190828 3878 190880 3884
rect 191748 3936 191800 3942
rect 191748 3878 191800 3884
rect 192024 3936 192076 3942
rect 192024 3878 192076 3884
rect 193128 3936 193180 3942
rect 193128 3878 193180 3884
rect 193220 3936 193272 3942
rect 193220 3878 193272 3884
rect 188540 480 188568 3878
rect 189736 480 189764 3878
rect 190840 480 190868 3878
rect 192036 480 192064 3878
rect 193232 480 193260 3878
rect 194428 480 194456 332930
rect 194520 3942 194548 335038
rect 195888 327548 195940 327554
rect 195888 327490 195940 327496
rect 195900 6914 195928 327490
rect 195624 6886 195928 6914
rect 194508 3936 194560 3942
rect 194508 3878 194560 3884
rect 195624 480 195652 6886
rect 197280 3942 197308 335106
rect 200028 331628 200080 331634
rect 200028 331570 200080 331576
rect 200040 3942 200068 331570
rect 201420 3942 201448 335242
rect 208308 335232 208360 335238
rect 208308 335174 208360 335180
rect 204168 334552 204220 334558
rect 204168 334494 204220 334500
rect 202788 332920 202840 332926
rect 202788 332862 202840 332868
rect 202696 330268 202748 330274
rect 202696 330210 202748 330216
rect 196808 3936 196860 3942
rect 196808 3878 196860 3884
rect 197268 3936 197320 3942
rect 197268 3878 197320 3884
rect 199108 3936 199160 3942
rect 199108 3878 199160 3884
rect 200028 3936 200080 3942
rect 200028 3878 200080 3884
rect 200304 3936 200356 3942
rect 200304 3878 200356 3884
rect 201408 3936 201460 3942
rect 201408 3878 201460 3884
rect 201500 3936 201552 3942
rect 201500 3878 201552 3884
rect 196820 480 196848 3878
rect 197912 3052 197964 3058
rect 197912 2994 197964 3000
rect 197924 480 197952 2994
rect 199120 480 199148 3878
rect 200316 480 200344 3878
rect 201512 480 201540 3878
rect 202708 480 202736 330210
rect 202800 3942 202828 332862
rect 204180 6914 204208 334494
rect 205548 332852 205600 332858
rect 205548 332794 205600 332800
rect 203904 6886 204208 6914
rect 202788 3936 202840 3942
rect 202788 3878 202840 3884
rect 203904 480 203932 6886
rect 205560 3942 205588 332794
rect 206928 330200 206980 330206
rect 206928 330142 206980 330148
rect 206940 3942 206968 330142
rect 208320 3942 208348 335174
rect 210976 334484 211028 334490
rect 210976 334426 211028 334432
rect 209780 5092 209832 5098
rect 209780 5034 209832 5040
rect 205088 3936 205140 3942
rect 205088 3878 205140 3884
rect 205548 3936 205600 3942
rect 205548 3878 205600 3884
rect 206192 3936 206244 3942
rect 206192 3878 206244 3884
rect 206928 3936 206980 3942
rect 206928 3878 206980 3884
rect 207388 3936 207440 3942
rect 207388 3878 207440 3884
rect 208308 3936 208360 3942
rect 208308 3878 208360 3884
rect 205100 480 205128 3878
rect 206204 480 206232 3878
rect 207400 480 207428 3878
rect 208584 3052 208636 3058
rect 208584 2994 208636 3000
rect 208596 480 208624 2994
rect 209792 480 209820 5034
rect 210988 480 211016 334426
rect 215208 334416 215260 334422
rect 215208 334358 215260 334364
rect 212448 331560 212500 331566
rect 212448 331502 212500 331508
rect 212460 6914 212488 331502
rect 213828 330132 213880 330138
rect 213828 330074 213880 330080
rect 212184 6886 212488 6914
rect 212184 480 212212 6886
rect 213840 3670 213868 330074
rect 215220 3670 215248 334358
rect 222108 334348 222160 334354
rect 222108 334290 222160 334296
rect 219348 334144 219400 334150
rect 219348 334086 219400 334092
rect 216588 332784 216640 332790
rect 216588 332726 216640 332732
rect 215944 327412 215996 327418
rect 215944 327354 215996 327360
rect 213368 3664 213420 3670
rect 213368 3606 213420 3612
rect 213828 3664 213880 3670
rect 213828 3606 213880 3612
rect 214472 3664 214524 3670
rect 214472 3606 214524 3612
rect 215208 3664 215260 3670
rect 215208 3606 215260 3612
rect 215668 3664 215720 3670
rect 215668 3606 215720 3612
rect 213380 480 213408 3606
rect 214484 480 214512 3606
rect 215680 480 215708 3606
rect 215956 2990 215984 327354
rect 216600 3670 216628 332726
rect 219256 332716 219308 332722
rect 219256 332658 219308 332664
rect 217968 331492 218020 331498
rect 217968 331434 218020 331440
rect 217980 3670 218008 331434
rect 216588 3664 216640 3670
rect 216588 3606 216640 3612
rect 216864 3664 216916 3670
rect 216864 3606 216916 3612
rect 217968 3664 218020 3670
rect 217968 3606 218020 3612
rect 218060 3664 218112 3670
rect 218060 3606 218112 3612
rect 215944 2984 215996 2990
rect 215944 2926 215996 2932
rect 216876 480 216904 3606
rect 218072 480 218100 3606
rect 219268 480 219296 332658
rect 219360 3670 219388 334086
rect 220728 330064 220780 330070
rect 220728 330006 220780 330012
rect 220740 6914 220768 330006
rect 220464 6886 220768 6914
rect 219348 3664 219400 3670
rect 219348 3606 219400 3612
rect 220464 480 220492 6886
rect 222120 3670 222148 334290
rect 226248 334280 226300 334286
rect 226248 334222 226300 334228
rect 223488 331424 223540 331430
rect 223488 331366 223540 331372
rect 223500 3670 223528 331366
rect 224868 329996 224920 330002
rect 224868 329938 224920 329944
rect 224880 3670 224908 329938
rect 226260 3670 226288 334222
rect 229008 334212 229060 334218
rect 229008 334154 229060 334160
rect 227628 331356 227680 331362
rect 227628 331298 227680 331304
rect 227536 329928 227588 329934
rect 227536 329870 227588 329876
rect 221556 3664 221608 3670
rect 221556 3606 221608 3612
rect 222108 3664 222160 3670
rect 222108 3606 222160 3612
rect 222752 3664 222804 3670
rect 222752 3606 222804 3612
rect 223488 3664 223540 3670
rect 223488 3606 223540 3612
rect 223948 3664 224000 3670
rect 223948 3606 224000 3612
rect 224868 3664 224920 3670
rect 224868 3606 224920 3612
rect 225144 3664 225196 3670
rect 225144 3606 225196 3612
rect 226248 3664 226300 3670
rect 226248 3606 226300 3612
rect 226340 3664 226392 3670
rect 226340 3606 226392 3612
rect 221568 480 221596 3606
rect 222764 480 222792 3606
rect 223960 480 223988 3606
rect 225156 480 225184 3606
rect 226352 480 226380 3606
rect 227548 480 227576 329870
rect 227640 3670 227668 331298
rect 229020 6914 229048 334154
rect 230388 332036 230440 332042
rect 230388 331978 230440 331984
rect 228744 6886 229048 6914
rect 227628 3664 227680 3670
rect 227628 3606 227680 3612
rect 228744 480 228772 6886
rect 230400 3534 230428 331978
rect 231136 3602 231164 335582
rect 231216 335436 231268 335442
rect 231216 335378 231268 335384
rect 231228 3670 231256 335378
rect 231306 334112 231362 334121
rect 231306 334047 231362 334056
rect 231400 334076 231452 334082
rect 231216 3664 231268 3670
rect 231216 3606 231268 3612
rect 231124 3596 231176 3602
rect 231124 3538 231176 3544
rect 229836 3528 229888 3534
rect 229836 3470 229888 3476
rect 230388 3528 230440 3534
rect 230388 3470 230440 3476
rect 231032 3528 231084 3534
rect 231032 3470 231084 3476
rect 229848 480 229876 3470
rect 231044 480 231072 3470
rect 231320 3466 231348 334047
rect 231400 334018 231452 334024
rect 231308 3460 231360 3466
rect 231308 3402 231360 3408
rect 231412 2922 231440 334018
rect 231768 327480 231820 327486
rect 231768 327422 231820 327428
rect 231780 3534 231808 327422
rect 232056 248402 232084 342751
rect 232148 338638 232176 349794
rect 232136 338632 232188 338638
rect 232136 338574 232188 338580
rect 232240 321842 232268 352407
rect 232332 337550 232360 358119
rect 232410 356280 232466 356289
rect 232410 356215 232466 356224
rect 232320 337544 232372 337550
rect 232320 337486 232372 337492
rect 232228 321836 232280 321842
rect 232228 321778 232280 321784
rect 232424 321774 232452 356215
rect 232516 337346 232544 363967
rect 232504 337340 232556 337346
rect 232504 337282 232556 337288
rect 232504 334008 232556 334014
rect 232504 333950 232556 333956
rect 232412 321768 232464 321774
rect 232412 321710 232464 321716
rect 232044 248396 232096 248402
rect 232044 248338 232096 248344
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 231400 2916 231452 2922
rect 231400 2858 231452 2864
rect 232240 480 232268 3470
rect 232516 3126 232544 333950
rect 232608 322726 232636 373487
rect 232700 322794 232728 379335
rect 232688 322788 232740 322794
rect 232688 322730 232740 322736
rect 232596 322720 232648 322726
rect 232596 322662 232648 322668
rect 232792 321910 232820 385047
rect 232870 381304 232926 381313
rect 232870 381239 232926 381248
rect 232884 349858 232912 381239
rect 233054 377496 233110 377505
rect 233054 377431 233110 377440
rect 232962 375456 233018 375465
rect 232962 375391 233018 375400
rect 232872 349852 232924 349858
rect 232872 349794 232924 349800
rect 232870 346624 232926 346633
rect 232870 346559 232926 346568
rect 232884 338570 232912 346559
rect 232872 338564 232924 338570
rect 232872 338506 232924 338512
rect 232872 335504 232924 335510
rect 232872 335446 232924 335452
rect 232884 331974 232912 335446
rect 232872 331968 232924 331974
rect 232872 331910 232924 331916
rect 232780 321904 232832 321910
rect 232780 321846 232832 321852
rect 232976 238950 233004 375391
rect 232964 238944 233016 238950
rect 232964 238886 233016 238892
rect 233068 238882 233096 377431
rect 233160 322402 233188 386951
rect 234434 383208 234490 383217
rect 234434 383143 234490 383152
rect 234342 371648 234398 371657
rect 234342 371583 234398 371592
rect 234158 369744 234214 369753
rect 234158 369679 234214 369688
rect 234066 365936 234122 365945
rect 234066 365871 234122 365880
rect 233974 361992 234030 362001
rect 233974 361927 234030 361936
rect 233882 360088 233938 360097
rect 233882 360023 233938 360032
rect 233790 354376 233846 354385
rect 233790 354311 233846 354320
rect 233698 350432 233754 350441
rect 233698 350367 233754 350376
rect 233514 344720 233570 344729
rect 233514 344655 233570 344664
rect 233238 338056 233294 338065
rect 233238 337991 233294 338000
rect 233252 329458 233280 337991
rect 233330 337920 233386 337929
rect 233330 337855 233386 337864
rect 233344 330449 233372 337855
rect 233528 337414 233556 344655
rect 233606 340912 233662 340921
rect 233606 340847 233662 340856
rect 233620 338026 233648 340847
rect 233608 338020 233660 338026
rect 233608 337962 233660 337968
rect 233516 337408 233568 337414
rect 233516 337350 233568 337356
rect 233608 336048 233660 336054
rect 233608 335990 233660 335996
rect 233620 331294 233648 335990
rect 233608 331288 233660 331294
rect 233608 331230 233660 331236
rect 233330 330440 233386 330449
rect 233330 330375 233386 330384
rect 233240 329452 233292 329458
rect 233240 329394 233292 329400
rect 233160 322374 233280 322402
rect 233148 322244 233200 322250
rect 233148 322186 233200 322192
rect 233056 238876 233108 238882
rect 233056 238818 233108 238824
rect 233160 3534 233188 322186
rect 233252 321978 233280 322374
rect 233240 321972 233292 321978
rect 233240 321914 233292 321920
rect 233712 237318 233740 350367
rect 233804 237386 233832 354311
rect 233896 238377 233924 360023
rect 233882 238368 233938 238377
rect 233882 238303 233938 238312
rect 233792 237380 233844 237386
rect 233792 237322 233844 237328
rect 233700 237312 233752 237318
rect 233700 237254 233752 237260
rect 233988 237153 234016 361927
rect 234080 238513 234108 365871
rect 234172 238649 234200 369679
rect 234250 367840 234306 367849
rect 234250 367775 234306 367784
rect 234158 238640 234214 238649
rect 234158 238575 234214 238584
rect 234066 238504 234122 238513
rect 234066 238439 234122 238448
rect 233974 237144 234030 237153
rect 233974 237079 234030 237088
rect 234264 237017 234292 367775
rect 234250 237008 234306 237017
rect 234250 236943 234306 236952
rect 234356 236473 234384 371583
rect 234448 238814 234476 383143
rect 285140 373994 285168 390118
rect 285048 373966 285168 373994
rect 234526 348528 234582 348537
rect 234526 348463 234582 348472
rect 234540 338706 234568 348463
rect 234710 339008 234766 339017
rect 234710 338943 234766 338952
rect 234528 338700 234580 338706
rect 234528 338642 234580 338648
rect 234620 338088 234672 338094
rect 234620 338030 234672 338036
rect 234632 336161 234660 338030
rect 234724 337482 234752 338943
rect 234816 338014 235060 338042
rect 234712 337476 234764 337482
rect 234712 337418 234764 337424
rect 234618 336152 234674 336161
rect 234618 336087 234674 336096
rect 234632 333577 234660 336087
rect 234618 333568 234674 333577
rect 234618 333503 234674 333512
rect 234816 333441 234844 338014
rect 234896 337952 234948 337958
rect 234896 337894 234948 337900
rect 234802 333432 234858 333441
rect 234802 333367 234858 333376
rect 234528 332648 234580 332654
rect 234528 332590 234580 332596
rect 234436 238808 234488 238814
rect 234436 238750 234488 238756
rect 234342 236464 234398 236473
rect 234342 236399 234398 236408
rect 234540 3534 234568 332590
rect 234712 331968 234764 331974
rect 234712 331910 234764 331916
rect 234724 326398 234752 331910
rect 234908 327826 234936 337894
rect 235138 337872 235166 338028
rect 235092 337844 235166 337872
rect 234988 337544 235040 337550
rect 234988 337486 235040 337492
rect 235000 336297 235028 337486
rect 234986 336288 235042 336297
rect 234986 336223 235042 336232
rect 234988 335436 235040 335442
rect 234988 335378 235040 335384
rect 234896 327820 234948 327826
rect 234896 327762 234948 327768
rect 235000 326398 235028 335378
rect 235092 331809 235120 337844
rect 235230 337770 235258 338028
rect 235322 337958 235350 338028
rect 235310 337952 235362 337958
rect 235310 337894 235362 337900
rect 235414 337804 235442 338028
rect 235506 337890 235534 338028
rect 235598 337958 235626 338028
rect 235586 337952 235638 337958
rect 235586 337894 235638 337900
rect 235494 337884 235546 337890
rect 235494 337826 235546 337832
rect 235690 337822 235718 338028
rect 235184 337742 235258 337770
rect 235368 337776 235442 337804
rect 235678 337816 235730 337822
rect 235538 337784 235594 337793
rect 235184 331945 235212 337742
rect 235368 337634 235396 337776
rect 235678 337758 235730 337764
rect 235782 337770 235810 338028
rect 235874 337890 235902 338028
rect 235862 337884 235914 337890
rect 235862 337826 235914 337832
rect 235966 337770 235994 338028
rect 235782 337742 235856 337770
rect 235538 337719 235594 337728
rect 235276 337606 235396 337634
rect 235448 337612 235500 337618
rect 235170 331936 235226 331945
rect 235170 331871 235226 331880
rect 235078 331800 235134 331809
rect 235276 331786 235304 337606
rect 235448 337554 235500 337560
rect 235460 332081 235488 337554
rect 235552 335889 235580 337719
rect 235632 337612 235684 337618
rect 235632 337554 235684 337560
rect 235538 335880 235594 335889
rect 235538 335815 235594 335824
rect 235446 332072 235502 332081
rect 235446 332007 235502 332016
rect 235078 331735 235134 331744
rect 235184 331758 235304 331786
rect 235184 328454 235212 331758
rect 235264 329860 235316 329866
rect 235264 329802 235316 329808
rect 235092 328426 235212 328454
rect 234712 326392 234764 326398
rect 234712 326334 234764 326340
rect 234988 326392 235040 326398
rect 234988 326334 235040 326340
rect 235092 324970 235120 328426
rect 235080 324964 235132 324970
rect 235080 324906 235132 324912
rect 234620 5160 234672 5166
rect 234620 5102 234672 5108
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233424 3528 233476 3534
rect 233424 3470 233476 3476
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 232504 3120 232556 3126
rect 232504 3062 232556 3068
rect 233436 480 233464 3470
rect 234632 480 234660 5102
rect 235276 3398 235304 329802
rect 235644 327758 235672 337554
rect 235828 331974 235856 337742
rect 235920 337742 235994 337770
rect 235816 331968 235868 331974
rect 235816 331910 235868 331916
rect 235920 329118 235948 337742
rect 236058 337634 236086 338028
rect 236012 337606 236086 337634
rect 236012 329186 236040 337606
rect 236150 337532 236178 338028
rect 236242 337770 236270 338028
rect 236334 337958 236362 338028
rect 236322 337952 236374 337958
rect 236426 337929 236454 338028
rect 236322 337894 236374 337900
rect 236412 337920 236468 337929
rect 236412 337855 236468 337864
rect 236518 337822 236546 338028
rect 236610 337822 236638 338028
rect 236506 337816 236558 337822
rect 236242 337742 236408 337770
rect 236506 337758 236558 337764
rect 236598 337816 236650 337822
rect 236702 337804 236730 338028
rect 236794 338008 236822 338028
rect 236932 338014 236992 338042
rect 236794 337980 236868 338008
rect 236702 337776 236776 337804
rect 236598 337758 236650 337764
rect 236104 337504 236178 337532
rect 236104 336025 236132 337504
rect 236184 337272 236236 337278
rect 236184 337214 236236 337220
rect 236090 336016 236146 336025
rect 236090 335951 236146 335960
rect 236196 335753 236224 337214
rect 236182 335744 236238 335753
rect 236182 335679 236238 335688
rect 236196 334665 236224 335679
rect 236380 335617 236408 337742
rect 236748 336025 236776 337776
rect 236734 336016 236790 336025
rect 236734 335951 236790 335960
rect 236366 335608 236422 335617
rect 236366 335543 236422 335552
rect 236182 334656 236238 334665
rect 236182 334591 236238 334600
rect 236748 334121 236776 335951
rect 236840 335646 236868 337980
rect 236932 336122 236960 338014
rect 237070 337940 237098 338028
rect 237162 337958 237190 338028
rect 237024 337912 237098 337940
rect 237150 337952 237202 337958
rect 236920 336116 236972 336122
rect 236920 336058 236972 336064
rect 237024 336002 237052 337912
rect 237150 337894 237202 337900
rect 237254 337770 237282 338028
rect 237346 337890 237374 338028
rect 237334 337884 237386 337890
rect 237334 337826 237386 337832
rect 237438 337770 237466 338028
rect 237530 337822 237558 338028
rect 236932 335974 237052 336002
rect 237208 337742 237282 337770
rect 237392 337742 237466 337770
rect 237518 337816 237570 337822
rect 237518 337758 237570 337764
rect 237622 337770 237650 338028
rect 237714 337958 237742 338028
rect 237702 337952 237754 337958
rect 237702 337894 237754 337900
rect 237806 337770 237834 338028
rect 237898 337958 237926 338028
rect 237886 337952 237938 337958
rect 237886 337894 237938 337900
rect 237990 337770 238018 338028
rect 238082 337890 238110 338028
rect 238070 337884 238122 337890
rect 238070 337826 238122 337832
rect 238174 337770 238202 338028
rect 237622 337742 237696 337770
rect 236828 335640 236880 335646
rect 236828 335582 236880 335588
rect 236826 335472 236882 335481
rect 236932 335458 236960 335974
rect 236882 335430 236960 335458
rect 236826 335407 236882 335416
rect 236734 334112 236790 334121
rect 236734 334047 236790 334056
rect 236366 333840 236422 333849
rect 236366 333775 236422 333784
rect 236642 333840 236698 333849
rect 236642 333775 236698 333784
rect 236380 333577 236408 333775
rect 236366 333568 236422 333577
rect 236366 333503 236422 333512
rect 236460 331968 236512 331974
rect 236460 331910 236512 331916
rect 236000 329180 236052 329186
rect 236000 329122 236052 329128
rect 235908 329112 235960 329118
rect 235908 329054 235960 329060
rect 235632 327752 235684 327758
rect 235632 327694 235684 327700
rect 236472 327418 236500 331910
rect 236460 327412 236512 327418
rect 236460 327354 236512 327360
rect 235356 326392 235408 326398
rect 235356 326334 235408 326340
rect 235368 325718 235396 326334
rect 235356 325712 235408 325718
rect 235356 325654 235408 325660
rect 235368 238921 235396 325654
rect 235354 238912 235410 238921
rect 235354 238847 235410 238856
rect 235816 3868 235868 3874
rect 235816 3810 235868 3816
rect 235264 3392 235316 3398
rect 235264 3334 235316 3340
rect 235828 480 235856 3810
rect 236656 2990 236684 333775
rect 236932 333169 236960 335430
rect 237010 335472 237066 335481
rect 237010 335407 237066 335416
rect 237024 333305 237052 335407
rect 237010 333296 237066 333305
rect 237010 333231 237066 333240
rect 236918 333160 236974 333169
rect 236918 333095 236974 333104
rect 237208 327962 237236 337742
rect 237392 336870 237420 337742
rect 237564 337272 237616 337278
rect 237564 337214 237616 337220
rect 237380 336864 237432 336870
rect 237380 336806 237432 336812
rect 237392 335481 237420 336806
rect 237378 335472 237434 335481
rect 237378 335407 237434 335416
rect 237470 333432 237526 333441
rect 237470 333367 237526 333376
rect 237288 331356 237340 331362
rect 237288 331298 237340 331304
rect 237196 327956 237248 327962
rect 237196 327898 237248 327904
rect 237300 326398 237328 331298
rect 237484 329254 237512 333367
rect 237472 329248 237524 329254
rect 237472 329190 237524 329196
rect 237576 326466 237604 337214
rect 237668 336433 237696 337742
rect 237760 337742 237834 337770
rect 237944 337742 238018 337770
rect 238128 337742 238202 337770
rect 238266 337770 238294 338028
rect 238358 337890 238386 338028
rect 238450 337890 238478 338028
rect 238542 337929 238570 338028
rect 238634 337958 238662 338028
rect 238726 337958 238754 338028
rect 238910 337958 238938 338028
rect 238622 337952 238674 337958
rect 238528 337920 238584 337929
rect 238346 337884 238398 337890
rect 238346 337826 238398 337832
rect 238438 337884 238490 337890
rect 238622 337894 238674 337900
rect 238714 337952 238766 337958
rect 238714 337894 238766 337900
rect 238898 337952 238950 337958
rect 238898 337894 238950 337900
rect 238528 337855 238584 337864
rect 238438 337826 238490 337832
rect 238668 337816 238720 337822
rect 238266 337742 238340 337770
rect 238668 337758 238720 337764
rect 238760 337816 238812 337822
rect 239002 337770 239030 338028
rect 239094 337822 239122 338028
rect 238760 337758 238812 337764
rect 237654 336424 237710 336433
rect 237654 336359 237710 336368
rect 237760 326534 237788 337742
rect 237840 337612 237892 337618
rect 237840 337554 237892 337560
rect 237852 336938 237880 337554
rect 237840 336932 237892 336938
rect 237840 336874 237892 336880
rect 237852 336258 237880 336874
rect 237840 336252 237892 336258
rect 237840 336194 237892 336200
rect 237944 336138 237972 337742
rect 238024 337612 238076 337618
rect 238024 337554 238076 337560
rect 238036 336569 238064 337554
rect 238022 336560 238078 336569
rect 238022 336495 238078 336504
rect 238128 336190 238156 337742
rect 237852 336110 237972 336138
rect 238116 336184 238168 336190
rect 238116 336126 238168 336132
rect 238208 336184 238260 336190
rect 238208 336126 238260 336132
rect 237852 334121 237880 336110
rect 237932 335504 237984 335510
rect 237932 335446 237984 335452
rect 237838 334112 237894 334121
rect 237838 334047 237894 334056
rect 237852 331906 237880 334047
rect 237944 333577 237972 335446
rect 238024 335368 238076 335374
rect 238024 335310 238076 335316
rect 237930 333568 237986 333577
rect 237930 333503 237986 333512
rect 237840 331900 237892 331906
rect 237840 331842 237892 331848
rect 237748 326528 237800 326534
rect 237748 326470 237800 326476
rect 237564 326460 237616 326466
rect 237564 326402 237616 326408
rect 236736 326392 236788 326398
rect 236736 326334 236788 326340
rect 237288 326392 237340 326398
rect 237288 326334 237340 326340
rect 236748 325786 236776 326334
rect 236736 325780 236788 325786
rect 236736 325722 236788 325728
rect 236748 238785 236776 325722
rect 236734 238776 236790 238785
rect 236734 238711 236790 238720
rect 238036 3738 238064 335310
rect 238220 333713 238248 336126
rect 238206 333704 238262 333713
rect 238206 333639 238262 333648
rect 238312 333441 238340 337742
rect 238576 337612 238628 337618
rect 238576 337554 238628 337560
rect 238298 333432 238354 333441
rect 238298 333367 238354 333376
rect 238312 332625 238340 333367
rect 238298 332616 238354 332625
rect 238298 332551 238354 332560
rect 238116 331968 238168 331974
rect 238116 331910 238168 331916
rect 238024 3732 238076 3738
rect 238024 3674 238076 3680
rect 238128 3670 238156 331910
rect 238588 13122 238616 337554
rect 238680 326874 238708 337758
rect 238772 336705 238800 337758
rect 238956 337742 239030 337770
rect 239082 337816 239134 337822
rect 239082 337758 239134 337764
rect 238758 336696 238814 336705
rect 238758 336631 238814 336640
rect 238852 336388 238904 336394
rect 238852 336330 238904 336336
rect 238760 336116 238812 336122
rect 238760 336058 238812 336064
rect 238772 334626 238800 336058
rect 238760 334620 238812 334626
rect 238760 334562 238812 334568
rect 238864 328030 238892 336330
rect 238956 335628 238984 337742
rect 239186 337634 239214 338028
rect 239278 337958 239306 338028
rect 239370 337958 239398 338028
rect 239266 337952 239318 337958
rect 239266 337894 239318 337900
rect 239358 337952 239410 337958
rect 239462 337929 239490 338028
rect 239554 337958 239582 338028
rect 239542 337952 239594 337958
rect 239358 337894 239410 337900
rect 239448 337920 239504 337929
rect 239646 337929 239674 338028
rect 239738 337958 239766 338028
rect 239726 337952 239778 337958
rect 239542 337894 239594 337900
rect 239632 337920 239688 337929
rect 239448 337855 239504 337864
rect 239830 337929 239858 338028
rect 239726 337894 239778 337900
rect 239816 337920 239872 337929
rect 239632 337855 239688 337864
rect 239922 337890 239950 338028
rect 239816 337855 239872 337864
rect 239910 337884 239962 337890
rect 239910 337826 239962 337832
rect 239772 337816 239824 337822
rect 239772 337758 239824 337764
rect 239862 337784 239918 337793
rect 239140 337606 239214 337634
rect 239494 337648 239550 337657
rect 239312 337612 239364 337618
rect 239140 337532 239168 337606
rect 239494 337583 239550 337592
rect 239312 337554 239364 337560
rect 239140 337504 239260 337532
rect 239128 335912 239180 335918
rect 239048 335860 239128 335866
rect 239048 335854 239180 335860
rect 239048 335838 239168 335854
rect 239048 335782 239076 335838
rect 239036 335776 239088 335782
rect 239036 335718 239088 335724
rect 238956 335600 239076 335628
rect 238944 331356 238996 331362
rect 238944 331298 238996 331304
rect 238956 328098 238984 331298
rect 239048 329390 239076 335600
rect 239128 334144 239180 334150
rect 239128 334086 239180 334092
rect 239036 329384 239088 329390
rect 239036 329326 239088 329332
rect 238944 328092 238996 328098
rect 238944 328034 238996 328040
rect 238852 328024 238904 328030
rect 238852 327966 238904 327972
rect 238668 326868 238720 326874
rect 238668 326810 238720 326816
rect 239140 326602 239168 334086
rect 239232 332217 239260 337504
rect 239218 332208 239274 332217
rect 239218 332143 239274 332152
rect 239324 327894 239352 337554
rect 239404 331968 239456 331974
rect 239404 331910 239456 331916
rect 239312 327888 239364 327894
rect 239312 327830 239364 327836
rect 239128 326596 239180 326602
rect 239128 326538 239180 326544
rect 238576 13116 238628 13122
rect 238576 13058 238628 13064
rect 239416 3806 239444 331910
rect 239508 331838 239536 337583
rect 239496 331832 239548 331838
rect 239496 331774 239548 331780
rect 239784 330585 239812 337758
rect 240014 337770 240042 338028
rect 239862 337719 239918 337728
rect 239968 337742 240042 337770
rect 239876 331362 239904 337719
rect 239864 331356 239916 331362
rect 239864 331298 239916 331304
rect 239968 330721 239996 337742
rect 240106 337634 240134 338028
rect 240198 337770 240226 338028
rect 240290 337890 240318 338028
rect 240278 337884 240330 337890
rect 240278 337826 240330 337832
rect 240382 337770 240410 338028
rect 240198 337742 240272 337770
rect 240060 337606 240134 337634
rect 240060 334150 240088 337606
rect 240140 336728 240192 336734
rect 240140 336670 240192 336676
rect 240152 335345 240180 336670
rect 240244 336394 240272 337742
rect 240336 337742 240410 337770
rect 240474 337770 240502 338028
rect 240566 337890 240594 338028
rect 240554 337884 240606 337890
rect 240554 337826 240606 337832
rect 240658 337770 240686 338028
rect 240474 337742 240548 337770
rect 240232 336388 240284 336394
rect 240232 336330 240284 336336
rect 240232 336252 240284 336258
rect 240232 336194 240284 336200
rect 240138 335336 240194 335345
rect 240138 335271 240194 335280
rect 240244 334762 240272 336194
rect 240232 334756 240284 334762
rect 240232 334698 240284 334704
rect 240048 334144 240100 334150
rect 240048 334086 240100 334092
rect 239954 330712 240010 330721
rect 239954 330647 240010 330656
rect 239770 330576 239826 330585
rect 239770 330511 239826 330520
rect 240336 328166 240364 337742
rect 240416 336796 240468 336802
rect 240416 336738 240468 336744
rect 240428 335578 240456 336738
rect 240416 335572 240468 335578
rect 240416 335514 240468 335520
rect 240416 334620 240468 334626
rect 240416 334562 240468 334568
rect 240428 332353 240456 334562
rect 240414 332344 240470 332353
rect 240414 332279 240470 332288
rect 240520 330970 240548 337742
rect 240428 330942 240548 330970
rect 240612 337742 240686 337770
rect 240796 338014 240856 338042
rect 240324 328160 240376 328166
rect 240324 328102 240376 328108
rect 240428 325694 240456 330942
rect 240612 328234 240640 337742
rect 240796 337498 240824 338014
rect 240934 337770 240962 338028
rect 240704 337470 240824 337498
rect 240888 337742 240962 337770
rect 241026 337770 241054 338028
rect 241118 337958 241146 338028
rect 241106 337952 241158 337958
rect 241210 337929 241238 338028
rect 241106 337894 241158 337900
rect 241196 337920 241252 337929
rect 241196 337855 241252 337864
rect 241302 337804 241330 338028
rect 241394 337958 241422 338028
rect 241382 337952 241434 337958
rect 241382 337894 241434 337900
rect 241164 337776 241330 337804
rect 241026 337742 241100 337770
rect 240704 336802 240732 337470
rect 240692 336796 240744 336802
rect 240692 336738 240744 336744
rect 240692 336456 240744 336462
rect 240692 336398 240744 336404
rect 240704 334150 240732 336398
rect 240888 334626 240916 337742
rect 240966 337648 241022 337657
rect 240966 337583 241022 337592
rect 240876 334620 240928 334626
rect 240876 334562 240928 334568
rect 240980 334506 241008 337583
rect 240888 334478 241008 334506
rect 240692 334144 240744 334150
rect 240692 334086 240744 334092
rect 240692 331356 240744 331362
rect 240692 331298 240744 331304
rect 240600 328228 240652 328234
rect 240600 328170 240652 328176
rect 240428 325666 240640 325694
rect 240612 4826 240640 325666
rect 240704 6186 240732 331298
rect 240888 328370 240916 334478
rect 240968 334144 241020 334150
rect 240968 334086 241020 334092
rect 240876 328364 240928 328370
rect 240876 328306 240928 328312
rect 240980 323610 241008 334086
rect 241072 328302 241100 337742
rect 241164 337657 241192 337776
rect 241150 337648 241206 337657
rect 241486 337634 241514 338028
rect 241578 337770 241606 338028
rect 241670 337890 241698 338028
rect 241658 337884 241710 337890
rect 241658 337826 241710 337832
rect 241762 337770 241790 338028
rect 241578 337742 241652 337770
rect 241150 337583 241206 337592
rect 241440 337606 241514 337634
rect 241152 337544 241204 337550
rect 241152 337486 241204 337492
rect 241164 330857 241192 337486
rect 241242 336016 241298 336025
rect 241242 335951 241298 335960
rect 241256 335374 241284 335951
rect 241244 335368 241296 335374
rect 241244 335310 241296 335316
rect 241244 334620 241296 334626
rect 241244 334562 241296 334568
rect 241150 330848 241206 330857
rect 241150 330783 241206 330792
rect 241256 330546 241284 334562
rect 241244 330540 241296 330546
rect 241244 330482 241296 330488
rect 241440 329526 241468 337606
rect 241624 336802 241652 337742
rect 241716 337742 241790 337770
rect 241612 336796 241664 336802
rect 241612 336738 241664 336744
rect 241716 330614 241744 337742
rect 241854 337634 241882 338028
rect 241946 337770 241974 338028
rect 242038 337895 242066 338028
rect 242024 337886 242080 337895
rect 242024 337821 242080 337830
rect 242130 337770 242158 338028
rect 242222 337929 242250 338028
rect 242208 337920 242264 337929
rect 242314 337890 242342 338028
rect 242406 337958 242434 338028
rect 242394 337952 242446 337958
rect 242394 337894 242446 337900
rect 242498 337906 242526 338028
rect 242590 338008 242618 338028
rect 242728 338026 242788 338042
rect 242716 338020 242788 338026
rect 242590 337980 242664 338008
rect 242208 337855 242264 337864
rect 242302 337884 242354 337890
rect 242498 337878 242572 337906
rect 242302 337826 242354 337832
rect 242440 337816 242492 337822
rect 241946 337742 242020 337770
rect 241808 337606 241882 337634
rect 241704 330608 241756 330614
rect 241704 330550 241756 330556
rect 241428 329520 241480 329526
rect 241428 329462 241480 329468
rect 241808 328438 241836 337606
rect 241886 337512 241942 337521
rect 241886 337447 241942 337456
rect 241900 329594 241928 337447
rect 241888 329588 241940 329594
rect 241888 329530 241940 329536
rect 241796 328432 241848 328438
rect 241796 328374 241848 328380
rect 241060 328296 241112 328302
rect 241060 328238 241112 328244
rect 240968 323604 241020 323610
rect 240968 323546 241020 323552
rect 240692 6180 240744 6186
rect 240692 6122 240744 6128
rect 240600 4820 240652 4826
rect 240600 4762 240652 4768
rect 241992 4010 242020 337742
rect 242084 337742 242158 337770
rect 242254 337784 242310 337793
rect 242084 335442 242112 337742
rect 242440 337758 242492 337764
rect 242254 337719 242310 337728
rect 242268 336054 242296 337719
rect 242256 336048 242308 336054
rect 242256 335990 242308 335996
rect 242164 335504 242216 335510
rect 242164 335446 242216 335452
rect 242072 335436 242124 335442
rect 242072 335378 242124 335384
rect 242072 334144 242124 334150
rect 242072 334086 242124 334092
rect 242084 4078 242112 334086
rect 242176 326738 242204 335446
rect 242256 335436 242308 335442
rect 242256 335378 242308 335384
rect 242268 333538 242296 335378
rect 242256 333532 242308 333538
rect 242256 333474 242308 333480
rect 242452 327690 242480 337758
rect 242544 334150 242572 337878
rect 242532 334144 242584 334150
rect 242532 334086 242584 334092
rect 242636 329730 242664 337980
rect 242768 338014 242788 338020
rect 242716 337962 242768 337968
rect 242866 337872 242894 338028
rect 242958 337929 242986 338028
rect 242820 337844 242894 337872
rect 242944 337920 243000 337929
rect 243050 337890 243078 338028
rect 243142 337958 243170 338028
rect 243130 337952 243182 337958
rect 243130 337894 243182 337900
rect 243234 337890 243262 338028
rect 242944 337855 243000 337864
rect 243038 337884 243090 337890
rect 242716 337000 242768 337006
rect 242716 336942 242768 336948
rect 242624 329724 242676 329730
rect 242624 329666 242676 329672
rect 242440 327684 242492 327690
rect 242440 327626 242492 327632
rect 242164 326732 242216 326738
rect 242164 326674 242216 326680
rect 242728 326670 242756 336942
rect 242820 336666 242848 337844
rect 243038 337826 243090 337832
rect 243222 337884 243274 337890
rect 243222 337826 243274 337832
rect 242898 337784 242954 337793
rect 242898 337719 242954 337728
rect 243174 337784 243230 337793
rect 243326 337770 243354 338028
rect 243174 337719 243230 337728
rect 243280 337742 243354 337770
rect 242808 336660 242860 336666
rect 242808 336602 242860 336608
rect 242806 336152 242862 336161
rect 242806 336087 242862 336096
rect 242820 336054 242848 336087
rect 242808 336048 242860 336054
rect 242808 335990 242860 335996
rect 242912 329798 242940 337719
rect 243188 330818 243216 337719
rect 243280 335050 243308 337742
rect 243418 337634 243446 338028
rect 243510 337770 243538 338028
rect 243602 337890 243630 338028
rect 243590 337884 243642 337890
rect 243590 337826 243642 337832
rect 243694 337770 243722 338028
rect 243786 337890 243814 338028
rect 243774 337884 243826 337890
rect 243774 337826 243826 337832
rect 243878 337770 243906 338028
rect 243510 337742 243584 337770
rect 243418 337606 243492 337634
rect 243360 337544 243412 337550
rect 243360 337486 243412 337492
rect 243372 335510 243400 337486
rect 243464 336530 243492 337606
rect 243452 336524 243504 336530
rect 243452 336466 243504 336472
rect 243452 336388 243504 336394
rect 243452 336330 243504 336336
rect 243360 335504 243412 335510
rect 243360 335446 243412 335452
rect 243280 335022 243400 335050
rect 243268 334960 243320 334966
rect 243268 334902 243320 334908
rect 243176 330812 243228 330818
rect 243176 330754 243228 330760
rect 242900 329792 242952 329798
rect 242900 329734 242952 329740
rect 243280 326942 243308 334902
rect 243372 333849 243400 335022
rect 243358 333840 243414 333849
rect 243358 333775 243414 333784
rect 243464 327010 243492 336330
rect 243556 334626 243584 337742
rect 243648 337742 243722 337770
rect 243832 337742 243906 337770
rect 243970 337770 243998 338028
rect 244062 337895 244090 338028
rect 244048 337886 244104 337895
rect 244048 337821 244104 337830
rect 244154 337770 244182 338028
rect 244246 337890 244274 338028
rect 244234 337884 244286 337890
rect 244234 337826 244286 337832
rect 244338 337770 244366 338028
rect 244430 337872 244458 338028
rect 244522 338008 244550 338028
rect 244522 337980 244596 338008
rect 244568 337890 244596 337980
rect 244556 337884 244608 337890
rect 244430 337844 244504 337872
rect 243970 337742 244044 337770
rect 244154 337742 244228 337770
rect 244338 337742 244412 337770
rect 243544 334620 243596 334626
rect 243544 334562 243596 334568
rect 243452 327004 243504 327010
rect 243452 326946 243504 326952
rect 243268 326936 243320 326942
rect 243268 326878 243320 326884
rect 243648 326806 243676 337742
rect 243726 337512 243782 337521
rect 243726 337447 243782 337456
rect 243740 336190 243768 337447
rect 243728 336184 243780 336190
rect 243728 336126 243780 336132
rect 243832 335646 243860 337742
rect 244016 337668 244044 337742
rect 243924 337640 244044 337668
rect 244094 337648 244150 337657
rect 243924 336938 243952 337640
rect 244094 337583 244150 337592
rect 244004 337544 244056 337550
rect 244004 337486 244056 337492
rect 243912 336932 243964 336938
rect 243912 336874 243964 336880
rect 243820 335640 243872 335646
rect 243820 335582 243872 335588
rect 244016 334966 244044 337486
rect 244004 334960 244056 334966
rect 244004 334902 244056 334908
rect 243728 334620 243780 334626
rect 243728 334562 243780 334568
rect 243740 329050 243768 334562
rect 243820 334144 243872 334150
rect 243820 334086 243872 334092
rect 243728 329044 243780 329050
rect 243728 328986 243780 328992
rect 243832 327622 243860 334086
rect 244108 328914 244136 337583
rect 244200 336462 244228 337742
rect 244188 336456 244240 336462
rect 244188 336398 244240 336404
rect 244188 335504 244240 335510
rect 244188 335446 244240 335452
rect 244200 335306 244228 335446
rect 244188 335300 244240 335306
rect 244188 335242 244240 335248
rect 244096 328908 244148 328914
rect 244096 328850 244148 328856
rect 244384 328846 244412 337742
rect 244476 335986 244504 337844
rect 244556 337826 244608 337832
rect 244554 337784 244610 337793
rect 244554 337719 244610 337728
rect 244464 335980 244516 335986
rect 244464 335922 244516 335928
rect 244464 335436 244516 335442
rect 244464 335378 244516 335384
rect 244476 334558 244504 335378
rect 244568 335073 244596 337719
rect 244706 337668 244734 338028
rect 244798 337770 244826 338028
rect 244890 337929 244918 338028
rect 244876 337920 244932 337929
rect 244876 337855 244932 337864
rect 244982 337822 245010 338028
rect 245074 337890 245102 338028
rect 245062 337884 245114 337890
rect 245062 337826 245114 337832
rect 244970 337816 245022 337822
rect 244798 337742 244872 337770
rect 245166 337770 245194 338028
rect 244970 337758 245022 337764
rect 244706 337640 244780 337668
rect 244554 335064 244610 335073
rect 244554 334999 244610 335008
rect 244648 334620 244700 334626
rect 244648 334562 244700 334568
rect 244464 334552 244516 334558
rect 244464 334494 244516 334500
rect 244372 328840 244424 328846
rect 244372 328782 244424 328788
rect 243820 327616 243872 327622
rect 243820 327558 243872 327564
rect 243636 326800 243688 326806
rect 243636 326742 243688 326748
rect 242716 326664 242768 326670
rect 242716 326606 242768 326612
rect 242072 4072 242124 4078
rect 242072 4014 242124 4020
rect 241980 4004 242032 4010
rect 241980 3946 242032 3952
rect 239404 3800 239456 3806
rect 239404 3742 239456 3748
rect 241704 3800 241756 3806
rect 241704 3742 241756 3748
rect 238116 3664 238168 3670
rect 238116 3606 238168 3612
rect 240508 3664 240560 3670
rect 240508 3606 240560 3612
rect 239312 3596 239364 3602
rect 239312 3538 239364 3544
rect 237012 3528 237064 3534
rect 237012 3470 237064 3476
rect 236644 2984 236696 2990
rect 236644 2926 236696 2932
rect 237024 480 237052 3470
rect 238116 3460 238168 3466
rect 238116 3402 238168 3408
rect 238128 480 238156 3402
rect 239324 480 239352 3538
rect 240520 480 240548 3606
rect 241716 480 241744 3742
rect 244096 3732 244148 3738
rect 244096 3674 244148 3680
rect 242900 3460 242952 3466
rect 242900 3402 242952 3408
rect 242912 480 242940 3402
rect 244108 480 244136 3674
rect 244660 3330 244688 334562
rect 244752 328778 244780 337640
rect 244844 337634 244872 337742
rect 245120 337742 245194 337770
rect 244844 337606 244964 337634
rect 244936 335714 244964 337606
rect 244924 335708 244976 335714
rect 244924 335650 244976 335656
rect 245016 335300 245068 335306
rect 245016 335242 245068 335248
rect 244924 333600 244976 333606
rect 244924 333542 244976 333548
rect 244740 328772 244792 328778
rect 244740 328714 244792 328720
rect 244648 3324 244700 3330
rect 244648 3266 244700 3272
rect 244936 3262 244964 333542
rect 245028 3874 245056 335242
rect 245120 327078 245148 337742
rect 245258 337668 245286 338028
rect 245350 337958 245378 338028
rect 245338 337952 245390 337958
rect 245338 337894 245390 337900
rect 245442 337822 245470 338028
rect 245534 337958 245562 338028
rect 245522 337952 245574 337958
rect 245522 337894 245574 337900
rect 245430 337816 245482 337822
rect 245626 337804 245654 338028
rect 245718 337929 245746 338028
rect 245704 337920 245760 337929
rect 245704 337855 245760 337864
rect 245430 337758 245482 337764
rect 245580 337776 245654 337804
rect 245212 337640 245286 337668
rect 245212 334626 245240 337640
rect 245292 335776 245344 335782
rect 245292 335718 245344 335724
rect 245200 334620 245252 334626
rect 245200 334562 245252 334568
rect 245200 334144 245252 334150
rect 245200 334086 245252 334092
rect 245212 333985 245240 334086
rect 245198 333976 245254 333985
rect 245198 333911 245254 333920
rect 245304 331214 245332 335718
rect 245476 334960 245528 334966
rect 245474 334928 245476 334937
rect 245528 334928 245530 334937
rect 245474 334863 245530 334872
rect 245580 333266 245608 337776
rect 245810 337770 245838 338028
rect 245902 337890 245930 338028
rect 245890 337884 245942 337890
rect 245890 337826 245942 337832
rect 245764 337742 245838 337770
rect 245994 337770 246022 338028
rect 246086 337929 246114 338028
rect 246072 337920 246128 337929
rect 246072 337855 246128 337864
rect 246178 337804 246206 338028
rect 246270 337929 246298 338028
rect 246362 337940 246390 338028
rect 246454 338008 246482 338028
rect 246454 337980 246528 338008
rect 246256 337920 246312 337929
rect 246362 337912 246436 337940
rect 246256 337855 246312 337864
rect 246132 337776 246206 337804
rect 245994 337742 246068 337770
rect 245658 337648 245714 337657
rect 245658 337583 245714 337592
rect 245568 333260 245620 333266
rect 245568 333202 245620 333208
rect 245474 332616 245530 332625
rect 245474 332551 245530 332560
rect 245212 331186 245332 331214
rect 245108 327072 245160 327078
rect 245108 327014 245160 327020
rect 245212 321554 245240 331186
rect 245120 321526 245240 321554
rect 245120 267034 245148 321526
rect 245488 316034 245516 332551
rect 245672 330750 245700 337583
rect 245764 333606 245792 337742
rect 245934 337648 245990 337657
rect 245934 337583 245990 337592
rect 245752 333600 245804 333606
rect 245752 333542 245804 333548
rect 245948 333402 245976 337583
rect 245936 333396 245988 333402
rect 245936 333338 245988 333344
rect 245660 330744 245712 330750
rect 245660 330686 245712 330692
rect 246040 326398 246068 337742
rect 246132 337668 246160 337776
rect 246132 337640 246252 337668
rect 246120 337544 246172 337550
rect 246120 337486 246172 337492
rect 246028 326392 246080 326398
rect 246028 326334 246080 326340
rect 245212 316006 245516 316034
rect 245212 272542 245240 316006
rect 245200 272536 245252 272542
rect 245200 272478 245252 272484
rect 245108 267028 245160 267034
rect 245108 266970 245160 266976
rect 245108 10328 245160 10334
rect 245108 10270 245160 10276
rect 245016 3868 245068 3874
rect 245016 3810 245068 3816
rect 245120 3466 245148 10270
rect 245200 4004 245252 4010
rect 245200 3946 245252 3952
rect 245108 3460 245160 3466
rect 245108 3402 245160 3408
rect 244924 3256 244976 3262
rect 244924 3198 244976 3204
rect 245212 480 245240 3946
rect 246132 3194 246160 337486
rect 246224 332246 246252 337640
rect 246408 335209 246436 337912
rect 246394 335200 246450 335209
rect 246394 335135 246450 335144
rect 246500 332314 246528 337980
rect 246638 337770 246666 338028
rect 246730 337890 246758 338028
rect 246718 337884 246770 337890
rect 246718 337826 246770 337832
rect 246822 337770 246850 338028
rect 246914 337890 246942 338028
rect 246902 337884 246954 337890
rect 246902 337826 246954 337832
rect 247006 337793 247034 338028
rect 246638 337742 246712 337770
rect 246488 332308 246540 332314
rect 246488 332250 246540 332256
rect 246212 332240 246264 332246
rect 246212 332182 246264 332188
rect 246304 331832 246356 331838
rect 246304 331774 246356 331780
rect 246212 326392 246264 326398
rect 246212 326334 246264 326340
rect 246224 4894 246252 326334
rect 246316 274650 246344 331774
rect 246684 330886 246712 337742
rect 246776 337742 246850 337770
rect 246992 337784 247048 337793
rect 246776 332382 246804 337742
rect 247098 337770 247126 338028
rect 247190 337890 247218 338028
rect 247178 337884 247230 337890
rect 247178 337826 247230 337832
rect 247282 337770 247310 338028
rect 247374 337895 247402 338028
rect 247360 337886 247416 337895
rect 247360 337821 247416 337830
rect 247466 337770 247494 338028
rect 247098 337742 247172 337770
rect 246992 337719 247048 337728
rect 246856 337544 246908 337550
rect 246856 337486 246908 337492
rect 247040 337544 247092 337550
rect 247040 337486 247092 337492
rect 246764 332376 246816 332382
rect 246764 332318 246816 332324
rect 246672 330880 246724 330886
rect 246672 330822 246724 330828
rect 246868 316034 246896 337486
rect 247052 330954 247080 337486
rect 247144 333538 247172 337742
rect 247236 337742 247310 337770
rect 247420 337742 247494 337770
rect 247236 335578 247264 337742
rect 247420 337668 247448 337742
rect 247558 337668 247586 338028
rect 247650 337804 247678 338028
rect 247742 337929 247770 338028
rect 247728 337920 247784 337929
rect 247728 337855 247784 337864
rect 247650 337776 247724 337804
rect 247328 337640 247448 337668
rect 247512 337640 247586 337668
rect 247224 335572 247276 335578
rect 247224 335514 247276 335520
rect 247132 333532 247184 333538
rect 247132 333474 247184 333480
rect 247328 331022 247356 337640
rect 247406 337512 247462 337521
rect 247406 337447 247462 337456
rect 247420 332450 247448 337447
rect 247512 333470 247540 337640
rect 247590 337512 247646 337521
rect 247590 337447 247646 337456
rect 247500 333464 247552 333470
rect 247500 333406 247552 333412
rect 247408 332444 247460 332450
rect 247408 332386 247460 332392
rect 247604 331090 247632 337447
rect 247696 332518 247724 337776
rect 247834 337770 247862 338028
rect 247926 337895 247954 338028
rect 247912 337886 247968 337895
rect 247912 337821 247968 337830
rect 247788 337742 247862 337770
rect 248018 337770 248046 338028
rect 248110 337890 248138 338028
rect 248098 337884 248150 337890
rect 248098 337826 248150 337832
rect 248202 337770 248230 338028
rect 248294 337958 248322 338028
rect 248282 337952 248334 337958
rect 248282 337894 248334 337900
rect 248386 337770 248414 338028
rect 248524 338014 248584 338042
rect 248524 337958 248552 338014
rect 248512 337952 248564 337958
rect 248662 337906 248690 338028
rect 248512 337894 248564 337900
rect 248616 337878 248690 337906
rect 248616 337804 248644 337878
rect 248018 337742 248092 337770
rect 247788 336734 247816 337742
rect 247958 337648 248014 337657
rect 247958 337583 248014 337592
rect 247776 336728 247828 336734
rect 247776 336670 247828 336676
rect 247972 332586 248000 337583
rect 247960 332580 248012 332586
rect 247960 332522 248012 332528
rect 247684 332512 247736 332518
rect 247684 332454 247736 332460
rect 247592 331084 247644 331090
rect 247592 331026 247644 331032
rect 247316 331016 247368 331022
rect 247316 330958 247368 330964
rect 247040 330948 247092 330954
rect 247040 330890 247092 330896
rect 248064 328642 248092 337742
rect 248156 337742 248230 337770
rect 248340 337742 248414 337770
rect 248524 337776 248644 337804
rect 248156 335850 248184 337742
rect 248144 335844 248196 335850
rect 248144 335786 248196 335792
rect 248340 334762 248368 337742
rect 248328 334756 248380 334762
rect 248328 334698 248380 334704
rect 248524 331770 248552 337776
rect 248754 337770 248782 338028
rect 248846 337890 248874 338028
rect 248938 337890 248966 338028
rect 248834 337884 248886 337890
rect 248834 337826 248886 337832
rect 248926 337884 248978 337890
rect 248926 337826 248978 337832
rect 248708 337742 248782 337770
rect 248708 336258 248736 337742
rect 249030 337668 249058 338028
rect 248892 337640 249058 337668
rect 249122 337668 249150 338028
rect 249214 337770 249242 338028
rect 249306 337890 249334 338028
rect 249398 337929 249426 338028
rect 249490 337958 249518 338028
rect 249478 337952 249530 337958
rect 249384 337920 249440 337929
rect 249294 337884 249346 337890
rect 249478 337894 249530 337900
rect 249384 337855 249440 337864
rect 249294 337826 249346 337832
rect 249430 337784 249486 337793
rect 249214 337742 249380 337770
rect 249122 337640 249196 337668
rect 248696 336252 248748 336258
rect 248696 336194 248748 336200
rect 248602 334112 248658 334121
rect 248892 334082 248920 337640
rect 249064 337544 249116 337550
rect 249064 337486 249116 337492
rect 249076 336784 249104 337486
rect 248984 336756 249104 336784
rect 248984 334694 249012 336756
rect 249064 336660 249116 336666
rect 249064 336602 249116 336608
rect 248972 334688 249024 334694
rect 248972 334630 249024 334636
rect 248602 334047 248658 334056
rect 248880 334076 248932 334082
rect 248512 331764 248564 331770
rect 248512 331706 248564 331712
rect 248052 328636 248104 328642
rect 248052 328578 248104 328584
rect 246684 316006 246896 316034
rect 246304 274644 246356 274650
rect 246304 274586 246356 274592
rect 246684 4962 246712 316006
rect 248616 271862 248644 334047
rect 248880 334018 248932 334024
rect 248788 326392 248840 326398
rect 248788 326334 248840 326340
rect 248604 271856 248656 271862
rect 248604 271798 248656 271804
rect 248800 5030 248828 326334
rect 249076 5166 249104 336602
rect 249168 333810 249196 337640
rect 249156 333804 249208 333810
rect 249156 333746 249208 333752
rect 249246 333296 249302 333305
rect 249246 333231 249302 333240
rect 249156 332716 249208 332722
rect 249156 332658 249208 332664
rect 249064 5160 249116 5166
rect 249064 5102 249116 5108
rect 248788 5024 248840 5030
rect 248788 4966 248840 4972
rect 246672 4956 246724 4962
rect 246672 4898 246724 4904
rect 246212 4888 246264 4894
rect 246212 4830 246264 4836
rect 247592 4140 247644 4146
rect 247592 4082 247644 4088
rect 246396 3868 246448 3874
rect 246396 3810 246448 3816
rect 246120 3188 246172 3194
rect 246120 3130 246172 3136
rect 246408 480 246436 3810
rect 247604 480 247632 4082
rect 249168 3534 249196 332658
rect 249260 236881 249288 333231
rect 249352 331226 249380 337742
rect 249582 337770 249610 338028
rect 249674 337890 249702 338028
rect 249662 337884 249714 337890
rect 249662 337826 249714 337832
rect 249766 337770 249794 338028
rect 249858 337958 249886 338028
rect 249950 337963 249978 338028
rect 249846 337952 249898 337958
rect 249846 337894 249898 337900
rect 249936 337954 249992 337963
rect 249936 337889 249992 337898
rect 249430 337719 249486 337728
rect 249536 337742 249610 337770
rect 249720 337742 249794 337770
rect 249890 337784 249946 337793
rect 249444 333878 249472 337719
rect 249536 334830 249564 337742
rect 249524 334824 249576 334830
rect 249524 334766 249576 334772
rect 249432 333872 249484 333878
rect 249432 333814 249484 333820
rect 249340 331220 249392 331226
rect 249340 331162 249392 331168
rect 249720 326398 249748 337742
rect 250042 337770 250070 338028
rect 250134 337890 250162 338028
rect 250122 337884 250174 337890
rect 250122 337826 250174 337832
rect 250226 337770 250254 338028
rect 249890 337719 249946 337728
rect 249996 337742 250070 337770
rect 250180 337742 250254 337770
rect 250318 337770 250346 338028
rect 250456 338014 250516 338042
rect 250318 337742 250392 337770
rect 249904 333198 249932 337719
rect 249892 333192 249944 333198
rect 249892 333134 249944 333140
rect 249996 333044 250024 337742
rect 250180 333130 250208 337742
rect 250364 337668 250392 337742
rect 250272 337640 250392 337668
rect 250168 333124 250220 333130
rect 250168 333066 250220 333072
rect 249904 333016 250024 333044
rect 249904 331702 249932 333016
rect 249984 332648 250036 332654
rect 249984 332590 250036 332596
rect 249892 331696 249944 331702
rect 249892 331638 249944 331644
rect 249708 326392 249760 326398
rect 249708 326334 249760 326340
rect 249246 236872 249302 236881
rect 249246 236807 249302 236816
rect 249996 3670 250024 332590
rect 250272 330410 250300 337640
rect 250456 335034 250484 338014
rect 250594 337804 250622 338028
rect 250686 337822 250714 338028
rect 250778 337958 250806 338028
rect 250766 337952 250818 337958
rect 250766 337894 250818 337900
rect 250548 337776 250622 337804
rect 250674 337816 250726 337822
rect 250444 335028 250496 335034
rect 250444 334970 250496 334976
rect 250548 334914 250576 337776
rect 250870 337770 250898 338028
rect 250962 337822 250990 338028
rect 251054 337963 251082 338028
rect 251040 337954 251096 337963
rect 251146 337958 251174 338028
rect 251238 337958 251266 338028
rect 251040 337889 251096 337898
rect 251134 337952 251186 337958
rect 251134 337894 251186 337900
rect 251226 337952 251278 337958
rect 251226 337894 251278 337900
rect 250674 337758 250726 337764
rect 250824 337742 250898 337770
rect 250950 337816 251002 337822
rect 251180 337816 251232 337822
rect 250950 337758 251002 337764
rect 251086 337784 251142 337793
rect 250628 335980 250680 335986
rect 250628 335922 250680 335928
rect 250456 334886 250576 334914
rect 250352 334076 250404 334082
rect 250352 334018 250404 334024
rect 250260 330404 250312 330410
rect 250260 330346 250312 330352
rect 250168 326392 250220 326398
rect 250168 326334 250220 326340
rect 250180 3942 250208 326334
rect 250364 321554 250392 334018
rect 250456 333062 250484 334886
rect 250536 334008 250588 334014
rect 250536 333950 250588 333956
rect 250444 333056 250496 333062
rect 250444 332998 250496 333004
rect 250364 321526 250484 321554
rect 250168 3936 250220 3942
rect 250168 3878 250220 3884
rect 250456 3806 250484 321526
rect 250444 3800 250496 3806
rect 250444 3742 250496 3748
rect 249984 3664 250036 3670
rect 249984 3606 250036 3612
rect 250548 3602 250576 333950
rect 250640 321554 250668 335922
rect 250824 332994 250852 337742
rect 251330 337804 251358 338028
rect 251422 337958 251450 338028
rect 251514 337958 251542 338028
rect 251410 337952 251462 337958
rect 251410 337894 251462 337900
rect 251502 337952 251554 337958
rect 251502 337894 251554 337900
rect 251180 337758 251232 337764
rect 251284 337776 251358 337804
rect 251086 337719 251142 337728
rect 251100 337498 251128 337719
rect 251008 337470 251128 337498
rect 250904 337340 250956 337346
rect 250904 337282 250956 337288
rect 250812 332988 250864 332994
rect 250812 332930 250864 332936
rect 250916 327554 250944 337282
rect 251008 335170 251036 337470
rect 251088 337340 251140 337346
rect 251088 337282 251140 337288
rect 250996 335164 251048 335170
rect 250996 335106 251048 335112
rect 250904 327548 250956 327554
rect 250904 327490 250956 327496
rect 251100 326398 251128 337282
rect 251192 331634 251220 337758
rect 251284 335714 251312 337776
rect 251606 337770 251634 338028
rect 251698 337958 251726 338028
rect 251686 337952 251738 337958
rect 251686 337894 251738 337900
rect 251560 337742 251634 337770
rect 251560 335918 251588 337742
rect 251790 337668 251818 338028
rect 251882 337822 251910 338028
rect 251870 337816 251922 337822
rect 251870 337758 251922 337764
rect 251974 337668 252002 338028
rect 252066 337770 252094 338028
rect 252158 338008 252186 338028
rect 252296 338014 252356 338042
rect 252158 337980 252232 338008
rect 252066 337742 252140 337770
rect 251790 337640 251864 337668
rect 251548 335912 251600 335918
rect 251548 335854 251600 335860
rect 251272 335708 251324 335714
rect 251272 335650 251324 335656
rect 251272 335096 251324 335102
rect 251272 335038 251324 335044
rect 251180 331628 251232 331634
rect 251180 331570 251232 331576
rect 251088 326392 251140 326398
rect 251088 326334 251140 326340
rect 250640 321526 250760 321554
rect 250732 270502 250760 321526
rect 251284 316034 251312 335038
rect 251836 334626 251864 337640
rect 251928 337640 252002 337668
rect 251824 334620 251876 334626
rect 251824 334562 251876 334568
rect 251928 333962 251956 337640
rect 252112 336954 252140 337742
rect 251836 333934 251956 333962
rect 252020 336926 252140 336954
rect 251836 331214 251864 333934
rect 251916 333192 251968 333198
rect 251916 333134 251968 333140
rect 251192 316006 251312 316034
rect 251560 331186 251864 331214
rect 250720 270496 250772 270502
rect 250720 270438 250772 270444
rect 251192 4146 251220 316006
rect 251180 4140 251232 4146
rect 251180 4082 251232 4088
rect 250536 3596 250588 3602
rect 250536 3538 250588 3544
rect 249156 3528 249208 3534
rect 249156 3470 249208 3476
rect 249984 3528 250036 3534
rect 249984 3470 250036 3476
rect 248788 3460 248840 3466
rect 248788 3402 248840 3408
rect 248800 480 248828 3402
rect 249996 480 250024 3470
rect 251180 3324 251232 3330
rect 251180 3266 251232 3272
rect 251192 480 251220 3266
rect 251560 3058 251588 331186
rect 251928 328454 251956 333134
rect 251836 328426 251956 328454
rect 251640 320204 251692 320210
rect 251640 320146 251692 320152
rect 251652 5098 251680 320146
rect 251836 318794 251864 328426
rect 252020 320210 252048 336926
rect 252100 334620 252152 334626
rect 252100 334562 252152 334568
rect 252112 330206 252140 334562
rect 252204 334490 252232 337980
rect 252192 334484 252244 334490
rect 252192 334426 252244 334432
rect 252296 331566 252324 338014
rect 252434 337906 252462 338028
rect 252526 337958 252554 338028
rect 252388 337878 252462 337906
rect 252514 337952 252566 337958
rect 252514 337894 252566 337900
rect 252284 331560 252336 331566
rect 252284 331502 252336 331508
rect 252100 330200 252152 330206
rect 252100 330142 252152 330148
rect 252388 330138 252416 337878
rect 252618 337804 252646 338028
rect 252572 337776 252646 337804
rect 252572 332790 252600 337776
rect 252710 337770 252738 338028
rect 252802 337890 252830 338028
rect 252894 337963 252922 338028
rect 252880 337954 252936 337963
rect 252790 337884 252842 337890
rect 252880 337889 252936 337898
rect 252790 337826 252842 337832
rect 252986 337770 253014 338028
rect 252710 337742 252784 337770
rect 252756 337668 252784 337742
rect 252664 337640 252784 337668
rect 252848 337742 253014 337770
rect 252560 332784 252612 332790
rect 252560 332726 252612 332732
rect 252468 332580 252520 332586
rect 252468 332522 252520 332528
rect 252376 330132 252428 330138
rect 252376 330074 252428 330080
rect 252008 320204 252060 320210
rect 252008 320146 252060 320152
rect 251836 318766 251956 318794
rect 251640 5092 251692 5098
rect 251640 5034 251692 5040
rect 251928 4010 251956 318766
rect 252480 6914 252508 332522
rect 252664 331498 252692 337640
rect 252744 334892 252796 334898
rect 252744 334834 252796 334840
rect 252652 331492 252704 331498
rect 252652 331434 252704 331440
rect 252756 331294 252784 334834
rect 252744 331288 252796 331294
rect 252744 331230 252796 331236
rect 252848 330070 252876 337742
rect 253078 337668 253106 338028
rect 253170 337770 253198 338028
rect 253262 337958 253290 338028
rect 253250 337952 253302 337958
rect 253250 337894 253302 337900
rect 253354 337770 253382 338028
rect 253446 337822 253474 338028
rect 253538 337958 253566 338028
rect 253526 337952 253578 337958
rect 253526 337894 253578 337900
rect 253170 337742 253244 337770
rect 252926 337648 252982 337657
rect 252926 337583 252982 337592
rect 253032 337640 253106 337668
rect 252940 333266 252968 337583
rect 253032 334354 253060 337640
rect 253112 337544 253164 337550
rect 253112 337486 253164 337492
rect 253020 334348 253072 334354
rect 253020 334290 253072 334296
rect 252928 333260 252980 333266
rect 252928 333202 252980 333208
rect 253124 331214 253152 337486
rect 253216 331430 253244 337742
rect 253308 337742 253382 337770
rect 253434 337816 253486 337822
rect 253630 337770 253658 338028
rect 253722 337822 253750 338028
rect 253814 337958 253842 338028
rect 253802 337952 253854 337958
rect 253802 337894 253854 337900
rect 253906 337890 253934 338028
rect 253894 337884 253946 337890
rect 253894 337826 253946 337832
rect 253434 337758 253486 337764
rect 253584 337742 253658 337770
rect 253710 337816 253762 337822
rect 253998 337770 254026 338028
rect 254090 338008 254118 338028
rect 254228 338014 254288 338042
rect 254090 337980 254164 338008
rect 253710 337758 253762 337764
rect 253952 337742 254026 337770
rect 253308 337634 253336 337742
rect 253308 337606 253428 337634
rect 253296 337544 253348 337550
rect 253296 337486 253348 337492
rect 253308 334898 253336 337486
rect 253296 334892 253348 334898
rect 253296 334834 253348 334840
rect 253400 334286 253428 337606
rect 253388 334280 253440 334286
rect 253388 334222 253440 334228
rect 253584 334218 253612 337742
rect 253756 337544 253808 337550
rect 253756 337486 253808 337492
rect 253572 334212 253624 334218
rect 253572 334154 253624 334160
rect 253388 333396 253440 333402
rect 253388 333338 253440 333344
rect 253204 331424 253256 331430
rect 253204 331366 253256 331372
rect 253204 331288 253256 331294
rect 253204 331230 253256 331236
rect 253032 331186 253152 331214
rect 252836 330064 252888 330070
rect 252836 330006 252888 330012
rect 253032 322250 253060 331186
rect 253020 322244 253072 322250
rect 253020 322186 253072 322192
rect 252652 9580 252704 9586
rect 252652 9522 252704 9528
rect 252388 6886 252508 6914
rect 251916 4004 251968 4010
rect 251916 3946 251968 3952
rect 251548 3052 251600 3058
rect 251548 2994 251600 3000
rect 252388 480 252416 6886
rect 252664 3874 252692 9522
rect 252652 3868 252704 3874
rect 252652 3810 252704 3816
rect 253216 3738 253244 331230
rect 253296 330200 253348 330206
rect 253296 330142 253348 330148
rect 253204 3732 253256 3738
rect 253204 3674 253256 3680
rect 253308 3398 253336 330142
rect 253400 3466 253428 333338
rect 253768 327486 253796 337486
rect 253952 333334 253980 337742
rect 254136 336666 254164 337980
rect 254124 336660 254176 336666
rect 254124 336602 254176 336608
rect 254228 335306 254256 338014
rect 254366 337872 254394 338028
rect 254458 337890 254486 338028
rect 254320 337844 254394 337872
rect 254446 337884 254498 337890
rect 254216 335300 254268 335306
rect 254216 335242 254268 335248
rect 254320 334744 254348 337844
rect 254446 337826 254498 337832
rect 254550 337793 254578 338028
rect 254642 337958 254670 338028
rect 254630 337952 254682 337958
rect 254630 337894 254682 337900
rect 254536 337784 254592 337793
rect 254734 337770 254762 338028
rect 254826 337958 254854 338028
rect 254918 337963 254946 338028
rect 254814 337952 254866 337958
rect 254814 337894 254866 337900
rect 254904 337954 254960 337963
rect 254904 337889 254960 337898
rect 255010 337890 255038 338028
rect 255102 337958 255130 338028
rect 255090 337952 255142 337958
rect 255090 337894 255142 337900
rect 254998 337884 255050 337890
rect 254998 337826 255050 337832
rect 255194 337804 255222 338028
rect 255286 337963 255314 338028
rect 255272 337954 255328 337963
rect 255378 337958 255406 338028
rect 255470 337963 255498 338028
rect 255272 337889 255328 337898
rect 255366 337952 255418 337958
rect 255366 337894 255418 337900
rect 255456 337954 255512 337963
rect 255456 337889 255512 337898
rect 255562 337890 255590 338028
rect 255654 337958 255682 338028
rect 255642 337952 255694 337958
rect 255642 337894 255694 337900
rect 255550 337884 255602 337890
rect 255550 337826 255602 337832
rect 255412 337816 255464 337822
rect 254536 337719 254592 337728
rect 254688 337742 254762 337770
rect 254858 337784 254914 337793
rect 254490 337648 254546 337657
rect 254490 337583 254546 337592
rect 254400 337340 254452 337346
rect 254400 337282 254452 337288
rect 254228 334716 254348 334744
rect 253940 333328 253992 333334
rect 253940 333270 253992 333276
rect 254228 332722 254256 334716
rect 254308 334620 254360 334626
rect 254308 334562 254360 334568
rect 254216 332716 254268 332722
rect 254216 332658 254268 332664
rect 253756 327480 253808 327486
rect 253756 327422 253808 327428
rect 254320 9586 254348 334562
rect 254412 330206 254440 337282
rect 254504 334014 254532 337583
rect 254582 335608 254638 335617
rect 254582 335543 254638 335552
rect 254492 334008 254544 334014
rect 254492 333950 254544 333956
rect 254400 330200 254452 330206
rect 254400 330142 254452 330148
rect 254596 326346 254624 335543
rect 254688 334082 254716 337742
rect 255194 337776 255268 337804
rect 254858 337719 254914 337728
rect 254872 337550 254900 337719
rect 254860 337544 254912 337550
rect 254860 337486 254912 337492
rect 254860 337340 254912 337346
rect 254860 337282 254912 337288
rect 254952 337340 255004 337346
rect 254952 337282 255004 337288
rect 254768 337204 254820 337210
rect 254768 337146 254820 337152
rect 254676 334076 254728 334082
rect 254676 334018 254728 334024
rect 254596 326318 254716 326346
rect 254584 326256 254636 326262
rect 254584 326198 254636 326204
rect 254492 323196 254544 323202
rect 254492 323138 254544 323144
rect 254504 10334 254532 323138
rect 254492 10328 254544 10334
rect 254492 10270 254544 10276
rect 254308 9580 254360 9586
rect 254308 9522 254360 9528
rect 253480 8492 253532 8498
rect 253480 8434 253532 8440
rect 253388 3460 253440 3466
rect 253388 3402 253440 3408
rect 253296 3392 253348 3398
rect 253296 3334 253348 3340
rect 253492 480 253520 8434
rect 254596 3534 254624 326198
rect 254688 239057 254716 326318
rect 254780 323202 254808 337146
rect 254872 332654 254900 337282
rect 254964 333198 254992 337282
rect 255240 336734 255268 337776
rect 255318 337784 255374 337793
rect 255746 337804 255774 338028
rect 255838 337963 255866 338028
rect 255824 337954 255880 337963
rect 255930 337958 255958 338028
rect 256022 338008 256050 338028
rect 256160 338014 256220 338042
rect 256022 337980 256096 338008
rect 255824 337889 255880 337898
rect 255918 337952 255970 337958
rect 255918 337894 255970 337900
rect 255412 337758 255464 337764
rect 255502 337784 255558 337793
rect 255318 337719 255374 337728
rect 255148 336706 255268 336734
rect 255148 335102 255176 336706
rect 255136 335096 255188 335102
rect 255136 335038 255188 335044
rect 255332 333402 255360 337719
rect 255320 333396 255372 333402
rect 255320 333338 255372 333344
rect 255228 333260 255280 333266
rect 255228 333202 255280 333208
rect 254952 333192 255004 333198
rect 254952 333134 255004 333140
rect 254860 332648 254912 332654
rect 254860 332590 254912 332596
rect 255240 326262 255268 333202
rect 255424 332586 255452 337758
rect 255502 337719 255558 337728
rect 255700 337776 255774 337804
rect 255964 337816 256016 337822
rect 255870 337784 255926 337793
rect 255412 332580 255464 332586
rect 255412 332522 255464 332528
rect 255412 326460 255464 326466
rect 255412 326402 255464 326408
rect 255228 326256 255280 326262
rect 255228 326198 255280 326204
rect 255424 326074 255452 326402
rect 255516 326346 255544 337719
rect 255596 337340 255648 337346
rect 255596 337282 255648 337288
rect 255608 326466 255636 337282
rect 255700 336734 255728 337776
rect 255964 337758 256016 337764
rect 255870 337719 255926 337728
rect 255700 336706 255820 336734
rect 255688 335368 255740 335374
rect 255688 335310 255740 335316
rect 255700 326534 255728 335310
rect 255688 326528 255740 326534
rect 255688 326470 255740 326476
rect 255596 326460 255648 326466
rect 255596 326402 255648 326408
rect 255516 326318 255728 326346
rect 255424 326046 255636 326074
rect 254768 323196 254820 323202
rect 254768 323138 254820 323144
rect 255504 322992 255556 322998
rect 255504 322934 255556 322940
rect 254674 239048 254730 239057
rect 254674 238983 254730 238992
rect 255516 3534 255544 322934
rect 255608 8498 255636 326046
rect 255596 8492 255648 8498
rect 255596 8434 255648 8440
rect 254584 3528 254636 3534
rect 254584 3470 254636 3476
rect 254676 3528 254728 3534
rect 254676 3470 254728 3476
rect 255504 3528 255556 3534
rect 255504 3470 255556 3476
rect 254688 480 254716 3470
rect 255700 3330 255728 326318
rect 255792 322998 255820 336706
rect 255884 326346 255912 337719
rect 255976 335918 256004 337758
rect 255964 335912 256016 335918
rect 255964 335854 256016 335860
rect 256068 333266 256096 337980
rect 256160 335850 256188 338014
rect 256298 337890 256326 338028
rect 256286 337884 256338 337890
rect 256286 337826 256338 337832
rect 256390 337770 256418 338028
rect 256482 337958 256510 338028
rect 256470 337952 256522 337958
rect 256470 337894 256522 337900
rect 256252 337742 256418 337770
rect 256148 335844 256200 335850
rect 256148 335786 256200 335792
rect 256146 335744 256202 335753
rect 256146 335679 256202 335688
rect 256056 333260 256108 333266
rect 256056 333202 256108 333208
rect 256160 330449 256188 335679
rect 256146 330440 256202 330449
rect 256146 330375 256202 330384
rect 256252 328454 256280 337742
rect 256574 337668 256602 338028
rect 256666 337890 256694 338028
rect 256654 337884 256706 337890
rect 256654 337826 256706 337832
rect 256758 337770 256786 338028
rect 256528 337640 256602 337668
rect 256712 337742 256786 337770
rect 256850 337770 256878 338028
rect 256942 337963 256970 338028
rect 256928 337954 256984 337963
rect 256928 337889 256984 337898
rect 257034 337890 257062 338028
rect 257126 337958 257154 338028
rect 257114 337952 257166 337958
rect 257114 337894 257166 337900
rect 257022 337884 257074 337890
rect 257022 337826 257074 337832
rect 257218 337822 257246 338028
rect 257310 337958 257338 338028
rect 257298 337952 257350 337958
rect 257298 337894 257350 337900
rect 257206 337816 257258 337822
rect 256974 337784 257030 337793
rect 256850 337742 256924 337770
rect 256424 337544 256476 337550
rect 256424 337486 256476 337492
rect 255976 328426 256280 328454
rect 255976 326466 256004 328426
rect 255964 326460 256016 326466
rect 255964 326402 256016 326408
rect 256332 326392 256384 326398
rect 255884 326318 256096 326346
rect 256332 326334 256384 326340
rect 255872 326256 255924 326262
rect 255872 326198 255924 326204
rect 255780 322992 255832 322998
rect 255780 322934 255832 322940
rect 255884 3466 255912 326198
rect 256068 321554 256096 326318
rect 256068 321526 256188 321554
rect 256160 6914 256188 321526
rect 255976 6886 256188 6914
rect 255872 3460 255924 3466
rect 255872 3402 255924 3408
rect 255976 3346 256004 6886
rect 256344 5370 256372 326334
rect 256332 5364 256384 5370
rect 256332 5306 256384 5312
rect 256436 3602 256464 337486
rect 256528 326398 256556 337640
rect 256608 333260 256660 333266
rect 256608 333202 256660 333208
rect 256516 326392 256568 326398
rect 256516 326334 256568 326340
rect 256620 316034 256648 333202
rect 256712 330954 256740 337742
rect 256792 336048 256844 336054
rect 256792 335990 256844 335996
rect 256804 332314 256832 335990
rect 256896 335374 256924 337742
rect 257402 337804 257430 338028
rect 257494 337958 257522 338028
rect 257586 337958 257614 338028
rect 257678 337963 257706 338028
rect 257482 337952 257534 337958
rect 257482 337894 257534 337900
rect 257574 337952 257626 337958
rect 257574 337894 257626 337900
rect 257664 337954 257720 337963
rect 257664 337889 257720 337898
rect 257402 337776 257476 337804
rect 257206 337758 257258 337764
rect 256974 337719 257030 337728
rect 256884 335368 256936 335374
rect 256884 335310 256936 335316
rect 256988 333334 257016 337719
rect 257252 335776 257304 335782
rect 257252 335718 257304 335724
rect 256976 333328 257028 333334
rect 256976 333270 257028 333276
rect 257068 333192 257120 333198
rect 257068 333134 257120 333140
rect 256792 332308 256844 332314
rect 256792 332250 256844 332256
rect 256700 330948 256752 330954
rect 256700 330890 256752 330896
rect 256528 316006 256648 316034
rect 256424 3596 256476 3602
rect 256424 3538 256476 3544
rect 256528 3534 256556 316006
rect 257080 5506 257108 333134
rect 257068 5500 257120 5506
rect 257068 5442 257120 5448
rect 257264 5098 257292 335718
rect 257344 335368 257396 335374
rect 257344 335310 257396 335316
rect 257252 5092 257304 5098
rect 257252 5034 257304 5040
rect 257356 4894 257384 335310
rect 257448 328454 257476 337776
rect 257664 337784 257720 337793
rect 257664 337719 257720 337728
rect 257678 337668 257706 337719
rect 257632 337640 257706 337668
rect 257770 337668 257798 338028
rect 257862 337958 257890 338028
rect 257850 337952 257902 337958
rect 257850 337894 257902 337900
rect 257954 337770 257982 338028
rect 257908 337742 257982 337770
rect 257770 337640 257844 337668
rect 257448 328426 257568 328454
rect 257436 326460 257488 326466
rect 257436 326402 257488 326408
rect 257448 5234 257476 326402
rect 257436 5228 257488 5234
rect 257436 5170 257488 5176
rect 257344 4888 257396 4894
rect 257344 4830 257396 4836
rect 257540 4418 257568 328426
rect 257632 326466 257660 337640
rect 257712 337544 257764 337550
rect 257712 337486 257764 337492
rect 257620 326460 257672 326466
rect 257620 326402 257672 326408
rect 257724 326346 257752 337486
rect 257632 326318 257752 326346
rect 257816 326346 257844 337640
rect 257908 335782 257936 337742
rect 258138 337668 258166 338028
rect 258230 337963 258258 338028
rect 258216 337954 258272 337963
rect 258216 337889 258272 337898
rect 258322 337822 258350 338028
rect 258414 337963 258442 338028
rect 258400 337954 258456 337963
rect 258400 337889 258456 337898
rect 258506 337890 258534 338028
rect 258598 337963 258626 338028
rect 258584 337954 258640 337963
rect 258690 337958 258718 338028
rect 258494 337884 258546 337890
rect 258584 337889 258640 337898
rect 258678 337952 258730 337958
rect 258678 337894 258730 337900
rect 258782 337890 258810 338028
rect 258874 337958 258902 338028
rect 258966 337963 258994 338028
rect 258862 337952 258914 337958
rect 258862 337894 258914 337900
rect 258952 337954 259008 337963
rect 258494 337826 258546 337832
rect 258770 337884 258822 337890
rect 258952 337889 259008 337898
rect 258770 337826 258822 337832
rect 258310 337816 258362 337822
rect 258310 337758 258362 337764
rect 258446 337784 258502 337793
rect 258446 337719 258502 337728
rect 258814 337784 258870 337793
rect 259058 337770 259086 338028
rect 259150 337963 259178 338028
rect 259136 337954 259192 337963
rect 259242 337958 259270 338028
rect 259334 337963 259362 338028
rect 259136 337889 259192 337898
rect 259230 337952 259282 337958
rect 259230 337894 259282 337900
rect 259320 337954 259376 337963
rect 259426 337958 259454 338028
rect 259518 337963 259546 338028
rect 259320 337889 259376 337898
rect 259414 337952 259466 337958
rect 259414 337894 259466 337900
rect 259504 337954 259560 337963
rect 259610 337958 259638 338028
rect 259504 337889 259560 337898
rect 259598 337952 259650 337958
rect 259598 337894 259650 337900
rect 259366 337784 259422 337793
rect 259058 337742 259132 337770
rect 258814 337719 258870 337728
rect 258138 337640 258212 337668
rect 257896 335776 257948 335782
rect 257896 335718 257948 335724
rect 257896 335640 257948 335646
rect 257896 335582 257948 335588
rect 257908 326466 257936 335582
rect 257988 333328 258040 333334
rect 257988 333270 258040 333276
rect 257896 326460 257948 326466
rect 257896 326402 257948 326408
rect 257816 326318 257936 326346
rect 257632 5166 257660 326318
rect 257712 326256 257764 326262
rect 257712 326198 257764 326204
rect 257804 326256 257856 326262
rect 257804 326198 257856 326204
rect 257620 5160 257672 5166
rect 257620 5102 257672 5108
rect 257724 5030 257752 326198
rect 257816 5302 257844 326198
rect 257804 5296 257856 5302
rect 257804 5238 257856 5244
rect 257712 5024 257764 5030
rect 257712 4966 257764 4972
rect 257908 4962 257936 326318
rect 258000 326262 258028 333270
rect 258184 329322 258212 337640
rect 258460 331430 258488 337719
rect 258632 337544 258684 337550
rect 258632 337486 258684 337492
rect 258448 331424 258500 331430
rect 258448 331366 258500 331372
rect 258264 331288 258316 331294
rect 258264 331230 258316 331236
rect 258172 329316 258224 329322
rect 258172 329258 258224 329264
rect 257988 326256 258040 326262
rect 257988 326198 258040 326204
rect 258276 16574 258304 331230
rect 258448 329316 258500 329322
rect 258448 329258 258500 329264
rect 258460 236774 258488 329258
rect 258448 236768 258500 236774
rect 258448 236710 258500 236716
rect 258276 16546 258396 16574
rect 257896 4956 257948 4962
rect 257896 4898 257948 4904
rect 257528 4412 257580 4418
rect 257528 4354 257580 4360
rect 257068 4072 257120 4078
rect 257068 4014 257120 4020
rect 256516 3528 256568 3534
rect 256516 3470 256568 3476
rect 255688 3324 255740 3330
rect 255688 3266 255740 3272
rect 255884 3318 256004 3346
rect 255884 480 255912 3318
rect 257080 480 257108 4014
rect 258264 3528 258316 3534
rect 258264 3470 258316 3476
rect 258276 480 258304 3470
rect 258368 3330 258396 16546
rect 258644 4826 258672 337486
rect 258724 335844 258776 335850
rect 258724 335786 258776 335792
rect 258632 4820 258684 4826
rect 258632 4762 258684 4768
rect 258736 3534 258764 335786
rect 258828 334830 258856 337719
rect 259104 337668 259132 337742
rect 259366 337719 259422 337728
rect 259550 337784 259606 337793
rect 259702 337770 259730 338028
rect 259794 337872 259822 338028
rect 259886 338008 259914 338028
rect 259886 337980 259960 338008
rect 259794 337844 259868 337872
rect 259702 337742 259776 337770
rect 259550 337719 259606 337728
rect 258998 337648 259054 337657
rect 259104 337640 259316 337668
rect 258998 337583 259054 337592
rect 258816 334824 258868 334830
rect 258816 334766 258868 334772
rect 258816 333940 258868 333946
rect 258816 333882 258868 333888
rect 258828 238066 258856 333882
rect 259012 330002 259040 337583
rect 259090 337512 259146 337521
rect 259090 337447 259146 337456
rect 259000 329996 259052 330002
rect 259000 329938 259052 329944
rect 259104 321554 259132 337447
rect 259182 337376 259238 337385
rect 259182 337311 259238 337320
rect 258920 321526 259132 321554
rect 258816 238060 258868 238066
rect 258816 238002 258868 238008
rect 258724 3528 258776 3534
rect 258724 3470 258776 3476
rect 258356 3324 258408 3330
rect 258356 3266 258408 3272
rect 258920 2922 258948 321526
rect 259196 316034 259224 337311
rect 259288 336666 259316 337640
rect 259380 337532 259408 337719
rect 259564 337668 259592 337719
rect 259564 337640 259684 337668
rect 259380 337504 259592 337532
rect 259276 336660 259328 336666
rect 259276 336602 259328 336608
rect 259460 335912 259512 335918
rect 259460 335854 259512 335860
rect 259104 316006 259224 316034
rect 259104 238134 259132 316006
rect 259092 238128 259144 238134
rect 259092 238070 259144 238076
rect 259472 4078 259500 335854
rect 259564 335714 259592 337504
rect 259552 335708 259604 335714
rect 259552 335650 259604 335656
rect 259552 333192 259604 333198
rect 259552 333134 259604 333140
rect 259564 6730 259592 333134
rect 259656 331702 259684 337640
rect 259748 332790 259776 337742
rect 259736 332784 259788 332790
rect 259736 332726 259788 332732
rect 259644 331696 259696 331702
rect 259644 331638 259696 331644
rect 259840 330070 259868 337844
rect 259932 336598 259960 337980
rect 260070 337958 260098 338028
rect 260058 337952 260110 337958
rect 260058 337894 260110 337900
rect 260162 337668 260190 338028
rect 260116 337640 260190 337668
rect 260254 337668 260282 338028
rect 260346 337958 260374 338028
rect 260334 337952 260386 337958
rect 260334 337894 260386 337900
rect 260438 337770 260466 338028
rect 260392 337742 260466 337770
rect 260530 337770 260558 338028
rect 260622 337890 260650 338028
rect 260610 337884 260662 337890
rect 260610 337826 260662 337832
rect 260714 337770 260742 338028
rect 260530 337742 260604 337770
rect 260254 337640 260328 337668
rect 259920 336592 259972 336598
rect 259920 336534 259972 336540
rect 260012 334688 260064 334694
rect 260012 334630 260064 334636
rect 259828 330064 259880 330070
rect 259828 330006 259880 330012
rect 260024 326466 260052 334630
rect 260012 326460 260064 326466
rect 260012 326402 260064 326408
rect 260116 326346 260144 337640
rect 260300 336122 260328 337640
rect 260288 336116 260340 336122
rect 260288 336058 260340 336064
rect 260392 335374 260420 337742
rect 260576 337634 260604 337742
rect 260484 337606 260604 337634
rect 260668 337742 260742 337770
rect 260380 335368 260432 335374
rect 260380 335310 260432 335316
rect 260196 326460 260248 326466
rect 260196 326402 260248 326408
rect 259932 326318 260144 326346
rect 259552 6724 259604 6730
rect 259552 6666 259604 6672
rect 259932 4350 259960 326318
rect 260012 326256 260064 326262
rect 260012 326198 260064 326204
rect 260024 4486 260052 326198
rect 260208 316034 260236 326402
rect 260484 326262 260512 337606
rect 260564 337544 260616 337550
rect 260564 337486 260616 337492
rect 260576 335510 260604 337486
rect 260564 335504 260616 335510
rect 260564 335446 260616 335452
rect 260564 335368 260616 335374
rect 260564 335310 260616 335316
rect 260576 330138 260604 335310
rect 260564 330132 260616 330138
rect 260564 330074 260616 330080
rect 260472 326256 260524 326262
rect 260472 326198 260524 326204
rect 260668 316034 260696 337742
rect 260806 337668 260834 338028
rect 260898 337822 260926 338028
rect 260886 337816 260938 337822
rect 260886 337758 260938 337764
rect 260760 337640 260834 337668
rect 260990 337668 261018 338028
rect 261082 337770 261110 338028
rect 261174 337890 261202 338028
rect 261266 337958 261294 338028
rect 261254 337952 261306 337958
rect 261254 337894 261306 337900
rect 261162 337884 261214 337890
rect 261162 337826 261214 337832
rect 261358 337770 261386 338028
rect 261450 337890 261478 338028
rect 261438 337884 261490 337890
rect 261438 337826 261490 337832
rect 261542 337770 261570 338028
rect 261634 337872 261662 338028
rect 261726 337940 261754 338028
rect 261818 338008 261846 338028
rect 261956 338014 262016 338042
rect 261818 337980 261892 338008
rect 261726 337912 261800 337940
rect 261634 337844 261708 337872
rect 261082 337742 261156 337770
rect 261358 337742 261478 337770
rect 261542 337742 261616 337770
rect 260990 337640 261064 337668
rect 260760 335646 260788 337640
rect 260840 336252 260892 336258
rect 260840 336194 260892 336200
rect 260748 335640 260800 335646
rect 260748 335582 260800 335588
rect 260748 335504 260800 335510
rect 260748 335446 260800 335452
rect 260760 332858 260788 335446
rect 260748 332852 260800 332858
rect 260748 332794 260800 332800
rect 260852 331906 260880 336194
rect 261036 335374 261064 337640
rect 261128 336394 261156 337742
rect 261450 337668 261478 337742
rect 261450 337640 261524 337668
rect 261496 337532 261524 337640
rect 261404 337504 261524 337532
rect 261116 336388 261168 336394
rect 261116 336330 261168 336336
rect 261116 335708 261168 335714
rect 261116 335650 261168 335656
rect 261024 335368 261076 335374
rect 261024 335310 261076 335316
rect 260840 331900 260892 331906
rect 260840 331842 260892 331848
rect 261128 331634 261156 335650
rect 261208 333192 261260 333198
rect 261208 333134 261260 333140
rect 261116 331628 261168 331634
rect 261116 331570 261168 331576
rect 261220 321554 261248 333134
rect 261404 328982 261432 337504
rect 261484 335368 261536 335374
rect 261484 335310 261536 335316
rect 261392 328976 261444 328982
rect 261392 328918 261444 328924
rect 261496 326346 261524 335310
rect 261588 326482 261616 337742
rect 261680 336326 261708 337844
rect 261668 336320 261720 336326
rect 261668 336262 261720 336268
rect 261772 335374 261800 337912
rect 261760 335368 261812 335374
rect 261760 335310 261812 335316
rect 261760 335096 261812 335102
rect 261760 335038 261812 335044
rect 261588 326454 261708 326482
rect 261496 326318 261616 326346
rect 261220 321526 261524 321554
rect 260116 316006 260236 316034
rect 260484 316006 260696 316034
rect 260116 232558 260144 316006
rect 260104 232552 260156 232558
rect 260104 232494 260156 232500
rect 260484 11014 260512 316006
rect 260472 11008 260524 11014
rect 260472 10950 260524 10956
rect 261496 10674 261524 321526
rect 261588 10946 261616 326318
rect 261576 10940 261628 10946
rect 261576 10882 261628 10888
rect 261680 10810 261708 326454
rect 261772 10878 261800 335038
rect 261760 10872 261812 10878
rect 261760 10814 261812 10820
rect 261668 10804 261720 10810
rect 261668 10746 261720 10752
rect 261864 10742 261892 337980
rect 261956 336190 261984 338014
rect 262094 337770 262122 338028
rect 262186 337890 262214 338028
rect 262278 337958 262306 338028
rect 262266 337952 262318 337958
rect 262266 337894 262318 337900
rect 262174 337884 262226 337890
rect 262174 337826 262226 337832
rect 262370 337770 262398 338028
rect 262462 337958 262490 338028
rect 262554 337958 262582 338028
rect 262450 337952 262502 337958
rect 262450 337894 262502 337900
rect 262542 337952 262594 337958
rect 262542 337894 262594 337900
rect 262646 337890 262674 338028
rect 262634 337884 262686 337890
rect 262634 337826 262686 337832
rect 262738 337770 262766 338028
rect 262830 337890 262858 338028
rect 262818 337884 262870 337890
rect 262818 337826 262870 337832
rect 262922 337770 262950 338028
rect 262094 337742 262168 337770
rect 261944 336184 261996 336190
rect 261944 336126 261996 336132
rect 262036 335980 262088 335986
rect 262036 335922 262088 335928
rect 261944 335368 261996 335374
rect 261944 335310 261996 335316
rect 261852 10736 261904 10742
rect 261852 10678 261904 10684
rect 261484 10668 261536 10674
rect 261484 10610 261536 10616
rect 261956 6594 261984 335310
rect 262048 6662 262076 335922
rect 262036 6656 262088 6662
rect 262036 6598 262088 6604
rect 261944 6588 261996 6594
rect 261944 6530 261996 6536
rect 262140 6526 262168 337742
rect 262324 337742 262398 337770
rect 262692 337742 262766 337770
rect 262876 337742 262950 337770
rect 263014 337770 263042 338028
rect 263106 337890 263134 338028
rect 263094 337884 263146 337890
rect 263094 337826 263146 337832
rect 263198 337770 263226 338028
rect 263014 337742 263088 337770
rect 262220 336252 262272 336258
rect 262220 336194 262272 336200
rect 262128 6520 262180 6526
rect 262128 6462 262180 6468
rect 262232 6186 262260 336194
rect 262324 326398 262352 337742
rect 262404 335640 262456 335646
rect 262404 335582 262456 335588
rect 262312 326392 262364 326398
rect 262312 326334 262364 326340
rect 262416 6254 262444 335582
rect 262588 335300 262640 335306
rect 262588 335242 262640 335248
rect 262600 330206 262628 335242
rect 262588 330200 262640 330206
rect 262588 330142 262640 330148
rect 262692 10538 262720 337742
rect 262772 337544 262824 337550
rect 262772 337486 262824 337492
rect 262784 10606 262812 337486
rect 262876 335442 262904 337742
rect 262956 337544 263008 337550
rect 262956 337486 263008 337492
rect 262968 336122 262996 337486
rect 262956 336116 263008 336122
rect 262956 336058 263008 336064
rect 262956 335844 263008 335850
rect 262956 335786 263008 335792
rect 262864 335436 262916 335442
rect 262864 335378 262916 335384
rect 262864 333192 262916 333198
rect 262864 333134 262916 333140
rect 262772 10600 262824 10606
rect 262772 10542 262824 10548
rect 262680 10532 262732 10538
rect 262680 10474 262732 10480
rect 262876 10334 262904 333134
rect 262968 10402 262996 335786
rect 263060 10470 263088 337742
rect 263152 337742 263226 337770
rect 263152 335646 263180 337742
rect 263290 337668 263318 338028
rect 263244 337640 263318 337668
rect 263244 335850 263272 337640
rect 263382 337634 263410 338028
rect 263474 337770 263502 338028
rect 263566 337929 263594 338028
rect 263552 337920 263608 337929
rect 263658 337890 263686 338028
rect 263750 338008 263778 338028
rect 263888 338014 263948 338042
rect 263750 337980 263824 338008
rect 263552 337855 263608 337864
rect 263646 337884 263698 337890
rect 263646 337826 263698 337832
rect 263690 337784 263746 337793
rect 263474 337742 263548 337770
rect 263382 337606 263456 337634
rect 263324 336728 263376 336734
rect 263324 336670 263376 336676
rect 263232 335844 263284 335850
rect 263232 335786 263284 335792
rect 263140 335640 263192 335646
rect 263140 335582 263192 335588
rect 263336 335594 263364 336670
rect 263428 336462 263456 337606
rect 263416 336456 263468 336462
rect 263416 336398 263468 336404
rect 263520 336258 263548 337742
rect 263690 337719 263746 337728
rect 263508 336252 263560 336258
rect 263508 336194 263560 336200
rect 263336 335566 263548 335594
rect 263324 335436 263376 335442
rect 263324 335378 263376 335384
rect 263232 332988 263284 332994
rect 263232 332930 263284 332936
rect 263140 326392 263192 326398
rect 263140 326334 263192 326340
rect 263048 10464 263100 10470
rect 263048 10406 263100 10412
rect 262956 10396 263008 10402
rect 262956 10338 263008 10344
rect 262864 10328 262916 10334
rect 262864 10270 262916 10276
rect 263152 6458 263180 326334
rect 263140 6452 263192 6458
rect 263140 6394 263192 6400
rect 263244 6390 263272 332930
rect 263232 6384 263284 6390
rect 263232 6326 263284 6332
rect 263336 6322 263364 335378
rect 263520 335354 263548 335566
rect 263520 335326 263640 335354
rect 263612 335186 263640 335326
rect 263520 335158 263640 335186
rect 263520 331498 263548 335158
rect 263704 333198 263732 337719
rect 263796 335442 263824 337980
rect 263784 335436 263836 335442
rect 263784 335378 263836 335384
rect 263888 335374 263916 338014
rect 264026 337770 264054 338028
rect 263980 337742 264054 337770
rect 263980 336666 264008 337742
rect 264118 337634 264146 338028
rect 264210 337958 264238 338028
rect 264302 337963 264330 338028
rect 264198 337952 264250 337958
rect 264198 337894 264250 337900
rect 264288 337954 264344 337963
rect 264288 337889 264344 337898
rect 264394 337890 264422 338028
rect 264382 337884 264434 337890
rect 264382 337826 264434 337832
rect 264486 337668 264514 338028
rect 264578 337770 264606 338028
rect 264670 337963 264698 338028
rect 264656 337954 264712 337963
rect 264762 337958 264790 338028
rect 264854 337963 264882 338028
rect 264656 337889 264712 337898
rect 264750 337952 264802 337958
rect 264750 337894 264802 337900
rect 264840 337954 264896 337963
rect 264946 337958 264974 338028
rect 265038 337958 265066 338028
rect 264840 337889 264896 337898
rect 264934 337952 264986 337958
rect 264934 337894 264986 337900
rect 265026 337952 265078 337958
rect 265026 337894 265078 337900
rect 264794 337784 264850 337793
rect 264578 337742 264652 337770
rect 264486 337640 264560 337668
rect 264118 337606 264192 337634
rect 263968 336660 264020 336666
rect 263968 336602 264020 336608
rect 263876 335368 263928 335374
rect 263876 335310 263928 335316
rect 263692 333192 263744 333198
rect 263692 333134 263744 333140
rect 264164 332994 264192 337606
rect 264532 336818 264560 337640
rect 264624 336938 264652 337742
rect 264794 337719 264850 337728
rect 264978 337784 265034 337793
rect 265130 337770 265158 338028
rect 265222 337958 265250 338028
rect 265210 337952 265262 337958
rect 265210 337894 265262 337900
rect 264978 337719 265034 337728
rect 265084 337742 265158 337770
rect 265314 337770 265342 338028
rect 265406 337958 265434 338028
rect 265394 337952 265446 337958
rect 265394 337894 265446 337900
rect 265498 337770 265526 338028
rect 265590 337872 265618 338028
rect 265682 338008 265710 338028
rect 265820 338014 265880 338042
rect 265682 337980 265756 338008
rect 265590 337844 265664 337872
rect 265314 337742 265388 337770
rect 265498 337742 265572 337770
rect 264612 336932 264664 336938
rect 264612 336874 264664 336880
rect 264532 336790 264652 336818
rect 264244 336320 264296 336326
rect 264244 336262 264296 336268
rect 264152 332988 264204 332994
rect 264152 332930 264204 332936
rect 263508 331492 263560 331498
rect 263508 331434 263560 331440
rect 263324 6316 263376 6322
rect 263324 6258 263376 6264
rect 262404 6248 262456 6254
rect 262404 6190 262456 6196
rect 262220 6180 262272 6186
rect 262220 6122 262272 6128
rect 264152 5364 264204 5370
rect 264152 5306 264204 5312
rect 260012 4480 260064 4486
rect 260012 4422 260064 4428
rect 259920 4344 259972 4350
rect 259920 4286 259972 4292
rect 259460 4072 259512 4078
rect 259460 4014 259512 4020
rect 260656 3596 260708 3602
rect 260656 3538 260708 3544
rect 259460 3528 259512 3534
rect 259460 3470 259512 3476
rect 258908 2916 258960 2922
rect 258908 2858 258960 2864
rect 259472 480 259500 3470
rect 260668 480 260696 3538
rect 261760 3460 261812 3466
rect 261760 3402 261812 3408
rect 261772 480 261800 3402
rect 262956 3324 263008 3330
rect 262956 3266 263008 3272
rect 262968 480 262996 3266
rect 264164 480 264192 5306
rect 264256 4554 264284 336262
rect 264520 335844 264572 335850
rect 264520 335786 264572 335792
rect 264336 335368 264388 335374
rect 264336 335310 264388 335316
rect 264348 330274 264376 335310
rect 264428 333328 264480 333334
rect 264428 333270 264480 333276
rect 264336 330268 264388 330274
rect 264336 330210 264388 330216
rect 264244 4548 264296 4554
rect 264244 4490 264296 4496
rect 264440 3262 264468 333270
rect 264532 93158 264560 335786
rect 264624 330410 264652 336790
rect 264808 333946 264836 337719
rect 264992 335918 265020 337719
rect 265084 337006 265112 337742
rect 265072 337000 265124 337006
rect 265072 336942 265124 336948
rect 264980 335912 265032 335918
rect 264980 335854 265032 335860
rect 264796 333940 264848 333946
rect 264796 333882 264848 333888
rect 264704 333260 264756 333266
rect 264704 333202 264756 333208
rect 264612 330404 264664 330410
rect 264612 330346 264664 330352
rect 264520 93152 264572 93158
rect 264520 93094 264572 93100
rect 264716 3534 264744 333202
rect 265360 331838 265388 337742
rect 265440 337544 265492 337550
rect 265440 337486 265492 337492
rect 265348 331832 265400 331838
rect 265348 331774 265400 331780
rect 265452 321554 265480 337486
rect 265544 334694 265572 337742
rect 265532 334688 265584 334694
rect 265532 334630 265584 334636
rect 265636 331226 265664 337844
rect 265728 336258 265756 337980
rect 265716 336252 265768 336258
rect 265716 336194 265768 336200
rect 265820 335594 265848 338014
rect 265958 337940 265986 338028
rect 265728 335566 265848 335594
rect 265912 337912 265986 337940
rect 265728 333810 265756 335566
rect 265912 334558 265940 337912
rect 266050 337770 266078 338028
rect 266142 337895 266170 338028
rect 266128 337886 266184 337895
rect 266128 337821 266184 337830
rect 266234 337770 266262 338028
rect 266004 337742 266078 337770
rect 266188 337742 266262 337770
rect 265900 334552 265952 334558
rect 265900 334494 265952 334500
rect 265716 333804 265768 333810
rect 265716 333746 265768 333752
rect 265624 331220 265676 331226
rect 265624 331162 265676 331168
rect 265452 321526 265756 321554
rect 265728 18630 265756 321526
rect 266004 316034 266032 337742
rect 266082 337648 266138 337657
rect 266082 337583 266138 337592
rect 266096 333742 266124 337583
rect 266084 333736 266136 333742
rect 266084 333678 266136 333684
rect 266188 331090 266216 337742
rect 266326 337634 266354 338028
rect 266280 337606 266354 337634
rect 266418 337634 266446 338028
rect 266510 337958 266538 338028
rect 266498 337952 266550 337958
rect 266498 337894 266550 337900
rect 266602 337770 266630 338028
rect 266694 337958 266722 338028
rect 266786 337958 266814 338028
rect 266682 337952 266734 337958
rect 266682 337894 266734 337900
rect 266774 337952 266826 337958
rect 266774 337894 266826 337900
rect 266878 337770 266906 338028
rect 266970 337890 266998 338028
rect 266958 337884 267010 337890
rect 266958 337826 267010 337832
rect 267062 337770 267090 338028
rect 266602 337742 266676 337770
rect 266878 337742 266952 337770
rect 266418 337606 266492 337634
rect 266280 336734 266308 337606
rect 266268 336728 266320 336734
rect 266268 336670 266320 336676
rect 266464 333606 266492 337606
rect 266452 333600 266504 333606
rect 266452 333542 266504 333548
rect 266176 331084 266228 331090
rect 266176 331026 266228 331032
rect 266360 330948 266412 330954
rect 266360 330890 266412 330896
rect 265820 316006 266032 316034
rect 265716 18624 265768 18630
rect 265716 18566 265768 18572
rect 265820 4758 265848 316006
rect 266372 16574 266400 330890
rect 266648 328370 266676 337742
rect 266924 337210 266952 337742
rect 267016 337742 267090 337770
rect 267154 337770 267182 338028
rect 267246 337890 267274 338028
rect 267338 337958 267366 338028
rect 267326 337952 267378 337958
rect 267326 337894 267378 337900
rect 267234 337884 267286 337890
rect 267234 337826 267286 337832
rect 267430 337770 267458 338028
rect 267522 337906 267550 338028
rect 267614 338008 267642 338028
rect 267614 337980 267688 338008
rect 267522 337878 267596 337906
rect 267154 337742 267228 337770
rect 267430 337742 267504 337770
rect 267016 337668 267044 337742
rect 267016 337640 267136 337668
rect 266912 337204 266964 337210
rect 266912 337146 266964 337152
rect 267004 336796 267056 336802
rect 267004 336738 267056 336744
rect 266636 328364 266688 328370
rect 266636 328306 266688 328312
rect 266372 16546 266584 16574
rect 265808 4752 265860 4758
rect 265808 4694 265860 4700
rect 264704 3528 264756 3534
rect 264704 3470 264756 3476
rect 265348 3528 265400 3534
rect 265348 3470 265400 3476
rect 264428 3256 264480 3262
rect 264428 3198 264480 3204
rect 265360 480 265388 3470
rect 266556 480 266584 16546
rect 267016 2990 267044 336738
rect 267108 330886 267136 337640
rect 267096 330880 267148 330886
rect 267096 330822 267148 330828
rect 267200 328302 267228 337742
rect 267476 336530 267504 337742
rect 267464 336524 267516 336530
rect 267464 336466 267516 336472
rect 267280 336184 267332 336190
rect 267280 336126 267332 336132
rect 267188 328296 267240 328302
rect 267188 328238 267240 328244
rect 267292 326534 267320 336126
rect 267568 333402 267596 337878
rect 267556 333396 267608 333402
rect 267556 333338 267608 333344
rect 267660 330750 267688 337980
rect 267798 337770 267826 338028
rect 267890 337890 267918 338028
rect 267878 337884 267930 337890
rect 267878 337826 267930 337832
rect 267982 337770 268010 338028
rect 267798 337742 267872 337770
rect 267740 336320 267792 336326
rect 267740 336262 267792 336268
rect 267752 336054 267780 336262
rect 267740 336048 267792 336054
rect 267740 335990 267792 335996
rect 267740 335368 267792 335374
rect 267740 335310 267792 335316
rect 267648 330744 267700 330750
rect 267648 330686 267700 330692
rect 267752 329866 267780 335310
rect 267740 329860 267792 329866
rect 267740 329802 267792 329808
rect 267844 328234 267872 337742
rect 267936 337742 268010 337770
rect 268074 337770 268102 338028
rect 268166 337890 268194 338028
rect 268154 337884 268206 337890
rect 268154 337826 268206 337832
rect 268258 337770 268286 338028
rect 268350 337958 268378 338028
rect 268338 337952 268390 337958
rect 268338 337894 268390 337900
rect 268442 337822 268470 338028
rect 268430 337816 268482 337822
rect 268074 337742 268148 337770
rect 268258 337742 268332 337770
rect 268430 337758 268482 337764
rect 267936 335374 267964 337742
rect 268016 337544 268068 337550
rect 268016 337486 268068 337492
rect 268028 336410 268056 337486
rect 268120 336666 268148 337742
rect 268108 336660 268160 336666
rect 268108 336602 268160 336608
rect 268028 336382 268148 336410
rect 268120 335510 268148 336382
rect 268108 335504 268160 335510
rect 268108 335446 268160 335452
rect 267924 335368 267976 335374
rect 267924 335310 267976 335316
rect 268304 330546 268332 337742
rect 268534 337668 268562 338028
rect 268626 337958 268654 338028
rect 268718 337963 268746 338028
rect 268614 337952 268666 337958
rect 268614 337894 268666 337900
rect 268704 337954 268760 337963
rect 268704 337889 268760 337898
rect 268810 337890 268838 338028
rect 268902 337929 268930 338028
rect 268888 337920 268944 337929
rect 268798 337884 268850 337890
rect 268994 337890 269022 338028
rect 269086 337958 269114 338028
rect 269074 337952 269126 337958
rect 269074 337894 269126 337900
rect 268888 337855 268944 337864
rect 268982 337884 269034 337890
rect 268798 337826 268850 337832
rect 268982 337826 269034 337832
rect 269026 337784 269082 337793
rect 269178 337770 269206 338028
rect 269270 337929 269298 338028
rect 269362 337958 269390 338028
rect 269350 337952 269402 337958
rect 269256 337920 269312 337929
rect 269350 337894 269402 337900
rect 269256 337855 269312 337864
rect 269454 337770 269482 338028
rect 269638 337929 269666 338028
rect 269624 337920 269680 337929
rect 269624 337855 269680 337864
rect 269730 337770 269758 338028
rect 269178 337742 269252 337770
rect 269454 337742 269528 337770
rect 269026 337719 269082 337728
rect 268534 337640 268700 337668
rect 268566 337512 268622 337521
rect 268566 337447 268622 337456
rect 268384 336320 268436 336326
rect 268384 336262 268436 336268
rect 268292 330540 268344 330546
rect 268292 330482 268344 330488
rect 267832 328228 267884 328234
rect 267832 328170 267884 328176
rect 267280 326528 267332 326534
rect 267280 326470 267332 326476
rect 267740 4888 267792 4894
rect 267740 4830 267792 4836
rect 267004 2984 267056 2990
rect 267004 2926 267056 2932
rect 267752 480 267780 4830
rect 268396 4690 268424 336262
rect 268476 335912 268528 335918
rect 268476 335854 268528 335860
rect 268384 4684 268436 4690
rect 268384 4626 268436 4632
rect 268488 4214 268516 335854
rect 268580 269822 268608 337447
rect 268672 330614 268700 337640
rect 269040 336569 269068 337719
rect 269224 336870 269252 337742
rect 269304 337204 269356 337210
rect 269304 337146 269356 337152
rect 269212 336864 269264 336870
rect 269212 336806 269264 336812
rect 269316 336734 269344 337146
rect 269224 336706 269344 336734
rect 269026 336560 269082 336569
rect 269026 336495 269082 336504
rect 268752 335300 268804 335306
rect 268752 335242 268804 335248
rect 268764 334082 268792 335242
rect 268752 334076 268804 334082
rect 268752 334018 268804 334024
rect 268660 330608 268712 330614
rect 268660 330550 268712 330556
rect 269224 329050 269252 336706
rect 269396 336252 269448 336258
rect 269396 336194 269448 336200
rect 269408 332518 269436 336194
rect 269500 336054 269528 337742
rect 269592 337742 269758 337770
rect 269822 337770 269850 338028
rect 269914 337890 269942 338028
rect 269902 337884 269954 337890
rect 269902 337826 269954 337832
rect 270006 337770 270034 338028
rect 269822 337742 269896 337770
rect 269488 336048 269540 336054
rect 269488 335990 269540 335996
rect 269488 332580 269540 332586
rect 269488 332522 269540 332528
rect 269396 332512 269448 332518
rect 269396 332454 269448 332460
rect 269212 329044 269264 329050
rect 269212 328986 269264 328992
rect 269500 326466 269528 332522
rect 269488 326460 269540 326466
rect 269488 326402 269540 326408
rect 269592 321554 269620 337742
rect 269670 337648 269726 337657
rect 269670 337583 269726 337592
rect 269684 335918 269712 337583
rect 269764 337544 269816 337550
rect 269764 337486 269816 337492
rect 269672 335912 269724 335918
rect 269672 335854 269724 335860
rect 269776 335594 269804 337486
rect 269868 336297 269896 337742
rect 269960 337742 270034 337770
rect 269854 336288 269910 336297
rect 269854 336223 269910 336232
rect 269856 335844 269908 335850
rect 269856 335786 269908 335792
rect 269684 335566 269804 335594
rect 269684 334286 269712 335566
rect 269764 335504 269816 335510
rect 269764 335446 269816 335452
rect 269672 334280 269724 334286
rect 269672 334222 269724 334228
rect 269672 324964 269724 324970
rect 269672 324906 269724 324912
rect 269316 321526 269620 321554
rect 268568 269816 268620 269822
rect 268568 269758 268620 269764
rect 269316 5438 269344 321526
rect 269304 5432 269356 5438
rect 269304 5374 269356 5380
rect 269684 5370 269712 324906
rect 269672 5364 269724 5370
rect 269672 5306 269724 5312
rect 268844 5296 268896 5302
rect 268844 5238 268896 5244
rect 268476 4208 268528 4214
rect 268476 4150 268528 4156
rect 268856 480 268884 5238
rect 269776 2854 269804 335446
rect 269868 331214 269896 335786
rect 269960 335374 269988 337742
rect 270098 337634 270126 338028
rect 270190 337890 270218 338028
rect 270178 337884 270230 337890
rect 270178 337826 270230 337832
rect 270282 337770 270310 338028
rect 270374 337929 270402 338028
rect 270466 337958 270494 338028
rect 270558 337958 270586 338028
rect 270454 337952 270506 337958
rect 270360 337920 270416 337929
rect 270454 337894 270506 337900
rect 270546 337952 270598 337958
rect 270546 337894 270598 337900
rect 270360 337855 270416 337864
rect 270052 337606 270126 337634
rect 270236 337742 270310 337770
rect 270406 337784 270462 337793
rect 269948 335368 270000 335374
rect 269948 335310 270000 335316
rect 269868 331186 269988 331214
rect 269856 326460 269908 326466
rect 269856 326402 269908 326408
rect 269868 4622 269896 326402
rect 269856 4616 269908 4622
rect 269856 4558 269908 4564
rect 269960 4282 269988 331186
rect 270052 324970 270080 337606
rect 270130 337512 270186 337521
rect 270130 337447 270186 337456
rect 270144 333849 270172 337447
rect 270130 333840 270186 333849
rect 270130 333775 270186 333784
rect 270040 324964 270092 324970
rect 270040 324906 270092 324912
rect 270236 5302 270264 337742
rect 270650 337770 270678 338028
rect 270742 337929 270770 338028
rect 270728 337920 270784 337929
rect 270728 337855 270784 337864
rect 270834 337770 270862 338028
rect 270406 337719 270462 337728
rect 270604 337742 270678 337770
rect 270788 337742 270862 337770
rect 270316 337544 270368 337550
rect 270316 337486 270368 337492
rect 270328 336258 270356 337486
rect 270316 336252 270368 336258
rect 270316 336194 270368 336200
rect 270420 336161 270448 337719
rect 270406 336152 270462 336161
rect 270406 336087 270462 336096
rect 270604 336025 270632 337742
rect 270788 337634 270816 337742
rect 270926 337634 270954 338028
rect 271018 337890 271046 338028
rect 271006 337884 271058 337890
rect 271006 337826 271058 337832
rect 271110 337770 271138 338028
rect 271202 337929 271230 338028
rect 271188 337920 271244 337929
rect 271188 337855 271244 337864
rect 271294 337770 271322 338028
rect 271386 337890 271414 338028
rect 271524 338014 271584 338042
rect 271524 337890 271552 338014
rect 271662 337890 271690 338028
rect 271374 337884 271426 337890
rect 271374 337826 271426 337832
rect 271512 337884 271564 337890
rect 271512 337826 271564 337832
rect 271650 337884 271702 337890
rect 271650 337826 271702 337832
rect 271510 337784 271566 337793
rect 271110 337742 271184 337770
rect 271294 337742 271460 337770
rect 270696 337606 270816 337634
rect 270880 337606 270954 337634
rect 271156 337634 271184 337742
rect 271156 337606 271276 337634
rect 270590 336016 270646 336025
rect 270590 335951 270646 335960
rect 270316 335912 270368 335918
rect 270696 335900 270724 337606
rect 270774 337512 270830 337521
rect 270774 337447 270830 337456
rect 270316 335854 270368 335860
rect 270604 335872 270724 335900
rect 270328 333713 270356 335854
rect 270408 335368 270460 335374
rect 270408 335310 270460 335316
rect 270314 333704 270370 333713
rect 270314 333639 270370 333648
rect 270420 330857 270448 335310
rect 270406 330848 270462 330857
rect 270406 330783 270462 330792
rect 270604 330721 270632 335872
rect 270684 335436 270736 335442
rect 270684 335378 270736 335384
rect 270590 330712 270646 330721
rect 270590 330647 270646 330656
rect 270224 5296 270276 5302
rect 270224 5238 270276 5244
rect 270696 5166 270724 335378
rect 270788 333577 270816 337447
rect 270774 333568 270830 333577
rect 270774 333503 270830 333512
rect 270880 232966 270908 337606
rect 271052 332648 271104 332654
rect 271052 332590 271104 332596
rect 270868 232960 270920 232966
rect 270868 232902 270920 232908
rect 271064 177410 271092 332590
rect 271248 234734 271276 337606
rect 271328 337544 271380 337550
rect 271328 337486 271380 337492
rect 271236 234728 271288 234734
rect 271236 234670 271288 234676
rect 271340 233714 271368 337486
rect 271432 334014 271460 337742
rect 271754 337770 271782 338028
rect 271510 337719 271566 337728
rect 271708 337742 271782 337770
rect 271420 334008 271472 334014
rect 271420 333950 271472 333956
rect 271420 326460 271472 326466
rect 271420 326402 271472 326408
rect 271432 233782 271460 326402
rect 271420 233776 271472 233782
rect 271420 233718 271472 233724
rect 271328 233708 271380 233714
rect 271328 233650 271380 233656
rect 271524 232898 271552 337719
rect 271708 326466 271736 337742
rect 271846 337634 271874 338028
rect 271800 337606 271874 337634
rect 271938 337634 271966 338028
rect 272030 337770 272058 338028
rect 272122 337929 272150 338028
rect 272214 337958 272242 338028
rect 272202 337952 272254 337958
rect 272108 337920 272164 337929
rect 272202 337894 272254 337900
rect 272108 337855 272164 337864
rect 272306 337770 272334 338028
rect 272398 337958 272426 338028
rect 272386 337952 272438 337958
rect 272386 337894 272438 337900
rect 272490 337770 272518 338028
rect 272030 337742 272104 337770
rect 272306 337742 272380 337770
rect 271938 337606 272012 337634
rect 271800 335442 271828 337606
rect 271880 337544 271932 337550
rect 271880 337486 271932 337492
rect 271788 335436 271840 335442
rect 271788 335378 271840 335384
rect 271788 334824 271840 334830
rect 271788 334766 271840 334772
rect 271800 333305 271828 334766
rect 271786 333296 271842 333305
rect 271786 333231 271842 333240
rect 271696 326460 271748 326466
rect 271696 326402 271748 326408
rect 271892 233850 271920 337486
rect 271984 335986 272012 337606
rect 271972 335980 272024 335986
rect 271972 335922 272024 335928
rect 271972 335572 272024 335578
rect 271972 335514 272024 335520
rect 271984 334830 272012 335514
rect 272076 335510 272104 337742
rect 272064 335504 272116 335510
rect 272064 335446 272116 335452
rect 271972 334824 272024 334830
rect 271972 334766 272024 334772
rect 272156 334416 272208 334422
rect 272156 334358 272208 334364
rect 272168 316034 272196 334358
rect 272352 332654 272380 337742
rect 272444 337742 272518 337770
rect 272444 333441 272472 337742
rect 272582 337634 272610 338028
rect 272674 337770 272702 338028
rect 272766 337958 272794 338028
rect 272754 337952 272806 337958
rect 272754 337894 272806 337900
rect 272858 337890 272886 338028
rect 272950 337963 272978 338028
rect 272936 337954 272992 337963
rect 272846 337884 272898 337890
rect 272936 337889 272992 337898
rect 272846 337826 272898 337832
rect 272890 337784 272946 337793
rect 272674 337742 272748 337770
rect 272582 337606 272656 337634
rect 272524 335980 272576 335986
rect 272524 335922 272576 335928
rect 272536 334762 272564 335922
rect 272524 334756 272576 334762
rect 272524 334698 272576 334704
rect 272430 333432 272486 333441
rect 272430 333367 272486 333376
rect 272340 332648 272392 332654
rect 272340 332590 272392 332596
rect 272628 323626 272656 337606
rect 272720 334150 272748 337742
rect 273042 337770 273070 338028
rect 273134 337895 273162 338028
rect 273120 337886 273176 337895
rect 273226 337872 273254 338028
rect 273318 338008 273346 338028
rect 273456 338014 273516 338042
rect 273318 337980 273392 338008
rect 273226 337844 273300 337872
rect 273120 337821 273176 337830
rect 273272 337770 273300 337844
rect 272890 337719 272946 337728
rect 272996 337742 273070 337770
rect 273180 337742 273300 337770
rect 272800 335504 272852 335510
rect 272800 335446 272852 335452
rect 272708 334144 272760 334150
rect 272708 334086 272760 334092
rect 272812 331214 272840 335446
rect 272904 334422 272932 337719
rect 272892 334416 272944 334422
rect 272892 334358 272944 334364
rect 272892 332648 272944 332654
rect 272892 332590 272944 332596
rect 272720 331186 272840 331214
rect 272720 326466 272748 331186
rect 272708 326460 272760 326466
rect 272708 326402 272760 326408
rect 272628 323598 272840 323626
rect 272708 322516 272760 322522
rect 272708 322458 272760 322464
rect 272076 316006 272196 316034
rect 271880 233844 271932 233850
rect 271880 233786 271932 233792
rect 271512 232892 271564 232898
rect 271512 232834 271564 232840
rect 272076 232830 272104 316006
rect 272720 239873 272748 322458
rect 272706 239864 272762 239873
rect 272706 239799 272762 239808
rect 272812 234870 272840 323598
rect 272800 234864 272852 234870
rect 272800 234806 272852 234812
rect 272904 234802 272932 332590
rect 272996 332450 273024 337742
rect 273074 337648 273130 337657
rect 273074 337583 273130 337592
rect 272984 332444 273036 332450
rect 272984 332386 273036 332392
rect 273088 316034 273116 337583
rect 273180 336433 273208 337742
rect 273166 336424 273222 336433
rect 273166 336359 273222 336368
rect 273364 329934 273392 337980
rect 273456 335209 273484 338014
rect 273594 337906 273622 338028
rect 273548 337878 273622 337906
rect 273548 337210 273576 337878
rect 273686 337804 273714 338028
rect 273778 337890 273806 338028
rect 273766 337884 273818 337890
rect 273766 337826 273818 337832
rect 273640 337776 273714 337804
rect 273536 337204 273588 337210
rect 273536 337146 273588 337152
rect 273442 335200 273498 335209
rect 273442 335135 273498 335144
rect 273640 332466 273668 337776
rect 273870 337770 273898 338028
rect 273962 337890 273990 338028
rect 273950 337884 274002 337890
rect 273950 337826 274002 337832
rect 274054 337770 274082 338028
rect 274146 337890 274174 338028
rect 274238 337958 274266 338028
rect 274226 337952 274278 337958
rect 274226 337894 274278 337900
rect 274134 337884 274186 337890
rect 274134 337826 274186 337832
rect 274330 337770 274358 338028
rect 274422 337804 274450 338028
rect 274514 337929 274542 338028
rect 274500 337920 274556 337929
rect 274500 337855 274556 337864
rect 274422 337776 274496 337804
rect 273870 337742 273944 337770
rect 273916 335850 273944 337742
rect 274008 337742 274082 337770
rect 274284 337742 274358 337770
rect 273904 335844 273956 335850
rect 273904 335786 273956 335792
rect 274008 335730 274036 337742
rect 274284 336954 274312 337742
rect 273824 335702 274036 335730
rect 274100 336926 274312 336954
rect 273720 335028 273772 335034
rect 273720 334970 273772 334976
rect 273456 332438 273668 332466
rect 273352 329928 273404 329934
rect 273352 329870 273404 329876
rect 273456 328454 273484 332438
rect 273732 330698 273760 334970
rect 272996 316006 273116 316034
rect 273272 328426 273484 328454
rect 273548 330670 273760 330698
rect 272892 234796 272944 234802
rect 272892 234738 272944 234744
rect 272996 234598 273024 316006
rect 273272 234938 273300 328426
rect 273548 316034 273576 330670
rect 273824 330562 273852 335702
rect 273904 335504 273956 335510
rect 273904 335446 273956 335452
rect 273364 316006 273576 316034
rect 273640 330534 273852 330562
rect 273916 330562 273944 335446
rect 273916 330534 274036 330562
rect 273260 234932 273312 234938
rect 273260 234874 273312 234880
rect 272984 234592 273036 234598
rect 272984 234534 273036 234540
rect 273364 234326 273392 316006
rect 273640 234394 273668 330534
rect 273720 329928 273772 329934
rect 273720 329870 273772 329876
rect 273732 239465 273760 329870
rect 273904 329792 273956 329798
rect 273904 329734 273956 329740
rect 273718 239456 273774 239465
rect 273718 239391 273774 239400
rect 273628 234388 273680 234394
rect 273628 234330 273680 234336
rect 273352 234320 273404 234326
rect 273352 234262 273404 234268
rect 272064 232824 272116 232830
rect 272064 232766 272116 232772
rect 271052 177404 271104 177410
rect 271052 177346 271104 177352
rect 273260 93152 273312 93158
rect 273260 93094 273312 93100
rect 270592 5160 270644 5166
rect 270592 5102 270644 5108
rect 270684 5160 270736 5166
rect 270684 5102 270736 5108
rect 269948 4276 270000 4282
rect 269948 4218 270000 4224
rect 270604 4214 270632 5102
rect 272432 5024 272484 5030
rect 272432 4966 272484 4972
rect 270592 4208 270644 4214
rect 270592 4150 270644 4156
rect 271236 4208 271288 4214
rect 271236 4150 271288 4156
rect 270040 3256 270092 3262
rect 270040 3198 270092 3204
rect 269764 2848 269816 2854
rect 269764 2790 269816 2796
rect 270052 480 270080 3198
rect 271248 480 271276 4150
rect 272444 480 272472 4966
rect 273272 490 273300 93094
rect 273916 5030 273944 329734
rect 274008 235210 274036 330534
rect 273996 235204 274048 235210
rect 273996 235146 274048 235152
rect 274100 235074 274128 336926
rect 274272 336796 274324 336802
rect 274272 336738 274324 336744
rect 274180 335844 274232 335850
rect 274180 335786 274232 335792
rect 274192 332178 274220 335786
rect 274180 332172 274232 332178
rect 274180 332114 274232 332120
rect 274180 332036 274232 332042
rect 274180 331978 274232 331984
rect 274088 235068 274140 235074
rect 274088 235010 274140 235016
rect 274192 235006 274220 331978
rect 274180 235000 274232 235006
rect 274180 234942 274232 234948
rect 274284 234462 274312 336738
rect 274468 335578 274496 337776
rect 274606 337770 274634 338028
rect 274560 337742 274634 337770
rect 274456 335572 274508 335578
rect 274456 335514 274508 335520
rect 274560 335510 274588 337742
rect 274698 337634 274726 338028
rect 274790 337770 274818 338028
rect 274882 337958 274910 338028
rect 274974 337963 275002 338028
rect 274870 337952 274922 337958
rect 274870 337894 274922 337900
rect 274960 337954 275016 337963
rect 274960 337889 275016 337898
rect 275066 337770 275094 338028
rect 275158 337958 275186 338028
rect 275146 337952 275198 337958
rect 275146 337894 275198 337900
rect 275250 337770 275278 338028
rect 274790 337742 274864 337770
rect 275066 337742 275140 337770
rect 274698 337606 274772 337634
rect 274638 337512 274694 337521
rect 274638 337447 274694 337456
rect 274548 335504 274600 335510
rect 274548 335446 274600 335452
rect 274362 335200 274418 335209
rect 274362 335135 274418 335144
rect 274376 234530 274404 335135
rect 274652 334626 274680 337447
rect 274744 336802 274772 337606
rect 274732 336796 274784 336802
rect 274732 336738 274784 336744
rect 274732 335912 274784 335918
rect 274732 335854 274784 335860
rect 274744 335374 274772 335854
rect 274836 335753 274864 337742
rect 275112 336870 275140 337742
rect 275204 337742 275278 337770
rect 275388 338014 275448 338042
rect 275100 336864 275152 336870
rect 275100 336806 275152 336812
rect 274822 335744 274878 335753
rect 274822 335679 274878 335688
rect 274824 335572 274876 335578
rect 274824 335514 274876 335520
rect 274732 335368 274784 335374
rect 274732 335310 274784 335316
rect 274640 334620 274692 334626
rect 274640 334562 274692 334568
rect 274836 235890 274864 335514
rect 274916 335368 274968 335374
rect 274916 335310 274968 335316
rect 274824 235884 274876 235890
rect 274824 235826 274876 235832
rect 274364 234524 274416 234530
rect 274364 234466 274416 234472
rect 274272 234456 274324 234462
rect 274272 234398 274324 234404
rect 274928 231198 274956 335310
rect 275204 328454 275232 337742
rect 275284 337544 275336 337550
rect 275284 337486 275336 337492
rect 275020 328426 275232 328454
rect 275020 234190 275048 328426
rect 275296 316034 275324 337486
rect 275388 336938 275416 338014
rect 275526 337940 275554 338028
rect 275480 337912 275554 337940
rect 275376 336932 275428 336938
rect 275376 336874 275428 336880
rect 275480 335578 275508 337912
rect 275618 337872 275646 338028
rect 275572 337844 275646 337872
rect 275572 336734 275600 337844
rect 275710 337668 275738 338028
rect 275802 337890 275830 338028
rect 275894 337963 275922 338028
rect 275880 337954 275936 337963
rect 275986 337958 276014 338028
rect 276078 337963 276106 338028
rect 275790 337884 275842 337890
rect 275880 337889 275936 337898
rect 275974 337952 276026 337958
rect 275974 337894 276026 337900
rect 276064 337954 276120 337963
rect 276170 337958 276198 338028
rect 276262 337963 276290 338028
rect 276064 337889 276120 337898
rect 276158 337952 276210 337958
rect 276158 337894 276210 337900
rect 276248 337954 276304 337963
rect 276248 337889 276304 337898
rect 276354 337890 276382 338028
rect 276446 337958 276474 338028
rect 276434 337952 276486 337958
rect 276434 337894 276486 337900
rect 275790 337826 275842 337832
rect 276342 337884 276394 337890
rect 276342 337826 276394 337832
rect 275926 337784 275982 337793
rect 275926 337719 275982 337728
rect 276202 337784 276258 337793
rect 276202 337719 276258 337728
rect 275664 337640 275738 337668
rect 275664 337346 275692 337640
rect 275744 337544 275796 337550
rect 275744 337486 275796 337492
rect 275834 337512 275890 337521
rect 275652 337340 275704 337346
rect 275652 337282 275704 337288
rect 275572 336706 275692 336734
rect 275468 335572 275520 335578
rect 275468 335514 275520 335520
rect 275468 335368 275520 335374
rect 275468 335310 275520 335316
rect 275560 335368 275612 335374
rect 275560 335310 275612 335316
rect 275376 334280 275428 334286
rect 275376 334222 275428 334228
rect 275204 316006 275324 316034
rect 275204 239737 275232 316006
rect 275190 239728 275246 239737
rect 275190 239663 275246 239672
rect 275388 235958 275416 334222
rect 275376 235952 275428 235958
rect 275376 235894 275428 235900
rect 275480 235142 275508 335310
rect 275572 235822 275600 335310
rect 275560 235816 275612 235822
rect 275560 235758 275612 235764
rect 275468 235136 275520 235142
rect 275468 235078 275520 235084
rect 275008 234184 275060 234190
rect 275008 234126 275060 234132
rect 275664 234122 275692 336706
rect 275756 335374 275784 337486
rect 275834 337447 275890 337456
rect 275744 335368 275796 335374
rect 275744 335310 275796 335316
rect 275848 316034 275876 337447
rect 275940 335918 275968 337719
rect 275928 335912 275980 335918
rect 275928 335854 275980 335860
rect 276216 335354 276244 337719
rect 276538 337668 276566 338028
rect 276630 337770 276658 338028
rect 276722 337963 276750 338028
rect 276708 337954 276764 337963
rect 276708 337889 276764 337898
rect 276630 337742 276704 337770
rect 276294 337648 276350 337657
rect 276294 337583 276350 337592
rect 276492 337640 276566 337668
rect 276308 337006 276336 337583
rect 276388 337544 276440 337550
rect 276492 337532 276520 337640
rect 276440 337504 276520 337532
rect 276388 337486 276440 337492
rect 276296 337000 276348 337006
rect 276296 336942 276348 336948
rect 276216 335326 276336 335354
rect 276308 334558 276336 335326
rect 276296 334552 276348 334558
rect 276296 334494 276348 334500
rect 276020 334144 276072 334150
rect 276020 334086 276072 334092
rect 276032 325694 276060 334086
rect 276480 332648 276532 332654
rect 276480 332590 276532 332596
rect 276388 332444 276440 332450
rect 276388 332386 276440 332392
rect 276296 329792 276348 329798
rect 276296 329734 276348 329740
rect 276032 325666 276152 325694
rect 275756 316006 275876 316034
rect 275756 234258 275784 316006
rect 275744 234252 275796 234258
rect 275744 234194 275796 234200
rect 275652 234116 275704 234122
rect 275652 234058 275704 234064
rect 276020 232552 276072 232558
rect 276020 232494 276072 232500
rect 274916 231192 274968 231198
rect 274916 231134 274968 231140
rect 276032 16574 276060 232494
rect 276124 231130 276152 325666
rect 276112 231124 276164 231130
rect 276112 231066 276164 231072
rect 276308 177342 276336 329734
rect 276400 239601 276428 332386
rect 276386 239592 276442 239601
rect 276386 239527 276442 239536
rect 276492 235618 276520 332590
rect 276572 332444 276624 332450
rect 276572 332386 276624 332392
rect 276584 235686 276612 332386
rect 276676 235754 276704 337742
rect 276814 337668 276842 338028
rect 276906 337770 276934 338028
rect 276998 337963 277026 338028
rect 276984 337954 277040 337963
rect 277090 337958 277118 338028
rect 277182 338008 277210 338028
rect 277320 338014 277380 338042
rect 277182 337980 277256 338008
rect 276984 337889 277040 337898
rect 277078 337952 277130 337958
rect 277078 337894 277130 337900
rect 277122 337784 277178 337793
rect 276906 337742 276980 337770
rect 276814 337640 276888 337668
rect 276756 337000 276808 337006
rect 276756 336942 276808 336948
rect 276664 235748 276716 235754
rect 276664 235690 276716 235696
rect 276572 235680 276624 235686
rect 276572 235622 276624 235628
rect 276480 235612 276532 235618
rect 276480 235554 276532 235560
rect 276768 235550 276796 336942
rect 276860 336734 276888 337640
rect 276952 337006 276980 337742
rect 277122 337719 277178 337728
rect 277136 337550 277164 337719
rect 277124 337544 277176 337550
rect 277124 337486 277176 337492
rect 277122 337376 277178 337385
rect 277122 337311 277178 337320
rect 276940 337000 276992 337006
rect 276940 336942 276992 336948
rect 276860 336706 276980 336734
rect 276952 334422 276980 336706
rect 277032 334892 277084 334898
rect 277032 334834 277084 334840
rect 276940 334416 276992 334422
rect 276940 334358 276992 334364
rect 276940 332240 276992 332246
rect 276940 332182 276992 332188
rect 276848 332104 276900 332110
rect 276848 332046 276900 332052
rect 276756 235544 276808 235550
rect 276756 235486 276808 235492
rect 276860 235482 276888 332046
rect 276848 235476 276900 235482
rect 276848 235418 276900 235424
rect 276952 234054 276980 332182
rect 276940 234048 276992 234054
rect 276940 233990 276992 233996
rect 277044 233986 277072 334834
rect 277032 233980 277084 233986
rect 277032 233922 277084 233928
rect 277136 232762 277164 337311
rect 277228 332654 277256 337980
rect 277216 332648 277268 332654
rect 277216 332590 277268 332596
rect 277320 329798 277348 338014
rect 277458 337770 277486 338028
rect 277412 337742 277486 337770
rect 277412 336870 277440 337742
rect 277550 337634 277578 338028
rect 277642 337770 277670 338028
rect 277734 337890 277762 338028
rect 277722 337884 277774 337890
rect 277722 337826 277774 337832
rect 277826 337770 277854 338028
rect 277918 337929 277946 338028
rect 277904 337920 277960 337929
rect 278010 337890 278038 338028
rect 278102 337958 278130 338028
rect 278090 337952 278142 337958
rect 278090 337894 278142 337900
rect 277904 337855 277960 337864
rect 277998 337884 278050 337890
rect 277998 337826 278050 337832
rect 277642 337742 277716 337770
rect 277550 337606 277624 337634
rect 277400 336864 277452 336870
rect 277400 336806 277452 336812
rect 277490 336424 277546 336433
rect 277490 336359 277546 336368
rect 277400 335912 277452 335918
rect 277504 335889 277532 336359
rect 277400 335854 277452 335860
rect 277490 335880 277546 335889
rect 277412 335730 277440 335854
rect 277490 335815 277546 335824
rect 277412 335702 277532 335730
rect 277400 335368 277452 335374
rect 277400 335310 277452 335316
rect 277308 329792 277360 329798
rect 277308 329734 277360 329740
rect 277412 235414 277440 335310
rect 277504 325694 277532 335702
rect 277596 329730 277624 337606
rect 277688 329934 277716 337742
rect 277780 337742 277854 337770
rect 277950 337784 278006 337793
rect 277780 335374 277808 337742
rect 278194 337770 278222 338028
rect 278286 337929 278314 338028
rect 278378 337958 278406 338028
rect 278470 337963 278498 338028
rect 278366 337952 278418 337958
rect 278272 337920 278328 337929
rect 278366 337894 278418 337900
rect 278456 337954 278512 337963
rect 278456 337889 278512 337898
rect 278272 337855 278328 337864
rect 278562 337770 278590 338028
rect 278654 337804 278682 338028
rect 278746 337958 278774 338028
rect 278838 337963 278866 338028
rect 278734 337952 278786 337958
rect 278734 337894 278786 337900
rect 278824 337954 278880 337963
rect 278824 337889 278880 337898
rect 278930 337822 278958 338028
rect 279022 337963 279050 338028
rect 279008 337954 279064 337963
rect 279114 337958 279142 338028
rect 279252 338014 279312 338042
rect 279008 337889 279064 337898
rect 279102 337952 279154 337958
rect 279102 337894 279154 337900
rect 278918 337816 278970 337822
rect 278654 337776 278774 337804
rect 277950 337719 278006 337728
rect 278148 337742 278222 337770
rect 278516 337742 278590 337770
rect 277858 337648 277914 337657
rect 277858 337583 277914 337592
rect 277768 335368 277820 335374
rect 277768 335310 277820 335316
rect 277676 329928 277728 329934
rect 277676 329870 277728 329876
rect 277584 329724 277636 329730
rect 277584 329666 277636 329672
rect 277872 328454 277900 337583
rect 277964 335578 277992 337719
rect 278148 337634 278176 337742
rect 278148 337606 278268 337634
rect 278136 337340 278188 337346
rect 278136 337282 278188 337288
rect 277952 335572 278004 335578
rect 277952 335514 278004 335520
rect 277952 335368 278004 335374
rect 277952 335310 278004 335316
rect 277964 334801 277992 335310
rect 277950 334792 278006 334801
rect 277950 334727 278006 334736
rect 278044 334008 278096 334014
rect 278044 333950 278096 333956
rect 277952 329724 278004 329730
rect 277952 329666 278004 329672
rect 277780 328426 277900 328454
rect 277504 325666 277624 325694
rect 277400 235408 277452 235414
rect 277400 235350 277452 235356
rect 277124 232756 277176 232762
rect 277124 232698 277176 232704
rect 276296 177336 276348 177342
rect 276296 177278 276348 177284
rect 276032 16546 276704 16574
rect 273904 5024 273956 5030
rect 273904 4966 273956 4972
rect 276020 4888 276072 4894
rect 276020 4830 276072 4836
rect 274824 4412 274876 4418
rect 274824 4354 274876 4360
rect 273456 598 273668 626
rect 273456 490 273484 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 462 273484 490
rect 273640 480 273668 598
rect 274836 480 274864 4354
rect 276032 480 276060 4830
rect 276676 490 276704 16546
rect 277596 4865 277624 325666
rect 277780 316034 277808 328426
rect 277688 316006 277808 316034
rect 277688 175982 277716 316006
rect 277964 235278 277992 329666
rect 277952 235272 278004 235278
rect 277952 235214 278004 235220
rect 277676 175976 277728 175982
rect 277676 175918 277728 175924
rect 277582 4856 277638 4865
rect 277582 4791 277638 4800
rect 278056 3126 278084 333950
rect 278148 235346 278176 337282
rect 278240 335442 278268 337606
rect 278320 337544 278372 337550
rect 278320 337486 278372 337492
rect 278228 335436 278280 335442
rect 278228 335378 278280 335384
rect 278332 335322 278360 337486
rect 278516 335918 278544 337742
rect 278746 337634 278774 337776
rect 278918 337758 278970 337764
rect 278962 337648 279018 337657
rect 278746 337606 278820 337634
rect 278596 337136 278648 337142
rect 278596 337078 278648 337084
rect 278504 335912 278556 335918
rect 278504 335854 278556 335860
rect 278504 335572 278556 335578
rect 278504 335514 278556 335520
rect 278412 335436 278464 335442
rect 278412 335378 278464 335384
rect 278240 335294 278360 335322
rect 278136 235340 278188 235346
rect 278136 235282 278188 235288
rect 278240 233918 278268 335294
rect 278320 329928 278372 329934
rect 278320 329870 278372 329876
rect 278228 233912 278280 233918
rect 278228 233854 278280 233860
rect 278332 232694 278360 329870
rect 278320 232688 278372 232694
rect 278320 232630 278372 232636
rect 278424 232558 278452 335378
rect 278516 232626 278544 335514
rect 278608 334150 278636 337078
rect 278596 334144 278648 334150
rect 278596 334086 278648 334092
rect 278792 331294 278820 337606
rect 278962 337583 279018 337592
rect 278976 337346 279004 337583
rect 278964 337340 279016 337346
rect 278964 337282 279016 337288
rect 279148 337068 279200 337074
rect 279148 337010 279200 337016
rect 278780 331288 278832 331294
rect 278780 331230 278832 331236
rect 279160 329798 279188 337010
rect 279252 332110 279280 338014
rect 279390 337770 279418 338028
rect 279344 337742 279418 337770
rect 279482 337770 279510 338028
rect 279574 337890 279602 338028
rect 279562 337884 279614 337890
rect 279562 337826 279614 337832
rect 279482 337742 279556 337770
rect 279344 337074 279372 337742
rect 279422 337648 279478 337657
rect 279422 337583 279478 337592
rect 279332 337068 279384 337074
rect 279332 337010 279384 337016
rect 279436 336274 279464 337583
rect 279528 337142 279556 337742
rect 279666 337634 279694 338028
rect 279758 337770 279786 338028
rect 279850 337929 279878 338028
rect 279836 337920 279892 337929
rect 279836 337855 279892 337864
rect 279942 337770 279970 338028
rect 279758 337742 279832 337770
rect 279666 337606 279740 337634
rect 279712 337362 279740 337606
rect 279804 337532 279832 337742
rect 279896 337742 279970 337770
rect 280034 337770 280062 338028
rect 280126 337890 280154 338028
rect 280218 337890 280246 338028
rect 280114 337884 280166 337890
rect 280114 337826 280166 337832
rect 280206 337884 280258 337890
rect 280206 337826 280258 337832
rect 280310 337804 280338 338028
rect 280402 337963 280430 338028
rect 280388 337954 280444 337963
rect 280388 337889 280444 337898
rect 280310 337776 280384 337804
rect 280034 337742 280108 337770
rect 279896 337634 279924 337742
rect 279896 337606 280016 337634
rect 279804 337504 279924 337532
rect 279712 337334 279832 337362
rect 279516 337136 279568 337142
rect 279516 337078 279568 337084
rect 279608 336864 279660 336870
rect 279608 336806 279660 336812
rect 279516 336796 279568 336802
rect 279516 336738 279568 336744
rect 279344 336246 279464 336274
rect 279240 332104 279292 332110
rect 279240 332046 279292 332052
rect 279344 332042 279372 336246
rect 279424 336116 279476 336122
rect 279424 336058 279476 336064
rect 279332 332036 279384 332042
rect 279332 331978 279384 331984
rect 279240 331968 279292 331974
rect 279240 331910 279292 331916
rect 279252 330585 279280 331910
rect 279238 330576 279294 330585
rect 279238 330511 279294 330520
rect 279148 329792 279200 329798
rect 279148 329734 279200 329740
rect 278504 232620 278556 232626
rect 278504 232562 278556 232568
rect 278412 232552 278464 232558
rect 278412 232494 278464 232500
rect 279436 6914 279464 336058
rect 279344 6886 279464 6914
rect 278320 5500 278372 5506
rect 278320 5442 278372 5448
rect 278044 3120 278096 3126
rect 278044 3062 278096 3068
rect 276952 598 277164 626
rect 276952 490 276980 598
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 462 276980 490
rect 277136 480 277164 598
rect 278332 480 278360 5442
rect 279344 3369 279372 6886
rect 279528 5930 279556 336738
rect 279620 332654 279648 336806
rect 279608 332648 279660 332654
rect 279608 332590 279660 332596
rect 279608 332172 279660 332178
rect 279608 332114 279660 332120
rect 279620 6066 279648 332114
rect 279804 329662 279832 337334
rect 279896 335345 279924 337504
rect 279882 335336 279938 335345
rect 279882 335271 279938 335280
rect 279988 329730 280016 337606
rect 280080 335209 280108 337742
rect 280356 335918 280384 337776
rect 280494 337770 280522 338028
rect 280586 337890 280614 338028
rect 280678 337895 280706 338028
rect 280574 337884 280626 337890
rect 280574 337826 280626 337832
rect 280664 337886 280720 337895
rect 280664 337821 280720 337830
rect 280770 337770 280798 338028
rect 280862 337890 280890 338028
rect 280850 337884 280902 337890
rect 280850 337826 280902 337832
rect 280954 337770 280982 338028
rect 281046 337906 281074 338028
rect 281184 338014 281244 338042
rect 281046 337878 281120 337906
rect 280494 337742 280568 337770
rect 280434 337648 280490 337657
rect 280434 337583 280490 337592
rect 280344 335912 280396 335918
rect 280344 335854 280396 335860
rect 280066 335200 280122 335209
rect 280066 335135 280122 335144
rect 280448 332489 280476 337583
rect 280434 332480 280490 332489
rect 280434 332415 280490 332424
rect 280160 331900 280212 331906
rect 280160 331842 280212 331848
rect 279976 329724 280028 329730
rect 279976 329666 280028 329672
rect 279700 329656 279752 329662
rect 279700 329598 279752 329604
rect 279792 329656 279844 329662
rect 279792 329598 279844 329604
rect 279712 16574 279740 329598
rect 280172 16574 280200 331842
rect 280540 329458 280568 337742
rect 280632 337742 280798 337770
rect 280908 337742 280982 337770
rect 280528 329452 280580 329458
rect 280528 329394 280580 329400
rect 280632 328778 280660 337742
rect 280908 335866 280936 337742
rect 280724 335838 280936 335866
rect 280724 332353 280752 335838
rect 280804 335776 280856 335782
rect 280804 335718 280856 335724
rect 280894 335744 280950 335753
rect 280710 332344 280766 332353
rect 280710 332279 280766 332288
rect 280620 328772 280672 328778
rect 280620 328714 280672 328720
rect 279712 16546 279832 16574
rect 280172 16546 280752 16574
rect 279620 6038 279740 6066
rect 279528 5902 279648 5930
rect 279620 4962 279648 5902
rect 279516 4956 279568 4962
rect 279516 4898 279568 4904
rect 279608 4956 279660 4962
rect 279608 4898 279660 4904
rect 279330 3360 279386 3369
rect 279330 3295 279386 3304
rect 279528 480 279556 4898
rect 279712 4146 279740 6038
rect 279700 4140 279752 4146
rect 279700 4082 279752 4088
rect 279804 3194 279832 16546
rect 279792 3188 279844 3194
rect 279792 3130 279844 3136
rect 280724 480 280752 16546
rect 280816 4078 280844 335718
rect 280894 335679 280950 335688
rect 280804 4072 280856 4078
rect 280804 4014 280856 4020
rect 280908 3874 280936 335679
rect 280988 334620 281040 334626
rect 280988 334562 281040 334568
rect 281000 3942 281028 334562
rect 281092 329390 281120 337878
rect 281184 335073 281212 338014
rect 281322 337958 281350 338028
rect 281310 337952 281362 337958
rect 281310 337894 281362 337900
rect 281414 337895 281442 338028
rect 281400 337886 281456 337895
rect 281400 337821 281456 337830
rect 281506 337770 281534 338028
rect 281460 337742 281534 337770
rect 281598 337770 281626 338028
rect 281690 337958 281718 338028
rect 281678 337952 281730 337958
rect 281678 337894 281730 337900
rect 281782 337770 281810 338028
rect 281874 337958 281902 338028
rect 281862 337952 281914 337958
rect 281862 337894 281914 337900
rect 281966 337770 281994 338028
rect 281598 337742 281672 337770
rect 281782 337742 281856 337770
rect 281262 337648 281318 337657
rect 281262 337583 281318 337592
rect 281170 335064 281226 335073
rect 281170 334999 281226 335008
rect 281080 329384 281132 329390
rect 281080 329326 281132 329332
rect 281276 329322 281304 337583
rect 281356 335504 281408 335510
rect 281356 335446 281408 335452
rect 281368 332217 281396 335446
rect 281460 334937 281488 337742
rect 281446 334928 281502 334937
rect 281446 334863 281502 334872
rect 281354 332208 281410 332217
rect 281354 332143 281410 332152
rect 281644 332081 281672 337742
rect 281828 336002 281856 337742
rect 281920 337742 281994 337770
rect 281920 336138 281948 337742
rect 282058 337532 282086 338028
rect 282150 337958 282178 338028
rect 282138 337952 282190 337958
rect 282138 337894 282190 337900
rect 282242 337770 282270 338028
rect 282334 337929 282362 338028
rect 282426 337958 282454 338028
rect 282518 337958 282546 338028
rect 282610 337963 282638 338028
rect 282414 337952 282466 337958
rect 282320 337920 282376 337929
rect 282414 337894 282466 337900
rect 282506 337952 282558 337958
rect 282506 337894 282558 337900
rect 282596 337954 282652 337963
rect 282596 337889 282652 337898
rect 282320 337855 282376 337864
rect 282550 337784 282606 337793
rect 282242 337742 282316 337770
rect 282288 337634 282316 337742
rect 282702 337770 282730 338028
rect 282794 337804 282822 338028
rect 282886 337872 282914 338028
rect 282978 337940 283006 338028
rect 282978 337912 283052 337940
rect 282886 337844 282960 337872
rect 282794 337776 282868 337804
rect 282550 337719 282606 337728
rect 282656 337742 282730 337770
rect 282288 337606 282500 337634
rect 282368 337544 282420 337550
rect 282058 337504 282132 337532
rect 281920 336110 282040 336138
rect 281828 335974 281948 336002
rect 281816 335572 281868 335578
rect 281816 335514 281868 335520
rect 281630 332072 281686 332081
rect 281630 332007 281686 332016
rect 281264 329316 281316 329322
rect 281264 329258 281316 329264
rect 281080 329112 281132 329118
rect 281080 329054 281132 329060
rect 280988 3936 281040 3942
rect 280988 3878 281040 3884
rect 280896 3868 280948 3874
rect 280896 3810 280948 3816
rect 281092 3262 281120 329054
rect 281828 236706 281856 335514
rect 281920 334801 281948 335974
rect 282012 335782 282040 336110
rect 282000 335776 282052 335782
rect 282104 335764 282132 337504
rect 282274 337512 282330 337521
rect 282368 337486 282420 337492
rect 282274 337447 282330 337456
rect 282104 335736 282224 335764
rect 282000 335718 282052 335724
rect 282000 335504 282052 335510
rect 282000 335446 282052 335452
rect 282092 335504 282144 335510
rect 282092 335446 282144 335452
rect 281906 334792 281962 334801
rect 281906 334727 281962 334736
rect 282012 331945 282040 335446
rect 281998 331936 282054 331945
rect 281998 331871 282054 331880
rect 282104 236842 282132 335446
rect 282196 334665 282224 335736
rect 282288 335481 282316 337447
rect 282380 336705 282408 337486
rect 282366 336696 282422 336705
rect 282366 336631 282422 336640
rect 282274 335472 282330 335481
rect 282274 335407 282330 335416
rect 282276 335300 282328 335306
rect 282276 335242 282328 335248
rect 282182 334656 282238 334665
rect 282182 334591 282238 334600
rect 282288 334540 282316 335242
rect 282196 334512 282316 334540
rect 282092 236836 282144 236842
rect 282092 236778 282144 236784
rect 281816 236700 281868 236706
rect 281816 236642 281868 236648
rect 281908 5092 281960 5098
rect 281908 5034 281960 5040
rect 281080 3256 281132 3262
rect 281080 3198 281132 3204
rect 281920 480 281948 5034
rect 282196 3330 282224 334512
rect 282276 334212 282328 334218
rect 282276 334154 282328 334160
rect 282368 334212 282420 334218
rect 282368 334154 282420 334160
rect 282184 3324 282236 3330
rect 282184 3266 282236 3272
rect 282288 3058 282316 334154
rect 282380 334082 282408 334154
rect 282368 334076 282420 334082
rect 282368 334018 282420 334024
rect 282368 332172 282420 332178
rect 282368 332114 282420 332120
rect 282380 331809 282408 332114
rect 282366 331800 282422 331809
rect 282366 331735 282422 331744
rect 282472 329118 282500 337606
rect 282564 335578 282592 337719
rect 282552 335572 282604 335578
rect 282552 335514 282604 335520
rect 282656 335510 282684 337742
rect 282840 337634 282868 337776
rect 282748 337606 282868 337634
rect 282644 335504 282696 335510
rect 282644 335446 282696 335452
rect 282552 335300 282604 335306
rect 282552 335242 282604 335248
rect 282460 329112 282512 329118
rect 282460 329054 282512 329060
rect 282564 328030 282592 335242
rect 282644 335232 282696 335238
rect 282644 335174 282696 335180
rect 282656 334121 282684 335174
rect 282642 334112 282698 334121
rect 282642 334047 282698 334056
rect 282552 328024 282604 328030
rect 282552 327966 282604 327972
rect 282748 316034 282776 337606
rect 282932 337550 282960 337844
rect 282920 337544 282972 337550
rect 282920 337486 282972 337492
rect 282920 337068 282972 337074
rect 282920 337010 282972 337016
rect 282932 336569 282960 337010
rect 283024 336938 283052 337912
rect 283162 337770 283190 338028
rect 283254 337963 283282 338028
rect 283240 337954 283296 337963
rect 283240 337889 283296 337898
rect 283346 337770 283374 338028
rect 283438 337929 283466 338028
rect 283424 337920 283480 337929
rect 283424 337855 283480 337864
rect 283530 337770 283558 338028
rect 283162 337742 283236 337770
rect 283208 336954 283236 337742
rect 283300 337742 283374 337770
rect 283484 337742 283558 337770
rect 283300 337074 283328 337742
rect 283378 337648 283434 337657
rect 283378 337583 283434 337592
rect 283288 337068 283340 337074
rect 283288 337010 283340 337016
rect 283012 336932 283064 336938
rect 283208 336926 283328 336954
rect 283012 336874 283064 336880
rect 282918 336560 282974 336569
rect 282918 336495 282974 336504
rect 283300 335918 283328 336926
rect 283288 335912 283340 335918
rect 283288 335854 283340 335860
rect 283196 335844 283248 335850
rect 283196 335786 283248 335792
rect 282828 335776 282880 335782
rect 282828 335718 282880 335724
rect 282840 329186 282868 335718
rect 283012 335096 283064 335102
rect 283012 335038 283064 335044
rect 283024 334257 283052 335038
rect 283208 334558 283236 335786
rect 283196 334552 283248 334558
rect 283196 334494 283248 334500
rect 283010 334248 283066 334257
rect 283010 334183 283066 334192
rect 282918 334112 282974 334121
rect 282918 334047 282974 334056
rect 282932 334014 282960 334047
rect 282920 334008 282972 334014
rect 282920 333950 282972 333956
rect 282828 329180 282880 329186
rect 282828 329122 282880 329128
rect 283392 327962 283420 337583
rect 283484 335850 283512 337742
rect 283622 337634 283650 338028
rect 283576 337606 283650 337634
rect 283472 335844 283524 335850
rect 283472 335786 283524 335792
rect 283472 335572 283524 335578
rect 283472 335514 283524 335520
rect 283484 328166 283512 335514
rect 283576 335442 283604 337606
rect 283714 337532 283742 338028
rect 283806 337634 283834 338028
rect 283898 337958 283926 338028
rect 283886 337952 283938 337958
rect 283886 337894 283938 337900
rect 283990 337895 284018 338028
rect 284082 337958 284110 338028
rect 284174 337963 284202 338028
rect 284070 337952 284122 337958
rect 283976 337886 284032 337895
rect 284070 337894 284122 337900
rect 284160 337954 284216 337963
rect 284160 337889 284216 337898
rect 284266 337890 284294 338028
rect 283976 337821 284032 337830
rect 284254 337884 284306 337890
rect 284254 337826 284306 337832
rect 284114 337784 284170 337793
rect 284358 337770 284386 338028
rect 284114 337719 284170 337728
rect 284312 337742 284386 337770
rect 283930 337648 283986 337657
rect 283806 337606 283880 337634
rect 283714 337504 283788 337532
rect 283656 337068 283708 337074
rect 283656 337010 283708 337016
rect 283564 335436 283616 335442
rect 283564 335378 283616 335384
rect 283564 332648 283616 332654
rect 283564 332590 283616 332596
rect 283472 328160 283524 328166
rect 283472 328102 283524 328108
rect 283380 327956 283432 327962
rect 283380 327898 283432 327904
rect 282656 316006 282776 316034
rect 282656 240786 282684 316006
rect 282644 240780 282696 240786
rect 282644 240722 282696 240728
rect 282920 236768 282972 236774
rect 282920 236710 282972 236716
rect 282932 16574 282960 236710
rect 282932 16546 283144 16574
rect 282276 3052 282328 3058
rect 282276 2994 282328 3000
rect 283116 480 283144 16546
rect 283576 3398 283604 332590
rect 283668 327894 283696 337010
rect 283760 335578 283788 337504
rect 283748 335572 283800 335578
rect 283748 335514 283800 335520
rect 283748 332648 283800 332654
rect 283748 332590 283800 332596
rect 283656 327888 283708 327894
rect 283656 327830 283708 327836
rect 283760 327758 283788 332590
rect 283852 328098 283880 337606
rect 283930 337583 283986 337592
rect 283944 332654 283972 337583
rect 284128 337550 284156 337719
rect 284116 337544 284168 337550
rect 284116 337486 284168 337492
rect 284312 335510 284340 337742
rect 284450 337634 284478 338028
rect 284542 337804 284570 338028
rect 284634 337929 284662 338028
rect 284620 337920 284676 337929
rect 284620 337855 284676 337864
rect 284542 337776 284616 337804
rect 284450 337606 284524 337634
rect 284390 335608 284446 335617
rect 284390 335543 284446 335552
rect 284300 335504 284352 335510
rect 284300 335446 284352 335452
rect 284024 335436 284076 335442
rect 284024 335378 284076 335384
rect 283932 332648 283984 332654
rect 283932 332590 283984 332596
rect 284036 331214 284064 335378
rect 284116 335368 284168 335374
rect 284404 335354 284432 335543
rect 284116 335310 284168 335316
rect 284312 335326 284432 335354
rect 284128 332654 284156 335310
rect 284116 332648 284168 332654
rect 284116 332590 284168 332596
rect 283944 331186 284064 331214
rect 283840 328092 283892 328098
rect 283840 328034 283892 328040
rect 283944 327826 283972 331186
rect 284312 329934 284340 335326
rect 284392 334008 284444 334014
rect 284392 333950 284444 333956
rect 284300 329928 284352 329934
rect 284300 329870 284352 329876
rect 283932 327820 283984 327826
rect 283932 327762 283984 327768
rect 283748 327752 283800 327758
rect 283748 327694 283800 327700
rect 284404 316034 284432 333950
rect 284496 329594 284524 337606
rect 284588 335442 284616 337776
rect 284726 337770 284754 338028
rect 284680 337742 284754 337770
rect 284576 335436 284628 335442
rect 284576 335378 284628 335384
rect 284680 335374 284708 337742
rect 284818 337634 284846 338028
rect 284772 337606 284846 337634
rect 284668 335368 284720 335374
rect 284668 335310 284720 335316
rect 284484 329588 284536 329594
rect 284484 329530 284536 329536
rect 284772 322522 284800 337606
rect 285048 337550 285076 373966
rect 285220 338020 285272 338026
rect 285220 337962 285272 337968
rect 285036 337544 285088 337550
rect 285036 337486 285088 337492
rect 284852 335368 284904 335374
rect 284852 335310 284904 335316
rect 284760 322516 284812 322522
rect 284760 322458 284812 322464
rect 284312 316006 284432 316034
rect 284312 3602 284340 316006
rect 284864 239698 284892 335310
rect 285036 335300 285088 335306
rect 285036 335242 285088 335248
rect 284944 329928 284996 329934
rect 284944 329870 284996 329876
rect 284852 239692 284904 239698
rect 284852 239634 284904 239640
rect 284392 238128 284444 238134
rect 284392 238070 284444 238076
rect 284300 3596 284352 3602
rect 284300 3538 284352 3544
rect 284404 3482 284432 238070
rect 284956 5234 284984 329870
rect 284944 5228 284996 5234
rect 284944 5170 284996 5176
rect 285048 4418 285076 335242
rect 285128 335232 285180 335238
rect 285128 335174 285180 335180
rect 285036 4412 285088 4418
rect 285036 4354 285088 4360
rect 285140 4214 285168 335174
rect 285232 237114 285260 337962
rect 285494 337920 285550 337929
rect 285494 337855 285550 337864
rect 285404 335504 285456 335510
rect 285404 335446 285456 335452
rect 285312 335436 285364 335442
rect 285312 335378 285364 335384
rect 285324 322454 285352 335378
rect 285312 322448 285364 322454
rect 285312 322390 285364 322396
rect 285416 322386 285444 335446
rect 285508 329934 285536 337855
rect 286322 335880 286378 335889
rect 286322 335815 286378 335824
rect 285586 334248 285642 334257
rect 285586 334183 285588 334192
rect 285640 334183 285642 334192
rect 285588 334154 285640 334160
rect 285680 331424 285732 331430
rect 285680 331366 285732 331372
rect 285496 329928 285548 329934
rect 285496 329870 285548 329876
rect 285404 322380 285456 322386
rect 285404 322322 285456 322328
rect 285220 237108 285272 237114
rect 285220 237050 285272 237056
rect 285692 16574 285720 331366
rect 285692 16546 286272 16574
rect 285128 4208 285180 4214
rect 285128 4150 285180 4156
rect 285404 3596 285456 3602
rect 285404 3538 285456 3544
rect 284312 3454 284432 3482
rect 283564 3392 283616 3398
rect 283564 3334 283616 3340
rect 284312 480 284340 3454
rect 285416 480 285444 3538
rect 286244 3482 286272 16546
rect 286336 5098 286364 335815
rect 286416 335164 286468 335170
rect 286416 335106 286468 335112
rect 286428 5506 286456 335106
rect 286520 219434 286548 390118
rect 288072 389768 288124 389774
rect 288072 389710 288124 389716
rect 287426 382256 287482 382265
rect 287426 382191 287482 382200
rect 287440 381750 287468 382191
rect 287428 381744 287480 381750
rect 287428 381686 287480 381692
rect 287426 377360 287482 377369
rect 287426 377295 287482 377304
rect 287440 376786 287468 377295
rect 287428 376780 287480 376786
rect 287428 376722 287480 376728
rect 287610 375864 287666 375873
rect 287610 375799 287666 375808
rect 287624 375426 287652 375799
rect 287612 375420 287664 375426
rect 287612 375362 287664 375368
rect 287794 372600 287850 372609
rect 287794 372535 287850 372544
rect 287808 371686 287836 372535
rect 287796 371680 287848 371686
rect 287796 371622 287848 371628
rect 287610 370968 287666 370977
rect 287610 370903 287666 370912
rect 287624 370598 287652 370903
rect 287612 370592 287664 370598
rect 287612 370534 287664 370540
rect 287978 367704 288034 367713
rect 287978 367639 288034 367648
rect 287992 367130 288020 367639
rect 287980 367124 288032 367130
rect 287980 367066 288032 367072
rect 287610 366072 287666 366081
rect 287610 366007 287666 366016
rect 287624 365770 287652 366007
rect 287612 365764 287664 365770
rect 287612 365706 287664 365712
rect 287610 362944 287666 362953
rect 287610 362879 287666 362888
rect 287624 362370 287652 362879
rect 287612 362364 287664 362370
rect 287612 362306 287664 362312
rect 287610 361312 287666 361321
rect 287610 361247 287666 361256
rect 287624 360670 287652 361247
rect 287612 360664 287664 360670
rect 287612 360606 287664 360612
rect 287610 359680 287666 359689
rect 287610 359615 287666 359624
rect 287624 359038 287652 359615
rect 287612 359032 287664 359038
rect 287612 358974 287664 358980
rect 287794 356416 287850 356425
rect 287794 356351 287850 356360
rect 287808 356114 287836 356351
rect 287796 356108 287848 356114
rect 287796 356050 287848 356056
rect 287518 353152 287574 353161
rect 287518 353087 287574 353096
rect 287532 351966 287560 353087
rect 287520 351960 287572 351966
rect 287520 351902 287572 351908
rect 287242 351520 287298 351529
rect 287242 351455 287244 351464
rect 287296 351455 287298 351464
rect 287244 351426 287296 351432
rect 287978 348392 288034 348401
rect 287978 348327 288034 348336
rect 287992 347818 288020 348327
rect 287980 347812 288032 347818
rect 287980 347754 288032 347760
rect 287978 346760 288034 346769
rect 287978 346695 288034 346704
rect 287992 346594 288020 346695
rect 287980 346588 288032 346594
rect 287980 346530 288032 346536
rect 287794 340232 287850 340241
rect 287794 340167 287850 340176
rect 287808 339522 287836 340167
rect 287796 339516 287848 339522
rect 287796 339458 287848 339464
rect 287426 338736 287482 338745
rect 287426 338671 287482 338680
rect 287440 338162 287468 338671
rect 287610 338192 287666 338201
rect 287428 338156 287480 338162
rect 287610 338127 287666 338136
rect 287428 338098 287480 338104
rect 287334 337512 287390 337521
rect 287334 337447 287390 337456
rect 286874 337376 286930 337385
rect 286874 337311 286930 337320
rect 286782 335472 286838 335481
rect 286782 335407 286838 335416
rect 286600 334552 286652 334558
rect 286600 334494 286652 334500
rect 286612 236910 286640 334494
rect 286692 332648 286744 332654
rect 286692 332590 286744 332596
rect 286704 236978 286732 332590
rect 286796 320890 286824 335407
rect 286888 331906 286916 337311
rect 286876 331900 286928 331906
rect 286876 331842 286928 331848
rect 287348 328454 287376 337447
rect 287624 337006 287652 338127
rect 287612 337000 287664 337006
rect 287612 336942 287664 336948
rect 287888 334484 287940 334490
rect 287888 334426 287940 334432
rect 287796 334144 287848 334150
rect 287796 334086 287848 334092
rect 287704 334076 287756 334082
rect 287704 334018 287756 334024
rect 287348 328426 287652 328454
rect 287624 322318 287652 328426
rect 287612 322312 287664 322318
rect 287612 322254 287664 322260
rect 286784 320884 286836 320890
rect 286784 320826 286836 320832
rect 287060 238060 287112 238066
rect 287060 238002 287112 238008
rect 286692 236972 286744 236978
rect 286692 236914 286744 236920
rect 286600 236904 286652 236910
rect 286600 236846 286652 236852
rect 286508 219428 286560 219434
rect 286508 219370 286560 219376
rect 287072 16574 287100 238002
rect 287072 16546 287376 16574
rect 286416 5500 286468 5506
rect 286416 5442 286468 5448
rect 286324 5092 286376 5098
rect 286324 5034 286376 5040
rect 286244 3454 286640 3482
rect 286612 480 286640 3454
rect 287348 490 287376 16546
rect 287716 3806 287744 334018
rect 287704 3800 287756 3806
rect 287704 3742 287756 3748
rect 287808 3670 287836 334086
rect 287900 3738 287928 334426
rect 287980 334212 288032 334218
rect 287980 334154 288032 334160
rect 287992 4010 288020 334154
rect 288084 239358 288112 389710
rect 288164 389360 288216 389366
rect 288164 389302 288216 389308
rect 288176 239426 288204 389302
rect 288346 387152 288402 387161
rect 288346 387087 288402 387096
rect 288360 387054 288388 387087
rect 288348 387048 288400 387054
rect 288348 386990 288400 386996
rect 288346 385520 288402 385529
rect 288346 385455 288402 385464
rect 288360 385082 288388 385455
rect 288348 385076 288400 385082
rect 288348 385018 288400 385024
rect 288346 383888 288402 383897
rect 288346 383823 288402 383832
rect 288360 383722 288388 383823
rect 288348 383716 288400 383722
rect 288348 383658 288400 383664
rect 288346 380624 288402 380633
rect 288346 380559 288402 380568
rect 288360 379574 288388 380559
rect 288348 379568 288400 379574
rect 288348 379510 288400 379516
rect 288346 378992 288402 379001
rect 288346 378927 288402 378936
rect 288360 378214 288388 378927
rect 288348 378208 288400 378214
rect 288348 378150 288400 378156
rect 288346 374232 288402 374241
rect 288346 374167 288348 374176
rect 288400 374167 288402 374176
rect 288348 374138 288400 374144
rect 288346 369336 288402 369345
rect 288346 369271 288402 369280
rect 288360 368558 288388 369271
rect 288348 368552 288400 368558
rect 288348 368494 288400 368500
rect 289096 365702 289124 390118
rect 291844 389904 291896 389910
rect 291844 389846 291896 389852
rect 290556 370592 290608 370598
rect 290556 370534 290608 370540
rect 289084 365696 289136 365702
rect 289084 365638 289136 365644
rect 288346 364440 288402 364449
rect 288346 364375 288348 364384
rect 288400 364375 288402 364384
rect 288348 364346 288400 364352
rect 289452 359032 289504 359038
rect 289452 358974 289504 358980
rect 288346 358048 288402 358057
rect 288346 357983 288402 357992
rect 288360 357474 288388 357983
rect 288348 357468 288400 357474
rect 288348 357410 288400 357416
rect 288346 354784 288402 354793
rect 288346 354719 288348 354728
rect 288400 354719 288402 354728
rect 288348 354690 288400 354696
rect 288346 350024 288402 350033
rect 288346 349959 288402 349968
rect 288360 349178 288388 349959
rect 288348 349172 288400 349178
rect 288348 349114 288400 349120
rect 288346 345128 288402 345137
rect 288346 345063 288348 345072
rect 288400 345063 288402 345072
rect 288348 345034 288400 345040
rect 288346 343496 288402 343505
rect 288346 343431 288402 343440
rect 288360 342310 288388 343431
rect 288348 342304 288400 342310
rect 288348 342246 288400 342252
rect 288346 341864 288402 341873
rect 288346 341799 288402 341808
rect 288360 340950 288388 341799
rect 288348 340944 288400 340950
rect 288348 340886 288400 340892
rect 288256 337952 288308 337958
rect 288256 337894 288308 337900
rect 288164 239420 288216 239426
rect 288164 239362 288216 239368
rect 288072 239352 288124 239358
rect 288072 239294 288124 239300
rect 288268 237046 288296 337894
rect 288440 335232 288492 335238
rect 288440 335174 288492 335180
rect 288348 329928 288400 329934
rect 288348 329870 288400 329876
rect 288360 237250 288388 329870
rect 288348 237244 288400 237250
rect 288348 237186 288400 237192
rect 288256 237040 288308 237046
rect 288256 236982 288308 236988
rect 288452 16574 288480 335174
rect 289360 335096 289412 335102
rect 289360 335038 289412 335044
rect 289268 334416 289320 334422
rect 289268 334358 289320 334364
rect 289084 334348 289136 334354
rect 289084 334290 289136 334296
rect 288452 16546 289032 16574
rect 287980 4004 288032 4010
rect 287980 3946 288032 3952
rect 287888 3732 287940 3738
rect 287888 3674 287940 3680
rect 287796 3664 287848 3670
rect 287796 3606 287848 3612
rect 287624 598 287836 626
rect 287624 490 287652 598
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 462 287652 490
rect 287808 480 287836 598
rect 289004 480 289032 16546
rect 289096 3534 289124 334290
rect 289176 334280 289228 334286
rect 289176 334222 289228 334228
rect 289188 3777 289216 334222
rect 289174 3768 289230 3777
rect 289174 3703 289230 3712
rect 289084 3528 289136 3534
rect 289084 3470 289136 3476
rect 289280 3466 289308 334358
rect 289372 3602 289400 335038
rect 289464 236638 289492 358974
rect 289544 338564 289596 338570
rect 289544 338506 289596 338512
rect 289452 236632 289504 236638
rect 289452 236574 289504 236580
rect 289556 236502 289584 338506
rect 290462 334384 290518 334393
rect 290462 334319 290518 334328
rect 289820 331492 289872 331498
rect 289820 331434 289872 331440
rect 289636 329588 289688 329594
rect 289636 329530 289688 329536
rect 289648 237182 289676 329530
rect 289636 237176 289688 237182
rect 289636 237118 289688 237124
rect 289544 236496 289596 236502
rect 289544 236438 289596 236444
rect 289360 3596 289412 3602
rect 289360 3538 289412 3544
rect 289268 3460 289320 3466
rect 289268 3402 289320 3408
rect 289832 490 289860 331434
rect 290476 3505 290504 334319
rect 290568 238474 290596 370534
rect 290648 334008 290700 334014
rect 290648 333950 290700 333956
rect 290556 238468 290608 238474
rect 290556 238410 290608 238416
rect 290660 3641 290688 333950
rect 291200 331424 291252 331430
rect 291200 331366 291252 331372
rect 291212 16574 291240 331366
rect 291856 238678 291884 389846
rect 291844 238672 291896 238678
rect 291844 238614 291896 238620
rect 291948 237930 291976 390458
rect 540428 390448 540480 390454
rect 540428 390390 540480 390396
rect 292212 390108 292264 390114
rect 292212 390050 292264 390056
rect 292028 390040 292080 390046
rect 292028 389982 292080 389988
rect 292040 238542 292068 389982
rect 292120 389700 292172 389706
rect 292120 389642 292172 389648
rect 292028 238536 292080 238542
rect 292028 238478 292080 238484
rect 292132 238270 292160 389642
rect 292224 239018 292252 390050
rect 395344 389972 395396 389978
rect 395344 389914 395396 389920
rect 296076 389836 296128 389842
rect 296076 389778 296128 389784
rect 294696 389632 294748 389638
rect 294696 389574 294748 389580
rect 293224 389224 293276 389230
rect 293224 389166 293276 389172
rect 292304 371680 292356 371686
rect 292304 371622 292356 371628
rect 292212 239012 292264 239018
rect 292212 238954 292264 238960
rect 292316 238406 292344 371622
rect 292396 339516 292448 339522
rect 292396 339458 292448 339464
rect 292304 238400 292356 238406
rect 292304 238342 292356 238348
rect 292120 238264 292172 238270
rect 292120 238206 292172 238212
rect 291936 237924 291988 237930
rect 291936 237866 291988 237872
rect 292408 237590 292436 339458
rect 292672 329996 292724 330002
rect 292672 329938 292724 329944
rect 292396 237584 292448 237590
rect 292396 237526 292448 237532
rect 292684 16574 292712 329938
rect 293236 238241 293264 389166
rect 293316 386436 293368 386442
rect 293316 386378 293368 386384
rect 293222 238232 293278 238241
rect 293222 238167 293278 238176
rect 293328 236745 293356 386378
rect 293408 376780 293460 376786
rect 293408 376722 293460 376728
rect 293420 238066 293448 376722
rect 293500 375420 293552 375426
rect 293500 375362 293552 375368
rect 293512 238202 293540 375362
rect 293592 374196 293644 374202
rect 293592 374138 293644 374144
rect 293604 238338 293632 374138
rect 294604 331356 294656 331362
rect 294604 331298 294656 331304
rect 293960 328840 294012 328846
rect 293960 328782 294012 328788
rect 293592 238332 293644 238338
rect 293592 238274 293644 238280
rect 293500 238196 293552 238202
rect 293500 238138 293552 238144
rect 293408 238060 293460 238066
rect 293408 238002 293460 238008
rect 293314 236736 293370 236745
rect 293314 236671 293370 236680
rect 293972 16574 294000 328782
rect 291212 16546 291424 16574
rect 292684 16546 293264 16574
rect 293972 16546 294552 16574
rect 290646 3632 290702 3641
rect 290646 3567 290702 3576
rect 290462 3496 290518 3505
rect 290462 3431 290518 3440
rect 290016 598 290228 626
rect 290016 490 290044 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 462 290044 490
rect 290200 480 290228 598
rect 291396 480 291424 16546
rect 292580 3324 292632 3330
rect 292580 3266 292632 3272
rect 292592 480 292620 3266
rect 293236 490 293264 16546
rect 294524 3210 294552 16546
rect 294616 3330 294644 331298
rect 294708 237658 294736 389574
rect 295984 389088 296036 389094
rect 295984 389030 296036 389036
rect 294788 381744 294840 381750
rect 294788 381686 294840 381692
rect 294800 238134 294828 381686
rect 294880 351484 294932 351490
rect 294880 351426 294932 351432
rect 294788 238128 294840 238134
rect 294788 238070 294840 238076
rect 294892 237794 294920 351426
rect 294972 346588 295024 346594
rect 294972 346530 295024 346536
rect 294880 237788 294932 237794
rect 294880 237730 294932 237736
rect 294696 237652 294748 237658
rect 294696 237594 294748 237600
rect 294984 236434 295012 346530
rect 295064 345092 295116 345098
rect 295064 345034 295116 345040
rect 295076 237522 295104 345034
rect 295064 237516 295116 237522
rect 295064 237458 295116 237464
rect 294972 236428 295024 236434
rect 294972 236370 295024 236376
rect 295996 46918 296024 389030
rect 296088 238610 296116 389778
rect 297364 389292 297416 389298
rect 297364 389234 297416 389240
rect 296168 365764 296220 365770
rect 296168 365706 296220 365712
rect 296076 238604 296128 238610
rect 296076 238546 296128 238552
rect 296180 236774 296208 365706
rect 296260 364404 296312 364410
rect 296260 364346 296312 364352
rect 296272 238746 296300 364346
rect 296352 362364 296404 362370
rect 296352 362306 296404 362312
rect 296260 238740 296312 238746
rect 296260 238682 296312 238688
rect 296364 237998 296392 362306
rect 296444 360664 296496 360670
rect 296444 360606 296496 360612
rect 296352 237992 296404 237998
rect 296352 237934 296404 237940
rect 296456 237862 296484 360606
rect 296536 338156 296588 338162
rect 296536 338098 296588 338104
rect 296444 237856 296496 237862
rect 296444 237798 296496 237804
rect 296548 237726 296576 338098
rect 297376 239154 297404 389234
rect 300124 389020 300176 389026
rect 300124 388962 300176 388968
rect 298744 385076 298796 385082
rect 298744 385018 298796 385024
rect 297456 378208 297508 378214
rect 297456 378150 297508 378156
rect 297468 239222 297496 378150
rect 297548 367124 297600 367130
rect 297548 367066 297600 367072
rect 297560 239290 297588 367066
rect 297732 340944 297784 340950
rect 297732 340886 297784 340892
rect 297640 338632 297692 338638
rect 297640 338574 297692 338580
rect 297548 239284 297600 239290
rect 297548 239226 297600 239232
rect 297456 239216 297508 239222
rect 297456 239158 297508 239164
rect 297364 239148 297416 239154
rect 297364 239090 297416 239096
rect 296536 237720 296588 237726
rect 296536 237662 296588 237668
rect 296168 236768 296220 236774
rect 296168 236710 296220 236716
rect 297652 236609 297680 338574
rect 297744 240038 297772 340886
rect 298100 331628 298152 331634
rect 298100 331570 298152 331576
rect 297732 240032 297784 240038
rect 297732 239974 297784 239980
rect 297638 236600 297694 236609
rect 297638 236535 297694 236544
rect 295984 46912 296036 46918
rect 295984 46854 296036 46860
rect 297272 4820 297324 4826
rect 297272 4762 297324 4768
rect 294604 3324 294656 3330
rect 294604 3266 294656 3272
rect 294524 3182 294920 3210
rect 293512 598 293724 626
rect 293512 490 293540 598
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 462 293540 490
rect 293696 480 293724 598
rect 294892 480 294920 3182
rect 296076 2916 296128 2922
rect 296076 2858 296128 2864
rect 296088 480 296116 2858
rect 297284 480 297312 4762
rect 298112 490 298140 331570
rect 298756 239086 298784 385018
rect 298928 356108 298980 356114
rect 298928 356050 298980 356056
rect 298836 354748 298888 354754
rect 298836 354690 298888 354696
rect 298744 239080 298796 239086
rect 298744 239022 298796 239028
rect 298848 236570 298876 354690
rect 298940 239494 298968 356050
rect 299020 347812 299072 347818
rect 299020 347754 299072 347760
rect 299032 239562 299060 347754
rect 299480 332716 299532 332722
rect 299480 332658 299532 332664
rect 299020 239556 299072 239562
rect 299020 239498 299072 239504
rect 298928 239488 298980 239494
rect 298928 239430 298980 239436
rect 298836 236564 298888 236570
rect 298836 236506 298888 236512
rect 299492 3482 299520 332658
rect 299572 331696 299624 331702
rect 299572 331638 299624 331644
rect 299584 4826 299612 331638
rect 300136 33114 300164 388962
rect 302884 388952 302936 388958
rect 302884 388894 302936 388900
rect 300216 335640 300268 335646
rect 300216 335582 300268 335588
rect 300124 33108 300176 33114
rect 300124 33050 300176 33056
rect 299572 4820 299624 4826
rect 299572 4762 299624 4768
rect 299492 3454 299704 3482
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3454
rect 300228 2922 300256 335582
rect 302240 332784 302292 332790
rect 302240 332726 302292 332732
rect 302252 16574 302280 332726
rect 302896 73166 302924 388894
rect 313924 388884 313976 388890
rect 313924 388826 313976 388832
rect 304262 336696 304318 336705
rect 304262 336631 304318 336640
rect 303620 330064 303672 330070
rect 303620 330006 303672 330012
rect 302884 73160 302936 73166
rect 302884 73102 302936 73108
rect 303632 16574 303660 330006
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 301964 4888 302016 4894
rect 301964 4830 302016 4836
rect 300768 4820 300820 4826
rect 300768 4762 300820 4768
rect 300216 2916 300268 2922
rect 300216 2858 300268 2864
rect 300780 480 300808 4762
rect 301976 480 302004 4830
rect 303172 480 303200 16546
rect 303908 490 303936 16546
rect 304276 4894 304304 336631
rect 304446 336560 304502 336569
rect 304446 336495 304502 336504
rect 304264 4888 304316 4894
rect 304264 4830 304316 4836
rect 304460 4826 304488 336495
rect 309140 332920 309192 332926
rect 309140 332862 309192 332868
rect 306380 332852 306432 332858
rect 306380 332794 306432 332800
rect 304448 4820 304500 4826
rect 304448 4762 304500 4768
rect 305552 2848 305604 2854
rect 305552 2790 305604 2796
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 2790
rect 306392 490 306420 332794
rect 309152 16574 309180 332862
rect 310520 330132 310572 330138
rect 310520 330074 310572 330080
rect 310532 16574 310560 330074
rect 313936 86970 313964 388826
rect 318064 388816 318116 388822
rect 318064 388758 318116 388764
rect 316684 335708 316736 335714
rect 316684 335650 316736 335656
rect 316040 335028 316092 335034
rect 316040 334970 316092 334976
rect 313924 86964 313976 86970
rect 313924 86906 313976 86912
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 307944 4344 307996 4350
rect 307944 4286 307996 4292
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 4286
rect 309048 4276 309100 4282
rect 309048 4218 309100 4224
rect 309060 480 309088 4218
rect 309796 490 309824 16546
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 16546
rect 314660 11008 314712 11014
rect 314660 10950 314712 10956
rect 313832 6724 313884 6730
rect 313832 6666 313884 6672
rect 312636 4480 312688 4486
rect 312636 4422 312688 4428
rect 312648 480 312676 4422
rect 313844 480 313872 6666
rect 314672 490 314700 10950
rect 316052 2854 316080 334970
rect 316132 330200 316184 330206
rect 316132 330142 316184 330148
rect 316144 16574 316172 330142
rect 316144 16546 316264 16574
rect 316040 2848 316092 2854
rect 316040 2790 316092 2796
rect 314856 598 315068 626
rect 314856 490 314884 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 462 314884 490
rect 315040 480 315068 598
rect 316236 480 316264 16546
rect 316696 2786 316724 335650
rect 317972 10940 318024 10946
rect 317972 10882 318024 10888
rect 317328 2848 317380 2854
rect 317328 2790 317380 2796
rect 316684 2780 316736 2786
rect 316684 2722 316736 2728
rect 317340 480 317368 2790
rect 317984 490 318012 10882
rect 318076 6866 318104 388758
rect 341524 336728 341576 336734
rect 341524 336670 341576 336676
rect 337384 335980 337436 335986
rect 337384 335922 337436 335928
rect 320180 333056 320232 333062
rect 320180 332998 320232 333004
rect 320192 16574 320220 332998
rect 322940 328908 322992 328914
rect 322940 328850 322992 328856
rect 320192 16546 320496 16574
rect 318064 6860 318116 6866
rect 318064 6802 318116 6808
rect 319720 4208 319772 4214
rect 319720 4150 319772 4156
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 317984 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 4150
rect 320468 490 320496 16546
rect 322112 10872 322164 10878
rect 322112 10814 322164 10820
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 10814
rect 322952 490 322980 328850
rect 329840 326460 329892 326466
rect 329840 326402 329892 326408
rect 329852 16574 329880 326402
rect 337396 16574 337424 335922
rect 329852 16546 330432 16574
rect 337396 16546 337608 16574
rect 324320 10804 324372 10810
rect 324320 10746 324372 10752
rect 324332 4214 324360 10746
rect 328736 10736 328788 10742
rect 328736 10678 328788 10684
rect 324412 6656 324464 6662
rect 324412 6598 324464 6604
rect 324320 4208 324372 4214
rect 324320 4150 324372 4156
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 6598
rect 328000 6588 328052 6594
rect 328000 6530 328052 6536
rect 326804 4480 326856 4486
rect 326804 4422 326856 4428
rect 325608 4208 325660 4214
rect 325608 4150 325660 4156
rect 325620 480 325648 4150
rect 326816 480 326844 4422
rect 328012 480 328040 6530
rect 328748 490 328776 10678
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 16546
rect 332692 10668 332744 10674
rect 332692 10610 332744 10616
rect 331588 6520 331640 6526
rect 331588 6462 331640 6468
rect 331600 480 331628 6462
rect 332704 480 332732 10610
rect 336280 10600 336332 10606
rect 336280 10542 336332 10548
rect 335084 6452 335136 6458
rect 335084 6394 335136 6400
rect 333888 4412 333940 4418
rect 333888 4354 333940 4360
rect 333900 480 333928 4354
rect 335096 480 335124 6394
rect 336292 480 336320 10542
rect 337580 2990 337608 16546
rect 339500 10532 339552 10538
rect 339500 10474 339552 10480
rect 338672 6384 338724 6390
rect 338672 6326 338724 6332
rect 337476 2984 337528 2990
rect 337476 2926 337528 2932
rect 337568 2984 337620 2990
rect 337568 2926 337620 2932
rect 337488 480 337516 2926
rect 338684 480 338712 6326
rect 339512 490 339540 10474
rect 341536 2990 341564 336670
rect 344284 336660 344336 336666
rect 344284 336602 344336 336608
rect 342904 10464 342956 10470
rect 342904 10406 342956 10412
rect 342168 6316 342220 6322
rect 342168 6258 342220 6264
rect 341524 2984 341576 2990
rect 341524 2926 341576 2932
rect 340972 2916 341024 2922
rect 340972 2858 341024 2864
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 2858
rect 342180 480 342208 6258
rect 342916 490 342944 10406
rect 344296 2922 344324 336602
rect 348424 336592 348476 336598
rect 348424 336534 348476 336540
rect 344560 335912 344612 335918
rect 344560 335854 344612 335860
rect 344468 335844 344520 335850
rect 344468 335786 344520 335792
rect 344376 335776 344428 335782
rect 344376 335718 344428 335724
rect 344388 236230 344416 335718
rect 344480 236298 344508 335786
rect 344572 236366 344600 335854
rect 344560 236360 344612 236366
rect 344560 236302 344612 236308
rect 344468 236292 344520 236298
rect 344468 236234 344520 236240
rect 344376 236224 344428 236230
rect 344376 236166 344428 236172
rect 346952 10396 347004 10402
rect 346952 10338 347004 10344
rect 345756 6248 345808 6254
rect 345756 6190 345808 6196
rect 344284 2916 344336 2922
rect 344284 2858 344336 2864
rect 344560 2848 344612 2854
rect 344560 2790 344612 2796
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 2790
rect 345768 480 345796 6190
rect 346964 480 346992 10338
rect 348436 2990 348464 336534
rect 355324 336524 355376 336530
rect 355324 336466 355376 336472
rect 351920 332988 351972 332994
rect 351920 332930 351972 332936
rect 351932 16574 351960 332930
rect 353300 330268 353352 330274
rect 353300 330210 353352 330216
rect 353312 16574 353340 330210
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 349160 10328 349212 10334
rect 349160 10270 349212 10276
rect 348056 2984 348108 2990
rect 348056 2926 348108 2932
rect 348424 2984 348476 2990
rect 348424 2926 348476 2932
rect 348068 480 348096 2926
rect 349172 1562 349200 10270
rect 349252 6180 349304 6186
rect 349252 6122 349304 6128
rect 349160 1556 349212 1562
rect 349160 1498 349212 1504
rect 349264 480 349292 6122
rect 351644 4616 351696 4622
rect 351644 4558 351696 4564
rect 350448 1556 350500 1562
rect 350448 1498 350500 1504
rect 350460 480 350488 1498
rect 351656 480 351684 4558
rect 352852 480 352880 16546
rect 353588 490 353616 16546
rect 355336 2922 355364 336466
rect 362224 336456 362276 336462
rect 362224 336398 362276 336404
rect 358820 333192 358872 333198
rect 358820 333134 358872 333140
rect 356060 333124 356112 333130
rect 356060 333066 356112 333072
rect 356072 16574 356100 333066
rect 357440 330336 357492 330342
rect 357440 330278 357492 330284
rect 356072 16546 356376 16574
rect 355232 2916 355284 2922
rect 355232 2858 355284 2864
rect 355324 2916 355376 2922
rect 355324 2858 355376 2864
rect 353864 598 354076 626
rect 353864 490 353892 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 462 353892 490
rect 354048 480 354076 598
rect 355244 480 355272 2858
rect 356348 480 356376 16546
rect 357452 6914 357480 330278
rect 357532 269816 357584 269822
rect 357532 269758 357584 269764
rect 357544 11762 357572 269758
rect 358832 16574 358860 333134
rect 360200 330404 360252 330410
rect 360200 330346 360252 330352
rect 360212 16574 360240 330346
rect 362236 16574 362264 336398
rect 369124 336388 369176 336394
rect 369124 336330 369176 336336
rect 362960 333940 363012 333946
rect 362960 333882 363012 333888
rect 362972 16574 363000 333882
rect 365720 333872 365772 333878
rect 365720 333814 365772 333820
rect 364340 330472 364392 330478
rect 364340 330414 364392 330420
rect 364352 16574 364380 330414
rect 358832 16546 359504 16574
rect 360212 16546 361160 16574
rect 362236 16546 362448 16574
rect 362972 16546 363552 16574
rect 364352 16546 364656 16574
rect 357532 11756 357584 11762
rect 357532 11698 357584 11704
rect 358728 11756 358780 11762
rect 358728 11698 358780 11704
rect 357452 6886 357572 6914
rect 357544 480 357572 6886
rect 358740 480 358768 11698
rect 359476 490 359504 16546
rect 359752 598 359964 626
rect 359752 490 359780 598
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 462 359780 490
rect 359936 480 359964 598
rect 361132 480 361160 16546
rect 362420 2854 362448 16546
rect 362316 2848 362368 2854
rect 362316 2790 362368 2796
rect 362408 2848 362460 2854
rect 362408 2790 362460 2796
rect 362328 480 362356 2790
rect 363524 480 363552 16546
rect 364628 480 364656 16546
rect 365732 2990 365760 333814
rect 367100 331764 367152 331770
rect 367100 331706 367152 331712
rect 367112 16574 367140 331706
rect 369136 16574 369164 336330
rect 376024 336320 376076 336326
rect 376024 336262 376076 336268
rect 369860 334960 369912 334966
rect 369860 334902 369912 334908
rect 369872 16574 369900 334902
rect 374000 334688 374052 334694
rect 374000 334630 374052 334636
rect 371240 331832 371292 331838
rect 371240 331774 371292 331780
rect 367112 16546 367784 16574
rect 369136 16546 369532 16574
rect 369872 16546 370176 16574
rect 365812 4616 365864 4622
rect 365812 4558 365864 4564
rect 365720 2984 365772 2990
rect 365720 2926 365772 2932
rect 365824 480 365852 4558
rect 367008 2984 367060 2990
rect 367008 2926 367060 2932
rect 367020 480 367048 2926
rect 367756 490 367784 16546
rect 369504 2990 369532 16546
rect 369400 2984 369452 2990
rect 369400 2926 369452 2932
rect 369492 2984 369544 2990
rect 369492 2926 369544 2932
rect 368032 598 368244 626
rect 368032 490 368060 598
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 462 368060 490
rect 368216 480 368244 598
rect 369412 480 369440 2926
rect 370148 490 370176 16546
rect 370424 598 370636 626
rect 370424 490 370452 598
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 462 370452 490
rect 370608 480 370636 598
rect 371252 490 371280 331774
rect 372620 18624 372672 18630
rect 372620 18566 372672 18572
rect 372632 16574 372660 18566
rect 372632 16546 372936 16574
rect 371528 598 371740 626
rect 371528 490 371556 598
rect 370566 -960 370678 480
rect 371252 462 371556 490
rect 371712 480 371740 598
rect 372908 480 372936 16546
rect 374012 6914 374040 334630
rect 374092 331220 374144 331226
rect 374092 331162 374144 331168
rect 374104 11762 374132 331162
rect 376036 16574 376064 336262
rect 382924 336252 382976 336258
rect 382924 336194 382976 336200
rect 376760 333804 376812 333810
rect 376760 333746 376812 333752
rect 376772 16574 376800 333746
rect 380900 333736 380952 333742
rect 380900 333678 380952 333684
rect 378140 331152 378192 331158
rect 378140 331094 378192 331100
rect 378152 16574 378180 331094
rect 380912 16574 380940 333678
rect 382372 331084 382424 331090
rect 382372 331026 382424 331032
rect 376036 16546 376616 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 380912 16546 381216 16574
rect 374092 11756 374144 11762
rect 374092 11698 374144 11704
rect 375288 11756 375340 11762
rect 375288 11698 375340 11704
rect 374012 6886 374132 6914
rect 374104 480 374132 6886
rect 375300 480 375328 11698
rect 376588 2922 376616 16546
rect 376484 2916 376536 2922
rect 376484 2858 376536 2864
rect 376576 2916 376628 2922
rect 376576 2858 376628 2864
rect 376496 480 376524 2858
rect 377692 480 377720 16546
rect 378428 490 378456 16546
rect 379980 4752 380032 4758
rect 379980 4694 380032 4700
rect 378704 598 378916 626
rect 378704 490 378732 598
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 462 378732 490
rect 378888 480 378916 598
rect 379992 480 380020 4694
rect 381188 480 381216 16546
rect 382384 480 382412 331026
rect 382936 2718 382964 336194
rect 391204 336184 391256 336190
rect 391204 336126 391256 336132
rect 387800 333668 387852 333674
rect 387800 333610 387852 333616
rect 383660 333600 383712 333606
rect 383660 333542 383712 333548
rect 383672 16574 383700 333542
rect 385040 331016 385092 331022
rect 385040 330958 385092 330964
rect 385052 16574 385080 330958
rect 386420 328364 386472 328370
rect 386420 328306 386472 328312
rect 386432 16574 386460 328306
rect 383672 16546 384344 16574
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 382924 2712 382976 2718
rect 382924 2654 382976 2660
rect 383568 2644 383620 2650
rect 383568 2586 383620 2592
rect 383580 480 383608 2586
rect 384316 490 384344 16546
rect 384592 598 384804 626
rect 384592 490 384620 598
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 462 384620 490
rect 384776 480 384804 598
rect 385972 480 386000 16546
rect 386708 490 386736 16546
rect 386984 598 387196 626
rect 386984 490 387012 598
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 462 387012 490
rect 387168 480 387196 598
rect 387812 490 387840 333610
rect 390652 333532 390704 333538
rect 390652 333474 390704 333480
rect 389180 330948 389232 330954
rect 389180 330890 389232 330896
rect 389192 16574 389220 330890
rect 390664 16574 390692 333474
rect 389192 16546 389496 16574
rect 390664 16546 391152 16574
rect 388088 598 388300 626
rect 388088 490 388116 598
rect 387126 -960 387238 480
rect 387812 462 388116 490
rect 388272 480 388300 598
rect 389468 480 389496 16546
rect 390652 2984 390704 2990
rect 390652 2926 390704 2932
rect 390664 480 390692 2926
rect 391124 2836 391152 16546
rect 391216 2990 391244 336126
rect 395356 334694 395384 389914
rect 418896 389564 418948 389570
rect 418896 389506 418948 389512
rect 398102 336424 398158 336433
rect 398102 336359 398158 336368
rect 395344 334688 395396 334694
rect 395344 334630 395396 334636
rect 394700 333464 394752 333470
rect 394700 333406 394752 333412
rect 391940 330880 391992 330886
rect 391940 330822 391992 330828
rect 391952 16574 391980 330822
rect 393320 328296 393372 328302
rect 393320 328238 393372 328244
rect 393332 16574 393360 328238
rect 394712 16574 394740 333406
rect 396080 330812 396132 330818
rect 396080 330754 396132 330760
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 391204 2984 391256 2990
rect 391204 2926 391256 2932
rect 391124 2808 391888 2836
rect 391860 480 391888 2808
rect 392596 490 392624 16546
rect 392872 598 393084 626
rect 392872 490 392900 598
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 462 392900 490
rect 393056 480 393084 598
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 396092 490 396120 330754
rect 398116 16574 398144 336359
rect 416042 336288 416098 336297
rect 416042 336223 416098 336232
rect 405004 336116 405056 336122
rect 405004 336058 405056 336064
rect 401600 334892 401652 334898
rect 401600 334834 401652 334840
rect 398840 333396 398892 333402
rect 398840 333338 398892 333344
rect 398116 16546 398328 16574
rect 397736 2916 397788 2922
rect 397736 2858 397788 2864
rect 396368 598 396580 626
rect 396368 490 396396 598
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 462 396396 490
rect 396552 480 396580 598
rect 397748 480 397776 2858
rect 398300 2854 398328 16546
rect 398852 6914 398880 333338
rect 398932 330744 398984 330750
rect 398932 330686 398984 330692
rect 398944 11762 398972 330686
rect 400220 328228 400272 328234
rect 400220 328170 400272 328176
rect 400232 16574 400260 328170
rect 401612 16574 401640 334834
rect 402980 330676 403032 330682
rect 402980 330618 403032 330624
rect 402992 16574 403020 330618
rect 400232 16546 400904 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 398932 11756 398984 11762
rect 398932 11698 398984 11704
rect 400128 11756 400180 11762
rect 400128 11698 400180 11704
rect 398852 6886 398972 6914
rect 398288 2848 398340 2854
rect 398288 2790 398340 2796
rect 398944 480 398972 6886
rect 400140 480 400168 11698
rect 400876 490 400904 16546
rect 401152 598 401364 626
rect 401152 490 401180 598
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 462 401180 490
rect 401336 480 401364 598
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 405016 2990 405044 336058
rect 407764 336048 407816 336054
rect 407764 335990 407816 335996
rect 405740 333328 405792 333334
rect 405740 333270 405792 333276
rect 405752 16574 405780 333270
rect 407212 330608 407264 330614
rect 407212 330550 407264 330556
rect 405752 16546 406056 16574
rect 404820 2984 404872 2990
rect 404820 2926 404872 2932
rect 405004 2984 405056 2990
rect 405004 2926 405056 2932
rect 405464 2984 405516 2990
rect 405516 2932 405688 2938
rect 405464 2926 405688 2932
rect 404832 480 404860 2926
rect 405476 2910 405688 2926
rect 405660 2854 405688 2910
rect 405648 2848 405700 2854
rect 405648 2790 405700 2796
rect 406028 480 406056 16546
rect 407224 480 407252 330550
rect 407776 2854 407804 335990
rect 415492 334824 415544 334830
rect 415492 334766 415544 334772
rect 412638 333976 412694 333985
rect 412638 333911 412694 333920
rect 408500 333260 408552 333266
rect 408500 333202 408552 333208
rect 408512 16574 408540 333202
rect 409880 330540 409932 330546
rect 409880 330482 409932 330488
rect 409892 16574 409920 330482
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 408408 2916 408460 2922
rect 408408 2858 408460 2864
rect 407764 2848 407816 2854
rect 407764 2790 407816 2796
rect 408420 480 408448 2858
rect 409156 490 409184 16546
rect 409432 598 409644 626
rect 409432 490 409460 598
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 462 409460 490
rect 409616 480 409644 598
rect 410812 480 410840 16546
rect 411904 5500 411956 5506
rect 411904 5442 411956 5448
rect 411916 480 411944 5442
rect 412652 490 412680 333911
rect 414020 328976 414072 328982
rect 414020 328918 414072 328924
rect 414032 16574 414060 328918
rect 415504 16574 415532 334766
rect 414032 16546 414336 16574
rect 415504 16546 415992 16574
rect 412928 598 413140 626
rect 412928 490 412956 598
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 462 412956 490
rect 413112 480 413140 598
rect 414308 480 414336 16546
rect 415492 2984 415544 2990
rect 415492 2926 415544 2932
rect 415504 480 415532 2926
rect 415964 2802 415992 16546
rect 416056 2990 416084 336223
rect 418802 333840 418858 333849
rect 418802 333775 418858 333784
rect 416780 329044 416832 329050
rect 416780 328986 416832 328992
rect 416792 16574 416820 328986
rect 416792 16546 417464 16574
rect 416044 2984 416096 2990
rect 416044 2926 416096 2932
rect 415964 2774 416728 2802
rect 416700 480 416728 2774
rect 417436 490 417464 16546
rect 418816 2990 418844 333775
rect 418908 234666 418936 389506
rect 439688 389496 439740 389502
rect 439688 389438 439740 389444
rect 540242 389464 540298 389473
rect 438308 389428 438360 389434
rect 438308 389370 438360 389376
rect 436744 337748 436796 337754
rect 436744 337690 436796 337696
rect 420920 337272 420972 337278
rect 420920 337214 420972 337220
rect 420182 336152 420238 336161
rect 420182 336087 420238 336096
rect 418896 234660 418948 234666
rect 418896 234602 418948 234608
rect 420196 16574 420224 336087
rect 420196 16546 420316 16574
rect 418804 2984 418856 2990
rect 418804 2926 418856 2932
rect 420184 2984 420236 2990
rect 420184 2926 420236 2932
rect 418988 2848 419040 2854
rect 418988 2790 419040 2796
rect 417712 598 417924 626
rect 417712 490 417740 598
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 462 417740 490
rect 417896 480 417924 598
rect 419000 480 419028 2790
rect 420196 480 420224 2926
rect 420288 2854 420316 16546
rect 420276 2848 420328 2854
rect 420276 2790 420328 2796
rect 420932 490 420960 337214
rect 422942 336016 422998 336025
rect 422942 335951 422998 335960
rect 422956 2922 422984 335951
rect 427082 334520 427138 334529
rect 427082 334455 427138 334464
rect 423678 333704 423734 333713
rect 423678 333639 423734 333648
rect 423692 16574 423720 333639
rect 423692 16546 423812 16574
rect 422576 2916 422628 2922
rect 422576 2858 422628 2864
rect 422944 2916 422996 2922
rect 422944 2858 422996 2864
rect 421208 598 421420 626
rect 421208 490 421236 598
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 462 421236 490
rect 421392 480 421420 598
rect 422588 480 422616 2858
rect 423784 480 423812 16546
rect 424968 5432 425020 5438
rect 424968 5374 425020 5380
rect 424980 480 425008 5374
rect 427096 3913 427124 334455
rect 432602 333568 432658 333577
rect 432602 333503 432658 333512
rect 429844 332580 429896 332586
rect 429844 332522 429896 332528
rect 427818 330848 427874 330857
rect 427818 330783 427874 330792
rect 427832 16574 427860 330783
rect 427832 16546 428504 16574
rect 427082 3904 427138 3913
rect 427082 3839 427138 3848
rect 427268 3052 427320 3058
rect 427268 2994 427320 3000
rect 426164 2984 426216 2990
rect 426164 2926 426216 2932
rect 426176 480 426204 2926
rect 427280 480 427308 2994
rect 428476 480 428504 16546
rect 429660 5364 429712 5370
rect 429660 5306 429712 5312
rect 429672 480 429700 5306
rect 429856 3058 429884 332522
rect 430580 332512 430632 332518
rect 430580 332454 430632 332460
rect 430592 16574 430620 332454
rect 430592 16546 430896 16574
rect 429844 3052 429896 3058
rect 429844 2994 429896 3000
rect 430868 480 430896 16546
rect 432052 5296 432104 5302
rect 432052 5238 432104 5244
rect 432064 480 432092 5238
rect 432616 2990 432644 333503
rect 434720 332444 434772 332450
rect 434720 332386 434772 332392
rect 434732 16574 434760 332386
rect 436650 272912 436706 272921
rect 436650 272847 436706 272856
rect 436664 272542 436692 272847
rect 436652 272536 436704 272542
rect 436652 272478 436704 272484
rect 436098 267472 436154 267481
rect 436098 267407 436154 267416
rect 436112 267034 436140 267407
rect 436100 267028 436152 267034
rect 436100 266970 436152 266976
rect 436112 266370 436140 266970
rect 436020 266342 436140 266370
rect 436020 239698 436048 266342
rect 436100 248396 436152 248402
rect 436100 248338 436152 248344
rect 436112 247353 436140 248338
rect 436098 247344 436154 247353
rect 436098 247279 436154 247288
rect 436756 245585 436784 337690
rect 438124 334756 438176 334762
rect 438124 334698 438176 334704
rect 436836 332308 436888 332314
rect 436836 332250 436888 332256
rect 436848 271946 436876 332250
rect 436928 326392 436980 326398
rect 436928 326334 436980 326340
rect 436940 287054 436968 326334
rect 436940 287026 437060 287054
rect 436848 271918 436968 271946
rect 436836 271856 436888 271862
rect 436836 271798 436888 271804
rect 436848 271289 436876 271798
rect 436834 271280 436890 271289
rect 436834 271215 436890 271224
rect 436836 270496 436888 270502
rect 436836 270438 436888 270444
rect 436848 270201 436876 270438
rect 436834 270192 436890 270201
rect 436834 270127 436890 270136
rect 436940 269074 436968 271918
rect 436928 269068 436980 269074
rect 436928 269010 436980 269016
rect 437032 267734 437060 287026
rect 437480 274644 437532 274650
rect 437480 274586 437532 274592
rect 437492 274281 437520 274586
rect 437478 274272 437534 274281
rect 437478 274207 437534 274216
rect 437386 272912 437442 272921
rect 437386 272847 437442 272856
rect 437296 269068 437348 269074
rect 437296 269010 437348 269016
rect 437308 268433 437336 269010
rect 437294 268424 437350 268433
rect 437294 268359 437350 268368
rect 437032 267706 437244 267734
rect 437216 265713 437244 267706
rect 437202 265704 437258 265713
rect 437202 265639 437258 265648
rect 436742 245576 436798 245585
rect 436742 245511 436798 245520
rect 436008 239692 436060 239698
rect 436008 239634 436060 239640
rect 437216 237969 437244 265639
rect 437308 238105 437336 268359
rect 437400 239630 437428 272847
rect 437388 239624 437440 239630
rect 437388 239566 437440 239572
rect 437294 238096 437350 238105
rect 437294 238031 437350 238040
rect 437202 237960 437258 237969
rect 437202 237895 437258 237904
rect 434732 16546 435128 16574
rect 434444 3052 434496 3058
rect 434444 2994 434496 3000
rect 432604 2984 432656 2990
rect 432604 2926 432656 2932
rect 433248 2848 433300 2854
rect 433248 2790 433300 2796
rect 433260 480 433288 2790
rect 434456 480 434484 2994
rect 435100 490 435128 16546
rect 437940 2984 437992 2990
rect 437940 2926 437992 2932
rect 436744 2916 436796 2922
rect 436744 2858 436796 2864
rect 435376 598 435588 626
rect 435376 490 435404 598
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 462 435404 490
rect 435560 480 435588 598
rect 436756 480 436784 2858
rect 437952 480 437980 2926
rect 438136 2854 438164 334698
rect 438214 333432 438270 333441
rect 438214 333367 438270 333376
rect 438228 2990 438256 333367
rect 438320 237454 438348 389370
rect 439502 333296 439558 333305
rect 439502 333231 439558 333240
rect 438858 330712 438914 330721
rect 438858 330647 438914 330656
rect 438766 274272 438822 274281
rect 438766 274207 438822 274216
rect 438674 271280 438730 271289
rect 438674 271215 438730 271224
rect 438582 270192 438638 270201
rect 438582 270127 438638 270136
rect 438596 239766 438624 270127
rect 438688 239902 438716 271215
rect 438676 239896 438728 239902
rect 438676 239838 438728 239844
rect 438780 239834 438808 274207
rect 438768 239828 438820 239834
rect 438768 239770 438820 239776
rect 438584 239760 438636 239766
rect 438584 239702 438636 239708
rect 438308 237448 438360 237454
rect 438308 237390 438360 237396
rect 438872 16574 438900 330647
rect 439136 240780 439188 240786
rect 439136 240722 439188 240728
rect 439148 236094 439176 240722
rect 439136 236088 439188 236094
rect 439136 236030 439188 236036
rect 438872 16546 439176 16574
rect 438216 2984 438268 2990
rect 438216 2926 438268 2932
rect 438124 2848 438176 2854
rect 438124 2790 438176 2796
rect 439148 480 439176 16546
rect 439516 2922 439544 333231
rect 439596 332376 439648 332382
rect 439596 332318 439648 332324
rect 439608 3058 439636 332318
rect 439700 237833 439728 389438
rect 540242 389399 540298 389408
rect 443644 388748 443696 388754
rect 443644 388690 443696 388696
rect 443656 325650 443684 388690
rect 447784 388136 447836 388142
rect 447784 388078 447836 388084
rect 446404 368552 446456 368558
rect 446404 368494 446456 368500
rect 446416 338774 446444 368494
rect 446404 338768 446456 338774
rect 446404 338710 446456 338716
rect 447048 328160 447100 328166
rect 447048 328102 447100 328108
rect 443644 325644 443696 325650
rect 443644 325586 443696 325592
rect 447060 322250 447088 328102
rect 447048 322244 447100 322250
rect 447048 322186 447100 322192
rect 447796 322114 447824 388078
rect 449164 388068 449216 388074
rect 449164 388010 449216 388016
rect 447784 322108 447836 322114
rect 447784 322050 447836 322056
rect 449176 322046 449204 388010
rect 481640 388000 481692 388006
rect 481640 387942 481692 387948
rect 471244 387048 471296 387054
rect 471244 386990 471296 386996
rect 468484 383716 468536 383722
rect 468484 383658 468536 383664
rect 465724 379568 465776 379574
rect 465724 379510 465776 379516
rect 464344 342304 464396 342310
rect 464344 342246 464396 342252
rect 464356 322658 464384 342246
rect 464344 322652 464396 322658
rect 464344 322594 464396 322600
rect 465736 322182 465764 379510
rect 467104 349172 467156 349178
rect 467104 349114 467156 349120
rect 467116 322930 467144 349114
rect 467840 338700 467892 338706
rect 467840 338642 467892 338648
rect 467104 322924 467156 322930
rect 467104 322866 467156 322872
rect 467852 322561 467880 338642
rect 468496 322590 468524 383658
rect 471256 322930 471284 386990
rect 474004 357468 474056 357474
rect 474004 357410 474056 357416
rect 472624 351960 472676 351966
rect 472624 351902 472676 351908
rect 471244 322924 471296 322930
rect 471244 322866 471296 322872
rect 472256 322856 472308 322862
rect 472256 322798 472308 322804
rect 469404 322652 469456 322658
rect 469404 322594 469456 322600
rect 468484 322584 468536 322590
rect 467838 322552 467894 322561
rect 469416 322561 469444 322594
rect 468484 322526 468536 322532
rect 469402 322552 469458 322561
rect 467838 322487 467894 322496
rect 469402 322487 469458 322496
rect 465724 322176 465776 322182
rect 465724 322118 465776 322124
rect 470692 322108 470744 322114
rect 470692 322050 470744 322056
rect 449164 322040 449216 322046
rect 449164 321982 449216 321988
rect 470704 321609 470732 322050
rect 471980 322040 472032 322046
rect 471980 321982 472032 321988
rect 471992 321609 472020 321982
rect 472268 321609 472296 322798
rect 472636 322658 472664 351902
rect 474016 322862 474044 357410
rect 479524 337680 479576 337686
rect 479524 337622 479576 337628
rect 476028 328092 476080 328098
rect 476028 328034 476080 328040
rect 474004 322856 474056 322862
rect 474004 322798 474056 322804
rect 472624 322652 472676 322658
rect 472624 322594 472676 322600
rect 474556 322652 474608 322658
rect 474556 322594 474608 322600
rect 474568 322561 474596 322594
rect 474554 322552 474610 322561
rect 474554 322487 474610 322496
rect 476040 322114 476068 328034
rect 476580 328024 476632 328030
rect 476580 327966 476632 327972
rect 476592 322561 476620 327966
rect 479536 322930 479564 337622
rect 479524 322924 479576 322930
rect 479524 322866 479576 322872
rect 480628 322924 480680 322930
rect 480628 322866 480680 322872
rect 479156 322856 479208 322862
rect 479156 322798 479208 322804
rect 479168 322561 479196 322798
rect 476578 322552 476634 322561
rect 476578 322487 476634 322496
rect 479154 322552 479210 322561
rect 479154 322487 479210 322496
rect 476028 322108 476080 322114
rect 476028 322050 476080 322056
rect 475476 321836 475528 321842
rect 475476 321778 475528 321784
rect 475488 321609 475516 321778
rect 478236 321768 478288 321774
rect 478236 321710 478288 321716
rect 478248 321609 478276 321710
rect 480640 321609 480668 322866
rect 481652 322561 481680 387942
rect 485780 387932 485832 387938
rect 485780 387874 485832 387880
rect 483020 337612 483072 337618
rect 483020 337554 483072 337560
rect 481732 327956 481784 327962
rect 481732 327898 481784 327904
rect 481638 322552 481694 322561
rect 481638 322487 481694 322496
rect 481744 321638 481772 327898
rect 483032 322561 483060 337554
rect 484860 327888 484912 327894
rect 484860 327830 484912 327836
rect 484872 322561 484900 327830
rect 483018 322552 483074 322561
rect 483018 322487 483074 322496
rect 484858 322552 484914 322561
rect 484858 322487 484914 322496
rect 484400 322312 484452 322318
rect 484400 322254 484452 322260
rect 481732 321632 481784 321638
rect 470690 321600 470746 321609
rect 470690 321535 470746 321544
rect 471978 321600 472034 321609
rect 471978 321535 472034 321544
rect 472254 321600 472310 321609
rect 472254 321535 472310 321544
rect 475474 321600 475530 321609
rect 475474 321535 475530 321544
rect 478234 321600 478290 321609
rect 478234 321535 478290 321544
rect 480626 321600 480682 321609
rect 484412 321609 484440 322254
rect 485792 322017 485820 387874
rect 537484 387864 537536 387870
rect 537484 387806 537536 387812
rect 488540 338768 488592 338774
rect 488540 338710 488592 338716
rect 488552 322561 488580 338710
rect 530676 337476 530728 337482
rect 530676 337418 530728 337424
rect 519542 330440 519598 330449
rect 519542 330375 519598 330384
rect 490564 327820 490616 327826
rect 490564 327762 490616 327768
rect 490576 322561 490604 327762
rect 492680 327752 492732 327758
rect 492680 327694 492732 327700
rect 492692 322561 492720 327694
rect 496820 322788 496872 322794
rect 496820 322730 496872 322736
rect 494244 322720 494296 322726
rect 494244 322662 494296 322668
rect 488538 322552 488594 322561
rect 488538 322487 488594 322496
rect 490562 322552 490618 322561
rect 490562 322487 490618 322496
rect 492678 322552 492734 322561
rect 492678 322487 492734 322496
rect 492220 322108 492272 322114
rect 492220 322050 492272 322056
rect 485778 322008 485834 322017
rect 485778 321943 485834 321952
rect 488172 321632 488224 321638
rect 481732 321574 481784 321580
rect 484398 321600 484454 321609
rect 480626 321535 480682 321544
rect 484398 321535 484454 321544
rect 488170 321600 488172 321609
rect 492232 321609 492260 322050
rect 494256 321609 494284 322662
rect 495532 322244 495584 322250
rect 495532 322186 495584 322192
rect 495544 321609 495572 322186
rect 496832 321609 496860 322730
rect 506940 322652 506992 322658
rect 506940 322594 506992 322600
rect 504180 322584 504232 322590
rect 504180 322526 504232 322532
rect 498660 322448 498712 322454
rect 498660 322390 498712 322396
rect 498200 322380 498252 322386
rect 498200 322322 498252 322328
rect 498212 321609 498240 322322
rect 498672 321609 498700 322390
rect 501052 322176 501104 322182
rect 501052 322118 501104 322124
rect 500684 321904 500736 321910
rect 500684 321846 500736 321852
rect 500696 321609 500724 321846
rect 501064 321609 501092 322118
rect 503260 321972 503312 321978
rect 503260 321914 503312 321920
rect 503272 321609 503300 321914
rect 504192 321609 504220 322526
rect 505468 322516 505520 322522
rect 505468 322458 505520 322464
rect 505480 321609 505508 322458
rect 506952 321609 506980 322594
rect 519556 322425 519584 330375
rect 519542 322416 519598 322425
rect 519542 322351 519598 322360
rect 519556 322250 519584 322351
rect 519544 322244 519596 322250
rect 519544 322186 519596 322192
rect 530688 321638 530716 337418
rect 536840 337204 536892 337210
rect 536840 337146 536892 337152
rect 530032 321632 530084 321638
rect 488224 321600 488226 321609
rect 488170 321535 488226 321544
rect 492218 321600 492274 321609
rect 492218 321535 492274 321544
rect 494242 321600 494298 321609
rect 494242 321535 494298 321544
rect 495530 321600 495586 321609
rect 495530 321535 495586 321544
rect 496818 321600 496874 321609
rect 496818 321535 496874 321544
rect 498198 321600 498254 321609
rect 498198 321535 498254 321544
rect 498658 321600 498714 321609
rect 498658 321535 498714 321544
rect 500682 321600 500738 321609
rect 500682 321535 500738 321544
rect 501050 321600 501106 321609
rect 501050 321535 501106 321544
rect 503258 321600 503314 321609
rect 503258 321535 503314 321544
rect 504178 321600 504234 321609
rect 504178 321535 504234 321544
rect 505466 321600 505522 321609
rect 505466 321535 505522 321544
rect 506938 321600 506994 321609
rect 506938 321535 506994 321544
rect 530030 321600 530032 321609
rect 530676 321632 530728 321638
rect 530084 321600 530086 321609
rect 530676 321574 530728 321580
rect 530030 321535 530086 321544
rect 439872 240032 439924 240038
rect 439872 239974 439924 239980
rect 439884 239850 439912 239974
rect 445668 239964 445720 239970
rect 445668 239906 445720 239912
rect 445574 239864 445630 239873
rect 439884 239822 440280 239850
rect 439686 237824 439742 237833
rect 439686 237759 439742 237768
rect 440252 236162 440280 239822
rect 445574 239799 445630 239808
rect 445588 239193 445616 239799
rect 445680 239329 445708 239906
rect 445760 239896 445812 239902
rect 522672 239896 522724 239902
rect 445760 239838 445812 239844
rect 445850 239864 445906 239873
rect 445772 239698 445800 239838
rect 445850 239799 445906 239808
rect 451094 239864 451150 239873
rect 451094 239799 451150 239808
rect 452750 239864 452806 239873
rect 452750 239799 452806 239808
rect 460938 239864 460994 239873
rect 460938 239799 460994 239808
rect 522670 239864 522672 239873
rect 522724 239864 522726 239873
rect 522670 239799 522726 239808
rect 523130 239864 523186 239873
rect 523130 239799 523132 239808
rect 445864 239698 445892 239799
rect 451108 239698 451136 239799
rect 445760 239692 445812 239698
rect 445760 239634 445812 239640
rect 445852 239692 445904 239698
rect 445852 239634 445904 239640
rect 451096 239692 451148 239698
rect 451096 239634 451148 239640
rect 451188 239692 451240 239698
rect 451188 239634 451240 239640
rect 451200 239578 451228 239634
rect 451108 239550 451228 239578
rect 452764 239562 452792 239799
rect 456064 239692 456116 239698
rect 456064 239634 456116 239640
rect 456076 239562 456104 239634
rect 460952 239562 460980 239799
rect 523184 239799 523186 239808
rect 523132 239770 523184 239776
rect 523040 239760 523092 239766
rect 462410 239728 462466 239737
rect 462410 239663 462466 239672
rect 473174 239728 473230 239737
rect 473174 239663 473230 239672
rect 475658 239728 475714 239737
rect 523130 239728 523186 239737
rect 523092 239708 523130 239714
rect 523040 239702 523130 239708
rect 523052 239686 523130 239702
rect 475658 239663 475714 239672
rect 523130 239663 523186 239672
rect 452752 239556 452804 239562
rect 451108 239329 451136 239550
rect 452752 239498 452804 239504
rect 456064 239556 456116 239562
rect 456064 239498 456116 239504
rect 460940 239556 460992 239562
rect 460940 239498 460992 239504
rect 461032 239556 461084 239562
rect 461032 239498 461084 239504
rect 452568 239488 452620 239494
rect 452568 239430 452620 239436
rect 452580 239329 452608 239430
rect 461044 239329 461072 239498
rect 445666 239320 445722 239329
rect 445666 239255 445722 239264
rect 451094 239320 451150 239329
rect 451094 239255 451150 239264
rect 452566 239320 452622 239329
rect 452566 239255 452622 239264
rect 461030 239320 461086 239329
rect 461030 239255 461086 239264
rect 445574 239184 445630 239193
rect 445574 239119 445630 239128
rect 452658 239184 452714 239193
rect 452658 239119 452714 239128
rect 440240 236156 440292 236162
rect 440240 236098 440292 236104
rect 441620 234728 441672 234734
rect 441620 234670 441672 234676
rect 440332 232960 440384 232966
rect 440332 232902 440384 232908
rect 439596 3052 439648 3058
rect 439596 2994 439648 3000
rect 439504 2916 439556 2922
rect 439504 2858 439556 2864
rect 440344 480 440372 232902
rect 441632 16574 441660 234670
rect 448612 233776 448664 233782
rect 448612 233718 448664 233724
rect 445760 233708 445812 233714
rect 445760 233650 445812 233656
rect 443000 232892 443052 232898
rect 443000 232834 443052 232840
rect 443012 16574 443040 232834
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 441528 3052 441580 3058
rect 441528 2994 441580 3000
rect 441540 480 441568 2994
rect 442644 480 442672 16546
rect 443380 490 443408 16546
rect 445024 3120 445076 3126
rect 445024 3062 445076 3068
rect 443656 598 443868 626
rect 443656 490 443684 598
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 462 443684 490
rect 443840 480 443868 598
rect 445036 480 445064 3062
rect 445772 490 445800 233650
rect 447140 177404 447192 177410
rect 447140 177346 447192 177352
rect 447152 16574 447180 177346
rect 447152 16546 447456 16574
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 16546
rect 448624 11762 448652 233718
rect 452672 16574 452700 239119
rect 462320 237584 462372 237590
rect 462320 237526 462372 237532
rect 462332 237289 462360 237526
rect 462318 237280 462374 237289
rect 462318 237215 462374 237224
rect 461122 236872 461178 236881
rect 461122 236807 461178 236816
rect 461136 236502 461164 236807
rect 461124 236496 461176 236502
rect 461124 236438 461176 236444
rect 459560 234864 459612 234870
rect 459560 234806 459612 234812
rect 456892 234796 456944 234802
rect 456892 234738 456944 234744
rect 452672 16546 453344 16574
rect 448612 11756 448664 11762
rect 448612 11698 448664 11704
rect 449808 11756 449860 11762
rect 449808 11698 449860 11704
rect 448612 2916 448664 2922
rect 448612 2858 448664 2864
rect 448624 480 448652 2858
rect 449820 480 449848 11698
rect 450912 5160 450964 5166
rect 450912 5102 450964 5108
rect 450924 480 450952 5102
rect 452108 2848 452160 2854
rect 452108 2790 452160 2796
rect 452120 480 452148 2790
rect 453316 480 453344 16546
rect 454500 5228 454552 5234
rect 454500 5170 454552 5176
rect 454512 480 454540 5170
rect 455696 5024 455748 5030
rect 455696 4966 455748 4972
rect 455708 480 455736 4966
rect 456904 480 456932 234738
rect 459572 16574 459600 234806
rect 462424 219434 462452 239663
rect 465262 239592 465318 239601
rect 465262 239527 465318 239536
rect 471978 239592 472034 239601
rect 473188 239562 473216 239663
rect 471978 239527 472034 239536
rect 473176 239556 473228 239562
rect 465080 237652 465132 237658
rect 465080 237594 465132 237600
rect 463700 237516 463752 237522
rect 463700 237458 463752 237464
rect 463712 237289 463740 237458
rect 465092 237289 465120 237594
rect 463698 237280 463754 237289
rect 463698 237215 463754 237224
rect 465078 237280 465134 237289
rect 465078 237215 465134 237224
rect 465078 236872 465134 236881
rect 465078 236807 465134 236816
rect 465092 236434 465120 236807
rect 465080 236428 465132 236434
rect 465080 236370 465132 236376
rect 463700 233844 463752 233850
rect 463700 233786 463752 233792
rect 462332 219406 462452 219434
rect 459572 16546 459968 16574
rect 458088 3188 458140 3194
rect 458088 3130 458140 3136
rect 458100 480 458128 3130
rect 459192 3052 459244 3058
rect 459192 2994 459244 3000
rect 459204 480 459232 2994
rect 459940 490 459968 16546
rect 461584 3256 461636 3262
rect 461584 3198 461636 3204
rect 460216 598 460428 626
rect 460216 490 460244 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 462 460244 490
rect 460400 480 460428 598
rect 461596 480 461624 3198
rect 462332 490 462360 219406
rect 463712 16574 463740 233786
rect 465172 232824 465224 232830
rect 465172 232766 465224 232772
rect 463712 16546 464016 16574
rect 462608 598 462820 626
rect 462608 490 462636 598
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462332 462 462636 490
rect 462792 480 462820 598
rect 463988 480 464016 16546
rect 465184 480 465212 232766
rect 465276 16574 465304 239527
rect 468482 239456 468538 239465
rect 471992 239426 472020 239527
rect 473176 239498 473228 239504
rect 468482 239391 468538 239400
rect 471980 239420 472032 239426
rect 467196 237788 467248 237794
rect 467196 237730 467248 237736
rect 467208 237697 467236 237730
rect 467840 237720 467892 237726
rect 467194 237688 467250 237697
rect 467194 237623 467250 237632
rect 467838 237688 467840 237697
rect 467892 237688 467894 237697
rect 467838 237623 467894 237632
rect 467840 237312 467892 237318
rect 467838 237280 467840 237289
rect 467892 237280 467894 237289
rect 467838 237215 467894 237224
rect 466460 234592 466512 234598
rect 466460 234534 466512 234540
rect 466472 16574 466500 234534
rect 465276 16546 465856 16574
rect 466472 16546 467512 16574
rect 465828 490 465856 16546
rect 466104 598 466316 626
rect 466104 490 466132 598
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 462 466132 490
rect 466288 480 466316 598
rect 467484 480 467512 16546
rect 468496 3398 468524 239391
rect 471980 239362 472032 239368
rect 475672 239358 475700 239663
rect 505008 239624 505060 239630
rect 479338 239592 479394 239601
rect 479338 239527 479394 239536
rect 487894 239592 487950 239601
rect 487894 239527 487950 239536
rect 495622 239592 495678 239601
rect 495622 239527 495678 239536
rect 496818 239592 496874 239601
rect 496818 239527 496874 239536
rect 500498 239592 500554 239601
rect 500498 239527 500554 239536
rect 501878 239592 501934 239601
rect 501878 239527 501934 239536
rect 503074 239592 503130 239601
rect 505008 239566 505060 239572
rect 505558 239592 505614 239601
rect 503074 239527 503130 239536
rect 479352 239494 479380 239527
rect 479340 239488 479392 239494
rect 479340 239430 479392 239436
rect 475660 239352 475712 239358
rect 475660 239294 475712 239300
rect 487908 239290 487936 239527
rect 487896 239284 487948 239290
rect 487896 239226 487948 239232
rect 495636 238950 495664 239527
rect 495624 238944 495676 238950
rect 495624 238886 495676 238892
rect 496832 238882 496860 239527
rect 496820 238876 496872 238882
rect 496820 238818 496872 238824
rect 500512 238814 500540 239527
rect 501892 239222 501920 239527
rect 501880 239216 501932 239222
rect 501880 239158 501932 239164
rect 503088 239154 503116 239527
rect 503076 239148 503128 239154
rect 503076 239090 503128 239096
rect 500500 238808 500552 238814
rect 500500 238750 500552 238756
rect 485412 238740 485464 238746
rect 485412 238682 485464 238688
rect 477684 238672 477736 238678
rect 477682 238640 477684 238649
rect 485424 238649 485452 238682
rect 477736 238640 477738 238649
rect 477682 238575 477738 238584
rect 483386 238640 483442 238649
rect 483386 238575 483442 238584
rect 484398 238640 484454 238649
rect 484398 238575 484400 238584
rect 483400 238542 483428 238575
rect 484452 238575 484454 238584
rect 485410 238640 485466 238649
rect 485410 238575 485466 238584
rect 484400 238546 484452 238552
rect 483388 238536 483440 238542
rect 482282 238504 482338 238513
rect 483388 238478 483440 238484
rect 484858 238504 484914 238513
rect 482282 238439 482284 238448
rect 482336 238439 482338 238448
rect 484858 238439 484914 238448
rect 482284 238410 482336 238416
rect 484872 238406 484900 238439
rect 484860 238400 484912 238406
rect 476578 238368 476634 238377
rect 476578 238303 476634 238312
rect 480626 238368 480682 238377
rect 480626 238303 480682 238312
rect 481730 238368 481786 238377
rect 484860 238342 484912 238348
rect 485962 238368 486018 238377
rect 481730 238303 481786 238312
rect 485962 238303 486018 238312
rect 488170 238368 488226 238377
rect 488170 238303 488172 238312
rect 476592 237930 476620 238303
rect 476580 237924 476632 237930
rect 476580 237866 476632 237872
rect 480640 237862 480668 238303
rect 481744 237998 481772 238303
rect 485976 238270 486004 238303
rect 488224 238303 488226 238312
rect 488172 238274 488224 238280
rect 485964 238264 486016 238270
rect 485964 238206 486016 238212
rect 491666 238232 491722 238241
rect 491666 238167 491668 238176
rect 491720 238167 491722 238176
rect 492770 238232 492826 238241
rect 492770 238167 492826 238176
rect 495162 238232 495218 238241
rect 495162 238167 495218 238176
rect 491668 238138 491720 238144
rect 492784 238066 492812 238167
rect 495176 238134 495204 238167
rect 495164 238128 495216 238134
rect 495164 238070 495216 238076
rect 492772 238060 492824 238066
rect 492772 238002 492824 238008
rect 481732 237992 481784 237998
rect 481732 237934 481784 237940
rect 480628 237856 480680 237862
rect 480628 237798 480680 237804
rect 485780 237448 485832 237454
rect 485780 237390 485832 237396
rect 470600 237380 470652 237386
rect 470600 237322 470652 237328
rect 470612 237289 470640 237322
rect 485792 237289 485820 237390
rect 505020 237386 505048 239566
rect 505558 239527 505614 239536
rect 506754 239592 506810 239601
rect 506754 239527 506810 239536
rect 505572 239086 505600 239527
rect 505560 239080 505612 239086
rect 505560 239022 505612 239028
rect 506768 239018 506796 239527
rect 506756 239012 506808 239018
rect 506756 238954 506808 238960
rect 505008 237380 505060 237386
rect 505008 237322 505060 237328
rect 521660 237380 521712 237386
rect 521660 237322 521712 237328
rect 521672 237289 521700 237322
rect 469218 237280 469274 237289
rect 469218 237215 469274 237224
rect 470598 237280 470654 237289
rect 470598 237215 470654 237224
rect 485778 237280 485834 237289
rect 485778 237215 485834 237224
rect 498198 237280 498254 237289
rect 498198 237215 498254 237224
rect 503718 237280 503774 237289
rect 503718 237215 503720 237224
rect 469232 236706 469260 237215
rect 498212 237182 498240 237215
rect 503772 237215 503774 237224
rect 521658 237280 521714 237289
rect 521658 237215 521714 237224
rect 503720 237186 503772 237192
rect 498200 237176 498252 237182
rect 490286 237144 490342 237153
rect 490286 237079 490342 237088
rect 492678 237144 492734 237153
rect 492678 237079 492680 237088
rect 490300 236910 490328 237079
rect 492732 237079 492734 237088
rect 494058 237144 494114 237153
rect 498200 237118 498252 237124
rect 494058 237079 494114 237088
rect 492680 237050 492732 237056
rect 494072 237046 494100 237079
rect 494060 237040 494112 237046
rect 491298 237008 491354 237017
rect 494060 236982 494112 236988
rect 491298 236943 491300 236952
rect 491352 236943 491354 236952
rect 491300 236914 491352 236920
rect 490288 236904 490340 236910
rect 471978 236872 472034 236881
rect 471978 236807 472034 236816
rect 473358 236872 473414 236881
rect 473358 236807 473360 236816
rect 469220 236700 469272 236706
rect 469220 236642 469272 236648
rect 471992 236638 472020 236807
rect 473412 236807 473414 236816
rect 474738 236872 474794 236881
rect 474738 236807 474794 236816
rect 476118 236872 476174 236881
rect 476118 236807 476174 236816
rect 485778 236872 485834 236881
rect 485778 236807 485834 236816
rect 488538 236872 488594 236881
rect 490288 236846 490340 236852
rect 488538 236807 488594 236816
rect 473360 236778 473412 236784
rect 471980 236632 472032 236638
rect 471980 236574 472032 236580
rect 470874 236328 470930 236337
rect 474752 236298 474780 236807
rect 476132 236570 476160 236807
rect 485792 236774 485820 236807
rect 485780 236768 485832 236774
rect 485780 236710 485832 236716
rect 476120 236564 476172 236570
rect 476120 236506 476172 236512
rect 488552 236366 488580 236807
rect 488540 236360 488592 236366
rect 488540 236302 488592 236308
rect 470874 236263 470930 236272
rect 474740 236292 474792 236298
rect 470888 236230 470916 236263
rect 474740 236234 474792 236240
rect 470876 236224 470928 236230
rect 469218 236192 469274 236201
rect 470876 236166 470928 236172
rect 477498 236192 477554 236201
rect 469218 236127 469274 236136
rect 477498 236127 477554 236136
rect 495438 236192 495494 236201
rect 495438 236127 495440 236136
rect 469232 236094 469260 236127
rect 469220 236088 469272 236094
rect 469220 236030 469272 236036
rect 475384 235000 475436 235006
rect 475384 234942 475436 234948
rect 472624 234932 472676 234938
rect 472624 234874 472676 234880
rect 470600 234524 470652 234530
rect 470600 234466 470652 234472
rect 468668 5092 468720 5098
rect 468668 5034 468720 5040
rect 468484 3392 468536 3398
rect 468484 3334 468536 3340
rect 468680 480 468708 5034
rect 469864 3392 469916 3398
rect 469864 3334 469916 3340
rect 469876 480 469904 3334
rect 470612 490 470640 234466
rect 472636 3398 472664 234874
rect 472716 234456 472768 234462
rect 472716 234398 472768 234404
rect 472624 3392 472676 3398
rect 472624 3334 472676 3340
rect 472256 3256 472308 3262
rect 472256 3198 472308 3204
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 3198
rect 472728 3126 472756 234398
rect 473452 3392 473504 3398
rect 473452 3334 473504 3340
rect 472716 3120 472768 3126
rect 472716 3062 472768 3068
rect 473464 480 473492 3334
rect 475396 3330 475424 234942
rect 477512 234666 477540 236127
rect 495492 236127 495494 236136
rect 495440 236098 495492 236104
rect 488540 235952 488592 235958
rect 488540 235894 488592 235900
rect 484400 235204 484452 235210
rect 484400 235146 484452 235152
rect 483664 235136 483716 235142
rect 483664 235078 483716 235084
rect 481732 235068 481784 235074
rect 481732 235010 481784 235016
rect 477500 234660 477552 234666
rect 477500 234602 477552 234608
rect 476764 234388 476816 234394
rect 476764 234330 476816 234336
rect 475752 4140 475804 4146
rect 475752 4082 475804 4088
rect 475384 3324 475436 3330
rect 475384 3266 475436 3272
rect 474556 3120 474608 3126
rect 474556 3062 474608 3068
rect 474568 480 474596 3062
rect 475764 480 475792 4082
rect 476776 3398 476804 234330
rect 479524 234320 479576 234326
rect 479524 234262 479576 234268
rect 476764 3392 476816 3398
rect 476764 3334 476816 3340
rect 478144 3392 478196 3398
rect 478144 3334 478196 3340
rect 476948 3324 477000 3330
rect 476948 3266 477000 3272
rect 476960 480 476988 3266
rect 478156 480 478184 3334
rect 479536 3330 479564 234262
rect 480536 3392 480588 3398
rect 480536 3334 480588 3340
rect 479524 3324 479576 3330
rect 479524 3266 479576 3272
rect 479340 3256 479392 3262
rect 479340 3198 479392 3204
rect 479352 480 479380 3198
rect 480548 480 480576 3334
rect 481744 480 481772 235010
rect 483676 4146 483704 235078
rect 484412 16574 484440 235146
rect 488552 16574 488580 235894
rect 490564 235884 490616 235890
rect 490564 235826 490616 235832
rect 490012 234252 490064 234258
rect 490012 234194 490064 234200
rect 484412 16546 484808 16574
rect 488552 16546 488856 16574
rect 483664 4140 483716 4146
rect 483664 4082 483716 4088
rect 484032 3936 484084 3942
rect 484032 3878 484084 3884
rect 482836 3324 482888 3330
rect 482836 3266 482888 3272
rect 482848 480 482876 3266
rect 484044 480 484072 3878
rect 484780 490 484808 16546
rect 486424 4956 486476 4962
rect 486424 4898 486476 4904
rect 485056 598 485268 626
rect 485056 490 485084 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 462 485084 490
rect 485240 480 485268 598
rect 486436 480 486464 4898
rect 487620 3868 487672 3874
rect 487620 3810 487672 3816
rect 487632 480 487660 3810
rect 488828 480 488856 16546
rect 490024 6914 490052 234194
rect 489932 6886 490052 6914
rect 489932 480 489960 6886
rect 490576 2922 490604 235826
rect 493324 235816 493376 235822
rect 493324 235758 493376 235764
rect 492680 234184 492732 234190
rect 492680 234126 492732 234132
rect 492692 16574 492720 234126
rect 492692 16546 493088 16574
rect 492312 4140 492364 4146
rect 492312 4082 492364 4088
rect 491116 4004 491168 4010
rect 491116 3946 491168 3952
rect 490564 2916 490616 2922
rect 490564 2858 490616 2864
rect 491128 480 491156 3946
rect 492324 480 492352 4082
rect 493060 490 493088 16546
rect 493336 3330 493364 235758
rect 497464 235748 497516 235754
rect 497464 235690 497516 235696
rect 496820 234116 496872 234122
rect 496820 234058 496872 234064
rect 496832 16574 496860 234058
rect 496832 16546 497136 16574
rect 494704 3800 494756 3806
rect 494704 3742 494756 3748
rect 493324 3324 493376 3330
rect 493324 3266 493376 3272
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 3742
rect 495900 2916 495952 2922
rect 495900 2858 495952 2864
rect 495912 480 495940 2858
rect 497108 480 497136 16546
rect 497476 3942 497504 235690
rect 500224 235680 500276 235686
rect 500224 235622 500276 235628
rect 499580 231192 499632 231198
rect 499580 231134 499632 231140
rect 499592 6914 499620 231134
rect 500236 16574 500264 235622
rect 501604 235612 501656 235618
rect 501604 235554 501656 235560
rect 500236 16546 500356 16574
rect 499592 6886 500264 6914
rect 497464 3936 497516 3942
rect 497464 3878 497516 3884
rect 498200 3732 498252 3738
rect 498200 3674 498252 3680
rect 498212 480 498240 3674
rect 500236 3482 500264 6886
rect 500328 3874 500356 16546
rect 500316 3868 500368 3874
rect 500316 3810 500368 3816
rect 501616 3738 501644 235554
rect 502340 235544 502392 235550
rect 502340 235486 502392 235492
rect 502352 16574 502380 235486
rect 506480 235476 506532 235482
rect 506480 235418 506532 235424
rect 503720 234048 503772 234054
rect 503720 233990 503772 233996
rect 502352 16546 503024 16574
rect 501604 3732 501656 3738
rect 501604 3674 501656 3680
rect 501788 3664 501840 3670
rect 501788 3606 501840 3612
rect 500236 3454 500632 3482
rect 499396 3324 499448 3330
rect 499396 3266 499448 3272
rect 499408 480 499436 3266
rect 500604 480 500632 3454
rect 501800 480 501828 3606
rect 502996 480 503024 16546
rect 503732 490 503760 233990
rect 505376 3596 505428 3602
rect 505376 3538 505428 3544
rect 504008 598 504220 626
rect 504008 490 504036 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 462 504036 490
rect 504192 480 504220 598
rect 505388 480 505416 3538
rect 506492 480 506520 235418
rect 508504 235408 508556 235414
rect 508504 235350 508556 235356
rect 506572 233980 506624 233986
rect 506572 233922 506624 233928
rect 506584 16574 506612 233922
rect 506584 16546 507256 16574
rect 507228 490 507256 16546
rect 508516 3602 508544 235350
rect 512644 235340 512696 235346
rect 512644 235282 512696 235288
rect 510620 232756 510672 232762
rect 510620 232698 510672 232704
rect 510632 16574 510660 232698
rect 510632 16546 511304 16574
rect 510068 3936 510120 3942
rect 510068 3878 510120 3884
rect 508504 3596 508556 3602
rect 508504 3538 508556 3544
rect 508872 3528 508924 3534
rect 508872 3470 508924 3476
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 3470
rect 510080 480 510108 3878
rect 511276 480 511304 16546
rect 512656 3466 512684 235282
rect 520280 235272 520332 235278
rect 520280 235214 520332 235220
rect 519544 233912 519596 233918
rect 519544 233854 519596 233860
rect 514760 231124 514812 231130
rect 514760 231066 514812 231072
rect 513564 3732 513616 3738
rect 513564 3674 513616 3680
rect 512460 3460 512512 3466
rect 512460 3402 512512 3408
rect 512644 3460 512696 3466
rect 512644 3402 512696 3408
rect 512472 480 512500 3402
rect 513576 480 513604 3674
rect 514772 480 514800 231066
rect 517520 177336 517572 177342
rect 517520 177278 517572 177284
rect 517532 16574 517560 177278
rect 519556 16574 519584 233854
rect 517532 16546 517928 16574
rect 519556 16546 519676 16574
rect 515954 3768 516010 3777
rect 515954 3703 516010 3712
rect 515968 480 515996 3703
rect 517152 3664 517204 3670
rect 517152 3606 517204 3612
rect 517164 480 517192 3606
rect 517900 490 517928 16546
rect 519542 3632 519598 3641
rect 519542 3567 519598 3576
rect 518176 598 518388 626
rect 518176 490 518204 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 3567
rect 519648 3534 519676 16546
rect 519636 3528 519688 3534
rect 519636 3470 519688 3476
rect 520292 490 520320 235214
rect 521660 232688 521712 232694
rect 521660 232630 521712 232636
rect 521672 16574 521700 232630
rect 524420 232620 524472 232626
rect 524420 232562 524472 232568
rect 524432 16574 524460 232562
rect 528560 232552 528612 232558
rect 528560 232494 528612 232500
rect 521672 16546 521884 16574
rect 524432 16546 525472 16574
rect 520568 598 520780 626
rect 520568 490 520596 598
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 462 520596 490
rect 520752 480 520780 598
rect 521856 480 521884 16546
rect 524236 3596 524288 3602
rect 524236 3538 524288 3544
rect 523038 3496 523094 3505
rect 523038 3431 523094 3440
rect 523052 480 523080 3431
rect 524248 480 524276 3538
rect 525444 480 525472 16546
rect 527824 3460 527876 3466
rect 527824 3402 527876 3408
rect 526626 3360 526682 3369
rect 526626 3295 526682 3304
rect 526640 480 526668 3295
rect 527836 480 527864 3402
rect 528572 490 528600 232494
rect 530584 175976 530636 175982
rect 530584 175918 530636 175924
rect 530122 3904 530178 3913
rect 530122 3839 530178 3848
rect 528848 598 529060 626
rect 528848 490 528876 598
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 462 528876 490
rect 529032 480 529060 598
rect 530136 480 530164 3839
rect 530596 3534 530624 175918
rect 533710 4856 533766 4865
rect 533710 4791 533766 4800
rect 530584 3528 530636 3534
rect 530584 3470 530636 3476
rect 532516 3528 532568 3534
rect 532516 3470 532568 3476
rect 531320 3460 531372 3466
rect 531320 3402 531372 3408
rect 531332 480 531360 3402
rect 532528 480 532556 3470
rect 533724 480 533752 4791
rect 534908 3596 534960 3602
rect 534908 3538 534960 3544
rect 534920 480 534948 3538
rect 536104 3528 536156 3534
rect 536104 3470 536156 3476
rect 536116 480 536144 3470
rect 536852 3346 536880 337146
rect 536932 332240 536984 332246
rect 536932 332182 536984 332188
rect 536944 3602 536972 332182
rect 537022 330576 537078 330585
rect 537022 330511 537078 330520
rect 536932 3596 536984 3602
rect 536932 3538 536984 3544
rect 537036 3534 537064 330511
rect 537116 322244 537168 322250
rect 537116 322186 537168 322192
rect 537128 239193 537156 322186
rect 537208 321632 537260 321638
rect 537208 321574 537260 321580
rect 537220 239698 537248 321574
rect 537496 299470 537524 387806
rect 538312 337408 538364 337414
rect 538312 337350 538364 337356
rect 538220 337136 538272 337142
rect 538220 337078 538272 337084
rect 537484 299464 537536 299470
rect 537484 299406 537536 299412
rect 537208 239692 537260 239698
rect 537208 239634 537260 239640
rect 537114 239184 537170 239193
rect 537114 239119 537170 239128
rect 538232 16574 538260 337078
rect 538324 316577 538352 337350
rect 538864 337068 538916 337074
rect 538864 337010 538916 337016
rect 538310 316568 538366 316577
rect 538310 316503 538366 316512
rect 538310 256592 538366 256601
rect 538310 256527 538366 256536
rect 538324 237969 538352 256527
rect 538494 254960 538550 254969
rect 538494 254895 538550 254904
rect 538402 253600 538458 253609
rect 538402 253535 538458 253544
rect 538416 238105 538444 253535
rect 538508 239970 538536 254895
rect 538496 239964 538548 239970
rect 538496 239906 538548 239912
rect 538402 238096 538458 238105
rect 538402 238031 538458 238040
rect 538310 237960 538366 237969
rect 538310 237895 538366 237904
rect 538232 16546 538444 16574
rect 537024 3528 537076 3534
rect 537024 3470 537076 3476
rect 536852 3318 537248 3346
rect 537220 480 537248 3318
rect 538416 480 538444 16546
rect 538876 3194 538904 337010
rect 538956 337000 539008 337006
rect 538956 336942 539008 336948
rect 538968 3466 538996 336942
rect 540256 20670 540284 389399
rect 540336 332172 540388 332178
rect 540336 332114 540388 332120
rect 540244 20664 540296 20670
rect 540244 20606 540296 20612
rect 540348 3534 540376 332114
rect 540440 273222 540468 390390
rect 544476 390380 544528 390386
rect 544476 390322 544528 390328
rect 543094 389600 543150 389609
rect 543094 389535 543150 389544
rect 543004 332104 543056 332110
rect 543004 332046 543056 332052
rect 542360 329792 542412 329798
rect 542360 329734 542412 329740
rect 540428 273216 540480 273222
rect 540428 273158 540480 273164
rect 542372 16574 542400 329734
rect 542372 16546 542768 16574
rect 540336 3528 540388 3534
rect 540336 3470 540388 3476
rect 541992 3528 542044 3534
rect 541992 3470 542044 3476
rect 538956 3460 539008 3466
rect 538956 3402 539008 3408
rect 539600 3460 539652 3466
rect 539600 3402 539652 3408
rect 538864 3188 538916 3194
rect 538864 3130 538916 3136
rect 539612 480 539640 3402
rect 540796 3188 540848 3194
rect 540796 3130 540848 3136
rect 540808 480 540836 3130
rect 542004 480 542032 3470
rect 542740 490 542768 16546
rect 543016 3194 543044 332046
rect 543108 179382 543136 389535
rect 543740 336932 543792 336938
rect 543740 336874 543792 336880
rect 543096 179376 543148 179382
rect 543096 179318 543148 179324
rect 543752 16574 543780 336874
rect 544384 329724 544436 329730
rect 544384 329666 544436 329672
rect 543752 16546 544332 16574
rect 544304 3482 544332 16546
rect 544396 4078 544424 329666
rect 544488 259418 544516 390322
rect 547236 390312 547288 390318
rect 547236 390254 547288 390260
rect 547144 332036 547196 332042
rect 547144 331978 547196 331984
rect 546500 329656 546552 329662
rect 546500 329598 546552 329604
rect 544476 259412 544528 259418
rect 544476 259354 544528 259360
rect 546512 16574 546540 329598
rect 546512 16546 546724 16574
rect 544384 4072 544436 4078
rect 544384 4014 544436 4020
rect 544304 3454 544424 3482
rect 543004 3188 543056 3194
rect 543004 3130 543056 3136
rect 543016 598 543228 626
rect 543016 490 543044 598
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 462 543044 490
rect 543200 480 543228 598
rect 544396 480 544424 3454
rect 545488 3188 545540 3194
rect 545488 3130 545540 3136
rect 545500 480 545528 3130
rect 546696 480 546724 16546
rect 547156 4146 547184 331978
rect 547248 313274 547276 390254
rect 569314 389328 569370 389337
rect 569314 389263 569370 389272
rect 555424 386980 555476 386986
rect 555424 386922 555476 386928
rect 547970 335336 548026 335345
rect 547970 335271 548026 335280
rect 547236 313268 547288 313274
rect 547236 313210 547288 313216
rect 547984 6914 548012 335271
rect 550638 335200 550694 335209
rect 550638 335135 550694 335144
rect 548524 331968 548576 331974
rect 548524 331910 548576 331916
rect 547892 6886 548012 6914
rect 547144 4140 547196 4146
rect 547144 4082 547196 4088
rect 547892 480 547920 6886
rect 548536 3534 548564 331910
rect 550652 16574 550680 335135
rect 554780 334620 554832 334626
rect 554780 334562 554832 334568
rect 551282 332480 551338 332489
rect 551282 332415 551338 332424
rect 550652 16546 551048 16574
rect 549076 4140 549128 4146
rect 549076 4082 549128 4088
rect 548524 3528 548576 3534
rect 548524 3470 548576 3476
rect 549088 480 549116 4082
rect 550272 4072 550324 4078
rect 550272 4014 550324 4020
rect 550284 480 550312 4014
rect 551020 490 551048 16546
rect 551296 3670 551324 332415
rect 553400 329588 553452 329594
rect 553400 329530 553452 329536
rect 553412 16574 553440 329530
rect 554792 16574 554820 334562
rect 555436 60722 555464 386922
rect 557540 336864 557592 336870
rect 557540 336806 557592 336812
rect 556160 331900 556212 331906
rect 556160 331842 556212 331848
rect 555424 60716 555476 60722
rect 555424 60658 555476 60664
rect 553412 16546 553808 16574
rect 554792 16546 555004 16574
rect 551284 3664 551336 3670
rect 551284 3606 551336 3612
rect 552664 3528 552716 3534
rect 552664 3470 552716 3476
rect 551296 598 551508 626
rect 551296 490 551324 598
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 462 551324 490
rect 551480 480 551508 598
rect 552676 480 552704 3470
rect 553780 480 553808 16546
rect 554976 480 555004 16546
rect 556172 480 556200 331842
rect 556252 329452 556304 329458
rect 556252 329394 556304 329400
rect 556264 16574 556292 329394
rect 556264 16546 556936 16574
rect 556908 490 556936 16546
rect 557552 6914 557580 336806
rect 561680 336796 561732 336802
rect 561680 336738 561732 336744
rect 558182 332344 558238 332353
rect 558182 332279 558238 332288
rect 558196 16574 558224 332279
rect 560300 329520 560352 329526
rect 560300 329462 560352 329468
rect 560312 16574 560340 329462
rect 561692 16574 561720 336738
rect 564438 335064 564494 335073
rect 564438 334999 564494 335008
rect 562322 332208 562378 332217
rect 562322 332143 562378 332152
rect 558196 16546 558316 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 557552 6886 558224 6914
rect 558196 2802 558224 6886
rect 558288 2922 558316 16546
rect 559748 3664 559800 3670
rect 559748 3606 559800 3612
rect 558276 2916 558328 2922
rect 558276 2858 558328 2864
rect 558196 2774 558592 2802
rect 557184 598 557396 626
rect 557184 490 557212 598
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 462 557212 490
rect 557368 480 557396 598
rect 558564 480 558592 2774
rect 559760 480 559788 3606
rect 560404 490 560432 16546
rect 560680 598 560892 626
rect 560680 490 560708 598
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560404 462 560708 490
rect 560864 480 560892 598
rect 562060 480 562088 16546
rect 562336 3534 562364 332143
rect 564452 3602 564480 334999
rect 568578 334928 568634 334937
rect 568578 334863 568634 334872
rect 564532 329384 564584 329390
rect 564532 329326 564584 329332
rect 564440 3596 564492 3602
rect 564440 3538 564492 3544
rect 562324 3528 562376 3534
rect 564544 3482 564572 329326
rect 566464 329316 566516 329322
rect 566464 329258 566516 329264
rect 566476 4146 566504 329258
rect 568592 16574 568620 334863
rect 569222 332072 569278 332081
rect 569222 332007 569278 332016
rect 568592 16546 568712 16574
rect 566464 4140 566516 4146
rect 566464 4082 566516 4088
rect 568028 4140 568080 4146
rect 568028 4082 568080 4088
rect 565636 3596 565688 3602
rect 565636 3538 565688 3544
rect 562324 3470 562376 3476
rect 564452 3454 564572 3482
rect 563244 2916 563296 2922
rect 563244 2858 563296 2864
rect 563256 480 563284 2858
rect 564452 480 564480 3454
rect 565648 480 565676 3538
rect 566832 3528 566884 3534
rect 566832 3470 566884 3476
rect 566844 480 566872 3470
rect 568040 480 568068 4082
rect 568684 490 568712 16546
rect 569236 3330 569264 332007
rect 569328 100706 569356 389263
rect 573362 389192 573418 389201
rect 573362 389127 573418 389136
rect 572718 334792 572774 334801
rect 572718 334727 572774 334736
rect 571340 329248 571392 329254
rect 571340 329190 571392 329196
rect 569316 100700 569368 100706
rect 569316 100642 569368 100648
rect 571352 16574 571380 329190
rect 571352 16546 571564 16574
rect 569224 3324 569276 3330
rect 569224 3266 569276 3272
rect 570328 3324 570380 3330
rect 570328 3266 570380 3272
rect 568960 598 569172 626
rect 568960 490 568988 598
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 462 568988 490
rect 569144 480 569172 598
rect 570340 480 570368 3266
rect 571536 480 571564 16546
rect 572732 480 572760 334727
rect 572810 331936 572866 331945
rect 572810 331871 572866 331880
rect 572824 16574 572852 331871
rect 573376 139398 573404 389127
rect 580356 387184 580408 387190
rect 580356 387126 580408 387132
rect 580264 386504 580316 386510
rect 580264 386446 580316 386452
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 575478 334656 575534 334665
rect 575478 334591 575534 334600
rect 574742 331800 574798 331809
rect 574742 331735 574798 331744
rect 574100 329180 574152 329186
rect 574100 329122 574152 329128
rect 573364 139392 573416 139398
rect 573364 139334 573416 139340
rect 572824 16546 573496 16574
rect 573468 490 573496 16546
rect 574112 6914 574140 329122
rect 574756 16574 574784 331735
rect 575492 16574 575520 334591
rect 576124 329112 576176 329118
rect 576124 329054 576176 329060
rect 574756 16546 574876 16574
rect 575492 16546 575888 16574
rect 574112 6886 574784 6914
rect 574756 3482 574784 6886
rect 574848 3602 574876 16546
rect 574836 3596 574888 3602
rect 574836 3538 574888 3544
rect 574756 3454 575152 3482
rect 573744 598 573956 626
rect 573744 490 573772 598
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573468 462 573772 490
rect 573928 480 573956 598
rect 575124 480 575152 3454
rect 575860 490 575888 16546
rect 576136 3806 576164 329054
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 579988 273216 580040 273222
rect 579988 273158 580040 273164
rect 580000 272241 580028 273158
rect 579986 272232 580042 272241
rect 579986 272167 580042 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579620 179376 579672 179382
rect 579620 179318 579672 179324
rect 579632 179217 579660 179318
rect 579618 179208 579674 179217
rect 579618 179143 579674 179152
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580276 112849 580304 386446
rect 580368 126041 580396 387126
rect 580908 386912 580960 386918
rect 580908 386854 580960 386860
rect 580724 386844 580776 386850
rect 580724 386786 580776 386792
rect 580632 386708 580684 386714
rect 580632 386650 580684 386656
rect 580448 386640 580500 386646
rect 580448 386582 580500 386588
rect 580460 152697 580488 386582
rect 580540 386572 580592 386578
rect 580540 386514 580592 386520
rect 580552 165889 580580 386514
rect 580644 205737 580672 386650
rect 580736 351937 580764 386786
rect 580816 386776 580868 386782
rect 580816 386718 580868 386724
rect 580722 351928 580778 351937
rect 580722 351863 580778 351872
rect 580724 334688 580776 334694
rect 580724 334630 580776 334636
rect 580630 205728 580686 205737
rect 580630 205663 580686 205672
rect 580736 192545 580764 334630
rect 580828 245585 580856 386718
rect 580920 378457 580948 386854
rect 580906 378448 580962 378457
rect 580906 378383 580962 378392
rect 580908 337544 580960 337550
rect 580908 337486 580960 337492
rect 580814 245576 580870 245585
rect 580814 245511 580870 245520
rect 580920 232393 580948 337486
rect 581000 320884 581052 320890
rect 581000 320826 581052 320832
rect 580906 232384 580962 232393
rect 580906 232319 580962 232328
rect 580722 192536 580778 192545
rect 580722 192471 580778 192480
rect 580538 165880 580594 165889
rect 580538 165815 580594 165824
rect 580446 152688 580502 152697
rect 580446 152623 580502 152632
rect 580354 126032 580410 126041
rect 580354 125967 580410 125976
rect 580262 112840 580318 112849
rect 580262 112775 580318 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 576124 3800 576176 3806
rect 576124 3742 576176 3748
rect 578608 3800 578660 3806
rect 578608 3742 578660 3748
rect 577412 3596 577464 3602
rect 577412 3538 577464 3544
rect 576136 598 576348 626
rect 576136 490 576164 598
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 462 576164 490
rect 576320 480 576348 598
rect 577424 480 577452 3538
rect 578620 480 578648 3742
rect 581012 480 581040 320826
rect 582196 4888 582248 4894
rect 582196 4830 582248 4836
rect 582208 480 582236 4830
rect 583392 2848 583444 2854
rect 583392 2790 583444 2796
rect 583404 480 583432 2790
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 3146 410488 3202 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3054 293120 3110 293176
rect 3146 254088 3202 254144
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3238 162832 3294 162888
rect 3146 110608 3202 110664
rect 2778 71612 2780 71632
rect 2780 71612 2832 71632
rect 2832 71612 2834 71632
rect 2778 71576 2834 71612
rect 3054 58520 3110 58576
rect 3514 345344 3570 345400
rect 3514 319232 3570 319288
rect 3514 306176 3570 306232
rect 3514 267144 3570 267200
rect 3514 241032 3570 241088
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3422 32408 3478 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 15106 335960 15162 336016
rect 15198 335552 15254 335608
rect 16578 334600 16634 334656
rect 24858 335416 24914 335472
rect 28998 333240 29054 333296
rect 25502 330384 25558 330440
rect 31666 336232 31722 336288
rect 32402 333376 32458 333432
rect 33046 336368 33102 336424
rect 36542 331744 36598 331800
rect 38566 336504 38622 336560
rect 39302 331880 39358 331936
rect 40682 333512 40738 333568
rect 50986 336640 51042 336696
rect 43442 332016 43498 332072
rect 48226 333648 48282 333704
rect 57886 335824 57942 335880
rect 55126 334736 55182 334792
rect 53102 332152 53158 332208
rect 62026 330656 62082 330712
rect 61382 330520 61438 330576
rect 66166 332288 66222 332344
rect 70306 330792 70362 330848
rect 81346 333784 81402 333840
rect 140686 335144 140742 335200
rect 136454 335008 136510 335064
rect 129646 334872 129702 334928
rect 128266 333920 128322 333976
rect 240690 389544 240746 389600
rect 235906 389408 235962 389464
rect 238390 389272 238446 389328
rect 239494 389136 239550 389192
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 233146 386960 233202 387016
rect 232778 385056 232834 385112
rect 232686 379344 232742 379400
rect 232594 373496 232650 373552
rect 232502 363976 232558 364032
rect 232318 358128 232374 358184
rect 232226 352416 232282 352472
rect 232042 342760 232098 342816
rect 158626 335280 158682 335336
rect 231306 334056 231362 334112
rect 232410 356224 232466 356280
rect 232870 381248 232926 381304
rect 233054 377440 233110 377496
rect 232962 375400 233018 375456
rect 232870 346568 232926 346624
rect 234434 383152 234490 383208
rect 234342 371592 234398 371648
rect 234158 369688 234214 369744
rect 234066 365880 234122 365936
rect 233974 361936 234030 361992
rect 233882 360032 233938 360088
rect 233790 354320 233846 354376
rect 233698 350376 233754 350432
rect 233514 344664 233570 344720
rect 233238 338000 233294 338056
rect 233330 337864 233386 337920
rect 233606 340856 233662 340912
rect 233330 330384 233386 330440
rect 233882 238312 233938 238368
rect 234250 367784 234306 367840
rect 234158 238584 234214 238640
rect 234066 238448 234122 238504
rect 233974 237088 234030 237144
rect 234250 236952 234306 237008
rect 234526 348472 234582 348528
rect 234710 338952 234766 339008
rect 234618 336096 234674 336152
rect 234618 333512 234674 333568
rect 234802 333376 234858 333432
rect 234342 236408 234398 236464
rect 234986 336232 235042 336288
rect 235538 337728 235594 337784
rect 235170 331880 235226 331936
rect 235078 331744 235134 331800
rect 235538 335824 235594 335880
rect 235446 332016 235502 332072
rect 236412 337864 236468 337920
rect 236090 335960 236146 336016
rect 236182 335688 236238 335744
rect 236734 335960 236790 336016
rect 236366 335552 236422 335608
rect 236182 334600 236238 334656
rect 236826 335416 236882 335472
rect 236734 334056 236790 334112
rect 236366 333784 236422 333840
rect 236642 333784 236698 333840
rect 236366 333512 236422 333568
rect 235354 238856 235410 238912
rect 237010 335416 237066 335472
rect 237010 333240 237066 333296
rect 236918 333104 236974 333160
rect 237378 335416 237434 335472
rect 237470 333376 237526 333432
rect 238528 337864 238584 337920
rect 237654 336368 237710 336424
rect 238022 336504 238078 336560
rect 237838 334056 237894 334112
rect 237930 333512 237986 333568
rect 236734 238720 236790 238776
rect 238206 333648 238262 333704
rect 238298 333376 238354 333432
rect 238298 332560 238354 332616
rect 238758 336640 238814 336696
rect 239448 337864 239504 337920
rect 239632 337864 239688 337920
rect 239816 337864 239872 337920
rect 239494 337592 239550 337648
rect 239218 332152 239274 332208
rect 239862 337728 239918 337784
rect 240138 335280 240194 335336
rect 239954 330656 240010 330712
rect 239770 330520 239826 330576
rect 240414 332288 240470 332344
rect 241196 337864 241252 337920
rect 240966 337592 241022 337648
rect 241150 337592 241206 337648
rect 241242 335960 241298 336016
rect 241150 330792 241206 330848
rect 242024 337830 242080 337886
rect 242208 337864 242264 337920
rect 241886 337456 241942 337512
rect 242254 337728 242310 337784
rect 242944 337864 243000 337920
rect 242898 337728 242954 337784
rect 243174 337728 243230 337784
rect 242806 336096 242862 336152
rect 243358 333784 243414 333840
rect 244048 337830 244104 337886
rect 243726 337456 243782 337512
rect 244094 337592 244150 337648
rect 244554 337728 244610 337784
rect 244876 337864 244932 337920
rect 244554 335008 244610 335064
rect 245704 337864 245760 337920
rect 245198 333920 245254 333976
rect 245474 334908 245476 334928
rect 245476 334908 245528 334928
rect 245528 334908 245530 334928
rect 245474 334872 245530 334908
rect 246072 337864 246128 337920
rect 246256 337864 246312 337920
rect 245658 337592 245714 337648
rect 245474 332560 245530 332616
rect 245934 337592 245990 337648
rect 246394 335144 246450 335200
rect 246992 337728 247048 337784
rect 247360 337830 247416 337886
rect 247728 337864 247784 337920
rect 247406 337456 247462 337512
rect 247590 337456 247646 337512
rect 247912 337830 247968 337886
rect 247958 337592 248014 337648
rect 249384 337864 249440 337920
rect 248602 334056 248658 334112
rect 249246 333240 249302 333296
rect 249430 337728 249486 337784
rect 249936 337898 249992 337954
rect 249890 337728 249946 337784
rect 249246 236816 249302 236872
rect 251040 337898 251096 337954
rect 251086 337728 251142 337784
rect 252880 337898 252936 337954
rect 252926 337592 252982 337648
rect 254536 337728 254592 337784
rect 254904 337898 254960 337954
rect 255272 337898 255328 337954
rect 255456 337898 255512 337954
rect 254490 337592 254546 337648
rect 254582 335552 254638 335608
rect 254858 337728 254914 337784
rect 255318 337728 255374 337784
rect 255824 337898 255880 337954
rect 255502 337728 255558 337784
rect 255870 337728 255926 337784
rect 254674 238992 254730 239048
rect 256146 335688 256202 335744
rect 256146 330384 256202 330440
rect 256928 337898 256984 337954
rect 256974 337728 257030 337784
rect 257664 337898 257720 337954
rect 257664 337728 257720 337784
rect 258216 337898 258272 337954
rect 258400 337898 258456 337954
rect 258584 337898 258640 337954
rect 258952 337898 259008 337954
rect 258446 337728 258502 337784
rect 258814 337728 258870 337784
rect 259136 337898 259192 337954
rect 259320 337898 259376 337954
rect 259504 337898 259560 337954
rect 259366 337728 259422 337784
rect 259550 337728 259606 337784
rect 258998 337592 259054 337648
rect 259090 337456 259146 337512
rect 259182 337320 259238 337376
rect 263552 337864 263608 337920
rect 263690 337728 263746 337784
rect 264288 337898 264344 337954
rect 264656 337898 264712 337954
rect 264840 337898 264896 337954
rect 264794 337728 264850 337784
rect 264978 337728 265034 337784
rect 266128 337830 266184 337886
rect 266082 337592 266138 337648
rect 268704 337898 268760 337954
rect 268888 337864 268944 337920
rect 269026 337728 269082 337784
rect 269256 337864 269312 337920
rect 269624 337864 269680 337920
rect 268566 337456 268622 337512
rect 269026 336504 269082 336560
rect 269670 337592 269726 337648
rect 269854 336232 269910 336288
rect 270360 337864 270416 337920
rect 270130 337456 270186 337512
rect 270130 333784 270186 333840
rect 270406 337728 270462 337784
rect 270728 337864 270784 337920
rect 270406 336096 270462 336152
rect 271188 337864 271244 337920
rect 270590 335960 270646 336016
rect 270774 337456 270830 337512
rect 270314 333648 270370 333704
rect 270406 330792 270462 330848
rect 270590 330656 270646 330712
rect 270774 333512 270830 333568
rect 271510 337728 271566 337784
rect 272108 337864 272164 337920
rect 271786 333240 271842 333296
rect 272936 337898 272992 337954
rect 272430 333376 272486 333432
rect 272890 337728 272946 337784
rect 273120 337830 273176 337886
rect 272706 239808 272762 239864
rect 273074 337592 273130 337648
rect 273166 336368 273222 336424
rect 273442 335144 273498 335200
rect 274500 337864 274556 337920
rect 273718 239400 273774 239456
rect 274960 337898 275016 337954
rect 274638 337456 274694 337512
rect 274362 335144 274418 335200
rect 274822 335688 274878 335744
rect 275880 337898 275936 337954
rect 276064 337898 276120 337954
rect 276248 337898 276304 337954
rect 275926 337728 275982 337784
rect 276202 337728 276258 337784
rect 275190 239672 275246 239728
rect 275834 337456 275890 337512
rect 276708 337898 276764 337954
rect 276294 337592 276350 337648
rect 276386 239536 276442 239592
rect 276984 337898 277040 337954
rect 277122 337728 277178 337784
rect 277122 337320 277178 337376
rect 277904 337864 277960 337920
rect 277490 336368 277546 336424
rect 277490 335824 277546 335880
rect 277950 337728 278006 337784
rect 278272 337864 278328 337920
rect 278456 337898 278512 337954
rect 278824 337898 278880 337954
rect 279008 337898 279064 337954
rect 277858 337592 277914 337648
rect 277950 334736 278006 334792
rect 277582 4800 277638 4856
rect 278962 337592 279018 337648
rect 279422 337592 279478 337648
rect 279836 337864 279892 337920
rect 280388 337898 280444 337954
rect 279238 330520 279294 330576
rect 279882 335280 279938 335336
rect 280664 337830 280720 337886
rect 280434 337592 280490 337648
rect 280066 335144 280122 335200
rect 280434 332424 280490 332480
rect 280710 332288 280766 332344
rect 279330 3304 279386 3360
rect 280894 335688 280950 335744
rect 281400 337830 281456 337886
rect 281262 337592 281318 337648
rect 281170 335008 281226 335064
rect 281446 334872 281502 334928
rect 281354 332152 281410 332208
rect 282320 337864 282376 337920
rect 282596 337898 282652 337954
rect 282550 337728 282606 337784
rect 281630 332016 281686 332072
rect 282274 337456 282330 337512
rect 281906 334736 281962 334792
rect 281998 331880 282054 331936
rect 282366 336640 282422 336696
rect 282274 335416 282330 335472
rect 282182 334600 282238 334656
rect 282366 331744 282422 331800
rect 282642 334056 282698 334112
rect 283240 337898 283296 337954
rect 283424 337864 283480 337920
rect 283378 337592 283434 337648
rect 282918 336504 282974 336560
rect 283010 334192 283066 334248
rect 282918 334056 282974 334112
rect 284160 337898 284216 337954
rect 283976 337830 284032 337886
rect 284114 337728 284170 337784
rect 283930 337592 283986 337648
rect 284620 337864 284676 337920
rect 284390 335552 284446 335608
rect 285494 337864 285550 337920
rect 286322 335824 286378 335880
rect 285586 334212 285642 334248
rect 285586 334192 285588 334212
rect 285588 334192 285640 334212
rect 285640 334192 285642 334212
rect 287426 382200 287482 382256
rect 287426 377304 287482 377360
rect 287610 375808 287666 375864
rect 287794 372544 287850 372600
rect 287610 370912 287666 370968
rect 287978 367648 288034 367704
rect 287610 366016 287666 366072
rect 287610 362888 287666 362944
rect 287610 361256 287666 361312
rect 287610 359624 287666 359680
rect 287794 356360 287850 356416
rect 287518 353096 287574 353152
rect 287242 351484 287298 351520
rect 287242 351464 287244 351484
rect 287244 351464 287296 351484
rect 287296 351464 287298 351484
rect 287978 348336 288034 348392
rect 287978 346704 288034 346760
rect 287794 340176 287850 340232
rect 287426 338680 287482 338736
rect 287610 338136 287666 338192
rect 287334 337456 287390 337512
rect 286874 337320 286930 337376
rect 286782 335416 286838 335472
rect 288346 387096 288402 387152
rect 288346 385464 288402 385520
rect 288346 383832 288402 383888
rect 288346 380568 288402 380624
rect 288346 378936 288402 378992
rect 288346 374196 288402 374232
rect 288346 374176 288348 374196
rect 288348 374176 288400 374196
rect 288400 374176 288402 374196
rect 288346 369280 288402 369336
rect 288346 364404 288402 364440
rect 288346 364384 288348 364404
rect 288348 364384 288400 364404
rect 288400 364384 288402 364404
rect 288346 357992 288402 358048
rect 288346 354748 288402 354784
rect 288346 354728 288348 354748
rect 288348 354728 288400 354748
rect 288400 354728 288402 354748
rect 288346 349968 288402 350024
rect 288346 345092 288402 345128
rect 288346 345072 288348 345092
rect 288348 345072 288400 345092
rect 288400 345072 288402 345092
rect 288346 343440 288402 343496
rect 288346 341808 288402 341864
rect 289174 3712 289230 3768
rect 290462 334328 290518 334384
rect 293222 238176 293278 238232
rect 293314 236680 293370 236736
rect 290646 3576 290702 3632
rect 290462 3440 290518 3496
rect 297638 236544 297694 236600
rect 304262 336640 304318 336696
rect 304446 336504 304502 336560
rect 398102 336368 398158 336424
rect 416042 336232 416098 336288
rect 412638 333920 412694 333976
rect 418802 333784 418858 333840
rect 420182 336096 420238 336152
rect 422942 335960 422998 336016
rect 427082 334464 427138 334520
rect 423678 333648 423734 333704
rect 432602 333512 432658 333568
rect 427818 330792 427874 330848
rect 427082 3848 427138 3904
rect 436650 272856 436706 272912
rect 436098 267416 436154 267472
rect 436098 247288 436154 247344
rect 436834 271224 436890 271280
rect 436834 270136 436890 270192
rect 437478 274216 437534 274272
rect 437386 272856 437442 272912
rect 437294 268368 437350 268424
rect 437202 265648 437258 265704
rect 436742 245520 436798 245576
rect 437294 238040 437350 238096
rect 437202 237904 437258 237960
rect 438214 333376 438270 333432
rect 439502 333240 439558 333296
rect 438858 330656 438914 330712
rect 438766 274216 438822 274272
rect 438674 271224 438730 271280
rect 438582 270136 438638 270192
rect 540242 389408 540298 389464
rect 467838 322496 467894 322552
rect 469402 322496 469458 322552
rect 474554 322496 474610 322552
rect 476578 322496 476634 322552
rect 479154 322496 479210 322552
rect 481638 322496 481694 322552
rect 483018 322496 483074 322552
rect 484858 322496 484914 322552
rect 470690 321544 470746 321600
rect 471978 321544 472034 321600
rect 472254 321544 472310 321600
rect 475474 321544 475530 321600
rect 478234 321544 478290 321600
rect 480626 321544 480682 321600
rect 519542 330384 519598 330440
rect 488538 322496 488594 322552
rect 490562 322496 490618 322552
rect 492678 322496 492734 322552
rect 485778 321952 485834 322008
rect 484398 321544 484454 321600
rect 519542 322360 519598 322416
rect 488170 321580 488172 321600
rect 488172 321580 488224 321600
rect 488224 321580 488226 321600
rect 488170 321544 488226 321580
rect 492218 321544 492274 321600
rect 494242 321544 494298 321600
rect 495530 321544 495586 321600
rect 496818 321544 496874 321600
rect 498198 321544 498254 321600
rect 498658 321544 498714 321600
rect 500682 321544 500738 321600
rect 501050 321544 501106 321600
rect 503258 321544 503314 321600
rect 504178 321544 504234 321600
rect 505466 321544 505522 321600
rect 506938 321544 506994 321600
rect 530030 321580 530032 321600
rect 530032 321580 530084 321600
rect 530084 321580 530086 321600
rect 530030 321544 530086 321580
rect 439686 237768 439742 237824
rect 445574 239808 445630 239864
rect 445850 239808 445906 239864
rect 451094 239808 451150 239864
rect 452750 239808 452806 239864
rect 460938 239808 460994 239864
rect 522670 239844 522672 239864
rect 522672 239844 522724 239864
rect 522724 239844 522726 239864
rect 522670 239808 522726 239844
rect 523130 239828 523186 239864
rect 523130 239808 523132 239828
rect 523132 239808 523184 239828
rect 523184 239808 523186 239828
rect 462410 239672 462466 239728
rect 473174 239672 473230 239728
rect 475658 239672 475714 239728
rect 523130 239672 523186 239728
rect 445666 239264 445722 239320
rect 451094 239264 451150 239320
rect 452566 239264 452622 239320
rect 461030 239264 461086 239320
rect 445574 239128 445630 239184
rect 452658 239128 452714 239184
rect 462318 237224 462374 237280
rect 461122 236816 461178 236872
rect 465262 239536 465318 239592
rect 471978 239536 472034 239592
rect 463698 237224 463754 237280
rect 465078 237224 465134 237280
rect 465078 236816 465134 236872
rect 468482 239400 468538 239456
rect 467194 237632 467250 237688
rect 467838 237668 467840 237688
rect 467840 237668 467892 237688
rect 467892 237668 467894 237688
rect 467838 237632 467894 237668
rect 467838 237260 467840 237280
rect 467840 237260 467892 237280
rect 467892 237260 467894 237280
rect 467838 237224 467894 237260
rect 479338 239536 479394 239592
rect 487894 239536 487950 239592
rect 495622 239536 495678 239592
rect 496818 239536 496874 239592
rect 500498 239536 500554 239592
rect 501878 239536 501934 239592
rect 503074 239536 503130 239592
rect 477682 238620 477684 238640
rect 477684 238620 477736 238640
rect 477736 238620 477738 238640
rect 477682 238584 477738 238620
rect 483386 238584 483442 238640
rect 484398 238604 484454 238640
rect 484398 238584 484400 238604
rect 484400 238584 484452 238604
rect 484452 238584 484454 238604
rect 485410 238584 485466 238640
rect 482282 238468 482338 238504
rect 482282 238448 482284 238468
rect 482284 238448 482336 238468
rect 482336 238448 482338 238468
rect 484858 238448 484914 238504
rect 476578 238312 476634 238368
rect 480626 238312 480682 238368
rect 481730 238312 481786 238368
rect 485962 238312 486018 238368
rect 488170 238332 488226 238368
rect 488170 238312 488172 238332
rect 488172 238312 488224 238332
rect 488224 238312 488226 238332
rect 491666 238196 491722 238232
rect 491666 238176 491668 238196
rect 491668 238176 491720 238196
rect 491720 238176 491722 238196
rect 492770 238176 492826 238232
rect 495162 238176 495218 238232
rect 505558 239536 505614 239592
rect 506754 239536 506810 239592
rect 469218 237224 469274 237280
rect 470598 237224 470654 237280
rect 485778 237224 485834 237280
rect 498198 237224 498254 237280
rect 503718 237244 503774 237280
rect 503718 237224 503720 237244
rect 503720 237224 503772 237244
rect 503772 237224 503774 237244
rect 521658 237224 521714 237280
rect 490286 237088 490342 237144
rect 492678 237108 492734 237144
rect 492678 237088 492680 237108
rect 492680 237088 492732 237108
rect 492732 237088 492734 237108
rect 494058 237088 494114 237144
rect 491298 236972 491354 237008
rect 491298 236952 491300 236972
rect 491300 236952 491352 236972
rect 491352 236952 491354 236972
rect 471978 236816 472034 236872
rect 473358 236836 473414 236872
rect 473358 236816 473360 236836
rect 473360 236816 473412 236836
rect 473412 236816 473414 236836
rect 474738 236816 474794 236872
rect 476118 236816 476174 236872
rect 485778 236816 485834 236872
rect 488538 236816 488594 236872
rect 470874 236272 470930 236328
rect 469218 236136 469274 236192
rect 477498 236136 477554 236192
rect 495438 236156 495494 236192
rect 495438 236136 495440 236156
rect 495440 236136 495492 236156
rect 495492 236136 495494 236156
rect 515954 3712 516010 3768
rect 519542 3576 519598 3632
rect 523038 3440 523094 3496
rect 526626 3304 526682 3360
rect 530122 3848 530178 3904
rect 533710 4800 533766 4856
rect 537022 330520 537078 330576
rect 537114 239128 537170 239184
rect 538310 316512 538366 316568
rect 538310 256536 538366 256592
rect 538494 254904 538550 254960
rect 538402 253544 538458 253600
rect 538402 238040 538458 238096
rect 538310 237904 538366 237960
rect 543094 389544 543150 389600
rect 569314 389272 569370 389328
rect 547970 335280 548026 335336
rect 550638 335144 550694 335200
rect 551282 332424 551338 332480
rect 558182 332288 558238 332344
rect 564438 335008 564494 335064
rect 562322 332152 562378 332208
rect 568578 334872 568634 334928
rect 569222 332016 569278 332072
rect 573362 389136 573418 389192
rect 572718 334736 572774 334792
rect 572810 331880 572866 331936
rect 580170 365064 580226 365120
rect 575478 334600 575534 334656
rect 574742 331744 574798 331800
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 579986 272176 580042 272232
rect 580170 258848 580226 258904
rect 580170 219000 580226 219056
rect 579618 179152 579674 179208
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580722 351872 580778 351928
rect 580630 205672 580686 205728
rect 580906 378392 580962 378448
rect 580814 245520 580870 245576
rect 580906 232328 580962 232384
rect 580722 192480 580778 192536
rect 580538 165824 580594 165880
rect 580446 152632 580502 152688
rect 580354 125976 580410 126032
rect 580262 112784 580318 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 583520 391628 584960 391868
rect 240685 389602 240751 389605
rect 543089 389602 543155 389605
rect 240685 389600 543155 389602
rect 240685 389544 240690 389600
rect 240746 389544 543094 389600
rect 543150 389544 543155 389600
rect 240685 389542 543155 389544
rect 240685 389539 240751 389542
rect 543089 389539 543155 389542
rect 235901 389466 235967 389469
rect 540237 389466 540303 389469
rect 235901 389464 540303 389466
rect 235901 389408 235906 389464
rect 235962 389408 540242 389464
rect 540298 389408 540303 389464
rect 235901 389406 540303 389408
rect 235901 389403 235967 389406
rect 540237 389403 540303 389406
rect 238385 389330 238451 389333
rect 569309 389330 569375 389333
rect 238385 389328 569375 389330
rect 238385 389272 238390 389328
rect 238446 389272 569314 389328
rect 569370 389272 569375 389328
rect 238385 389270 569375 389272
rect 238385 389267 238451 389270
rect 569309 389267 569375 389270
rect 239489 389194 239555 389197
rect 573357 389194 573423 389197
rect 239489 389192 573423 389194
rect 239489 389136 239494 389192
rect 239550 389136 573362 389192
rect 573418 389136 573423 389192
rect 239489 389134 573423 389136
rect 239489 389131 239555 389134
rect 573357 389131 573423 389134
rect 288341 387154 288407 387157
rect 284924 387152 288407 387154
rect 284924 387096 288346 387152
rect 288402 387096 288407 387152
rect 284924 387094 288407 387096
rect 288341 387091 288407 387094
rect 233141 387018 233207 387021
rect 233141 387016 235060 387018
rect 233141 386960 233146 387016
rect 233202 386960 235060 387016
rect 233141 386958 235060 386960
rect 233141 386955 233207 386958
rect 288341 385522 288407 385525
rect 284924 385520 288407 385522
rect 284924 385464 288346 385520
rect 288402 385464 288407 385520
rect 284924 385462 288407 385464
rect 288341 385459 288407 385462
rect 232773 385114 232839 385117
rect 232773 385112 235060 385114
rect 232773 385056 232778 385112
rect 232834 385056 235060 385112
rect 232773 385054 235060 385056
rect 232773 385051 232839 385054
rect -960 384284 480 384524
rect 288341 383890 288407 383893
rect 284924 383888 288407 383890
rect 284924 383832 288346 383888
rect 288402 383832 288407 383888
rect 284924 383830 288407 383832
rect 288341 383827 288407 383830
rect 234429 383210 234495 383213
rect 234429 383208 235060 383210
rect 234429 383152 234434 383208
rect 234490 383152 235060 383208
rect 234429 383150 235060 383152
rect 234429 383147 234495 383150
rect 287421 382258 287487 382261
rect 284924 382256 287487 382258
rect 284924 382200 287426 382256
rect 287482 382200 287487 382256
rect 284924 382198 287487 382200
rect 287421 382195 287487 382198
rect 232865 381306 232931 381309
rect 232865 381304 235060 381306
rect 232865 381248 232870 381304
rect 232926 381248 235060 381304
rect 232865 381246 235060 381248
rect 232865 381243 232931 381246
rect 288341 380626 288407 380629
rect 284924 380624 288407 380626
rect 284924 380568 288346 380624
rect 288402 380568 288407 380624
rect 284924 380566 288407 380568
rect 288341 380563 288407 380566
rect 232681 379402 232747 379405
rect 232681 379400 235060 379402
rect 232681 379344 232686 379400
rect 232742 379344 235060 379400
rect 232681 379342 235060 379344
rect 232681 379339 232747 379342
rect 288341 378994 288407 378997
rect 284924 378992 288407 378994
rect 284924 378936 288346 378992
rect 288402 378936 288407 378992
rect 284924 378934 288407 378936
rect 288341 378931 288407 378934
rect 580901 378450 580967 378453
rect 583520 378450 584960 378540
rect 580901 378448 584960 378450
rect 580901 378392 580906 378448
rect 580962 378392 584960 378448
rect 580901 378390 584960 378392
rect 580901 378387 580967 378390
rect 583520 378300 584960 378390
rect 233049 377498 233115 377501
rect 233049 377496 235060 377498
rect 233049 377440 233054 377496
rect 233110 377440 235060 377496
rect 233049 377438 235060 377440
rect 233049 377435 233115 377438
rect 287421 377362 287487 377365
rect 284924 377360 287487 377362
rect 284924 377304 287426 377360
rect 287482 377304 287487 377360
rect 284924 377302 287487 377304
rect 287421 377299 287487 377302
rect 287605 375866 287671 375869
rect 284924 375864 287671 375866
rect 284924 375808 287610 375864
rect 287666 375808 287671 375864
rect 284924 375806 287671 375808
rect 287605 375803 287671 375806
rect 232957 375458 233023 375461
rect 232957 375456 235060 375458
rect 232957 375400 232962 375456
rect 233018 375400 235060 375456
rect 232957 375398 235060 375400
rect 232957 375395 233023 375398
rect 288341 374234 288407 374237
rect 284924 374232 288407 374234
rect 284924 374176 288346 374232
rect 288402 374176 288407 374232
rect 284924 374174 288407 374176
rect 288341 374171 288407 374174
rect 232589 373554 232655 373557
rect 232589 373552 235060 373554
rect 232589 373496 232594 373552
rect 232650 373496 235060 373552
rect 232589 373494 235060 373496
rect 232589 373491 232655 373494
rect 287789 372602 287855 372605
rect 284924 372600 287855 372602
rect 284924 372544 287794 372600
rect 287850 372544 287855 372600
rect 284924 372542 287855 372544
rect 287789 372539 287855 372542
rect 234337 371650 234403 371653
rect 234337 371648 235060 371650
rect 234337 371592 234342 371648
rect 234398 371592 235060 371648
rect 234337 371590 235060 371592
rect 234337 371587 234403 371590
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 287605 370970 287671 370973
rect 284924 370968 287671 370970
rect 284924 370912 287610 370968
rect 287666 370912 287671 370968
rect 284924 370910 287671 370912
rect 287605 370907 287671 370910
rect 234153 369746 234219 369749
rect 234153 369744 235060 369746
rect 234153 369688 234158 369744
rect 234214 369688 235060 369744
rect 234153 369686 235060 369688
rect 234153 369683 234219 369686
rect 288341 369338 288407 369341
rect 284924 369336 288407 369338
rect 284924 369280 288346 369336
rect 288402 369280 288407 369336
rect 284924 369278 288407 369280
rect 288341 369275 288407 369278
rect 234245 367842 234311 367845
rect 234245 367840 235060 367842
rect 234245 367784 234250 367840
rect 234306 367784 235060 367840
rect 234245 367782 235060 367784
rect 234245 367779 234311 367782
rect 287973 367706 288039 367709
rect 284924 367704 288039 367706
rect 284924 367648 287978 367704
rect 288034 367648 288039 367704
rect 284924 367646 288039 367648
rect 287973 367643 288039 367646
rect 287605 366074 287671 366077
rect 284924 366072 287671 366074
rect 284924 366016 287610 366072
rect 287666 366016 287671 366072
rect 284924 366014 287671 366016
rect 287605 366011 287671 366014
rect 234061 365938 234127 365941
rect 234061 365936 235060 365938
rect 234061 365880 234066 365936
rect 234122 365880 235060 365936
rect 234061 365878 235060 365880
rect 234061 365875 234127 365878
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 288341 364442 288407 364445
rect 284924 364440 288407 364442
rect 284924 364384 288346 364440
rect 288402 364384 288407 364440
rect 284924 364382 288407 364384
rect 288341 364379 288407 364382
rect 232497 364034 232563 364037
rect 232497 364032 235060 364034
rect 232497 363976 232502 364032
rect 232558 363976 235060 364032
rect 232497 363974 235060 363976
rect 232497 363971 232563 363974
rect 287605 362946 287671 362949
rect 284924 362944 287671 362946
rect 284924 362888 287610 362944
rect 287666 362888 287671 362944
rect 284924 362886 287671 362888
rect 287605 362883 287671 362886
rect 233969 361994 234035 361997
rect 233969 361992 235060 361994
rect 233969 361936 233974 361992
rect 234030 361936 235060 361992
rect 233969 361934 235060 361936
rect 233969 361931 234035 361934
rect 287605 361314 287671 361317
rect 284924 361312 287671 361314
rect 284924 361256 287610 361312
rect 287666 361256 287671 361312
rect 284924 361254 287671 361256
rect 287605 361251 287671 361254
rect 233877 360090 233943 360093
rect 233877 360088 235060 360090
rect 233877 360032 233882 360088
rect 233938 360032 235060 360088
rect 233877 360030 235060 360032
rect 233877 360027 233943 360030
rect 287605 359682 287671 359685
rect 284924 359680 287671 359682
rect 284924 359624 287610 359680
rect 287666 359624 287671 359680
rect 284924 359622 287671 359624
rect 287605 359619 287671 359622
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 232313 358186 232379 358189
rect 232313 358184 235060 358186
rect 232313 358128 232318 358184
rect 232374 358128 235060 358184
rect 232313 358126 235060 358128
rect 232313 358123 232379 358126
rect 288341 358050 288407 358053
rect 284924 358048 288407 358050
rect 284924 357992 288346 358048
rect 288402 357992 288407 358048
rect 284924 357990 288407 357992
rect 288341 357987 288407 357990
rect 287789 356418 287855 356421
rect 284924 356416 287855 356418
rect 284924 356360 287794 356416
rect 287850 356360 287855 356416
rect 284924 356358 287855 356360
rect 287789 356355 287855 356358
rect 232405 356282 232471 356285
rect 232405 356280 235060 356282
rect 232405 356224 232410 356280
rect 232466 356224 235060 356280
rect 232405 356222 235060 356224
rect 232405 356219 232471 356222
rect 288341 354786 288407 354789
rect 284924 354784 288407 354786
rect 284924 354728 288346 354784
rect 288402 354728 288407 354784
rect 284924 354726 288407 354728
rect 288341 354723 288407 354726
rect 233785 354378 233851 354381
rect 233785 354376 235060 354378
rect 233785 354320 233790 354376
rect 233846 354320 235060 354376
rect 233785 354318 235060 354320
rect 233785 354315 233851 354318
rect 287513 353154 287579 353157
rect 284924 353152 287579 353154
rect 284924 353096 287518 353152
rect 287574 353096 287579 353152
rect 284924 353094 287579 353096
rect 287513 353091 287579 353094
rect 232221 352474 232287 352477
rect 232221 352472 235060 352474
rect 232221 352416 232226 352472
rect 232282 352416 235060 352472
rect 232221 352414 235060 352416
rect 232221 352411 232287 352414
rect 580717 351930 580783 351933
rect 583520 351930 584960 352020
rect 580717 351928 584960 351930
rect 580717 351872 580722 351928
rect 580778 351872 584960 351928
rect 580717 351870 584960 351872
rect 580717 351867 580783 351870
rect 583520 351780 584960 351870
rect 287237 351522 287303 351525
rect 284924 351520 287303 351522
rect 284924 351464 287242 351520
rect 287298 351464 287303 351520
rect 284924 351462 287303 351464
rect 287237 351459 287303 351462
rect 233693 350434 233759 350437
rect 233693 350432 235060 350434
rect 233693 350376 233698 350432
rect 233754 350376 235060 350432
rect 233693 350374 235060 350376
rect 233693 350371 233759 350374
rect 288341 350026 288407 350029
rect 284924 350024 288407 350026
rect 284924 349968 288346 350024
rect 288402 349968 288407 350024
rect 284924 349966 288407 349968
rect 288341 349963 288407 349966
rect 234521 348530 234587 348533
rect 234521 348528 235060 348530
rect 234521 348472 234526 348528
rect 234582 348472 235060 348528
rect 234521 348470 235060 348472
rect 234521 348467 234587 348470
rect 287973 348394 288039 348397
rect 284924 348392 288039 348394
rect 284924 348336 287978 348392
rect 288034 348336 288039 348392
rect 284924 348334 288039 348336
rect 287973 348331 288039 348334
rect 287973 346762 288039 346765
rect 284924 346760 288039 346762
rect 284924 346704 287978 346760
rect 288034 346704 288039 346760
rect 284924 346702 288039 346704
rect 287973 346699 288039 346702
rect 232865 346626 232931 346629
rect 232865 346624 235060 346626
rect 232865 346568 232870 346624
rect 232926 346568 235060 346624
rect 232865 346566 235060 346568
rect 232865 346563 232931 346566
rect -960 345402 480 345492
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 288341 345130 288407 345133
rect 284924 345128 288407 345130
rect 284924 345072 288346 345128
rect 288402 345072 288407 345128
rect 284924 345070 288407 345072
rect 288341 345067 288407 345070
rect 233509 344722 233575 344725
rect 233509 344720 235060 344722
rect 233509 344664 233514 344720
rect 233570 344664 235060 344720
rect 233509 344662 235060 344664
rect 233509 344659 233575 344662
rect 288341 343498 288407 343501
rect 284924 343496 288407 343498
rect 284924 343440 288346 343496
rect 288402 343440 288407 343496
rect 284924 343438 288407 343440
rect 288341 343435 288407 343438
rect 232037 342818 232103 342821
rect 232037 342816 235060 342818
rect 232037 342760 232042 342816
rect 232098 342760 235060 342816
rect 232037 342758 235060 342760
rect 232037 342755 232103 342758
rect 288341 341866 288407 341869
rect 284924 341864 288407 341866
rect 284924 341808 288346 341864
rect 288402 341808 288407 341864
rect 284924 341806 288407 341808
rect 288341 341803 288407 341806
rect 233601 340914 233667 340917
rect 233601 340912 235060 340914
rect 233601 340856 233606 340912
rect 233662 340856 235060 340912
rect 233601 340854 235060 340856
rect 233601 340851 233667 340854
rect 287789 340234 287855 340237
rect 284924 340232 287855 340234
rect 284924 340176 287794 340232
rect 287850 340176 287855 340232
rect 284924 340174 287855 340176
rect 287789 340171 287855 340174
rect 234705 339010 234771 339013
rect 234705 339008 235060 339010
rect 234705 338952 234710 339008
rect 234766 338952 235060 339008
rect 234705 338950 235060 338952
rect 234705 338947 234771 338950
rect 287421 338738 287487 338741
rect 284924 338736 287487 338738
rect 284924 338680 287426 338736
rect 287482 338680 287487 338736
rect 284924 338678 287487 338680
rect 287421 338675 287487 338678
rect 583520 338452 584960 338692
rect 287605 338194 287671 338197
rect 279006 338192 287671 338194
rect 279006 338136 287610 338192
rect 287666 338136 287671 338192
rect 279006 338134 287671 338136
rect 233233 338058 233299 338061
rect 233233 338056 241208 338058
rect 233233 338000 233238 338056
rect 233294 338000 241208 338056
rect 233233 337998 241208 338000
rect 233233 337995 233299 337998
rect 241148 337925 241208 337998
rect 243862 337998 246314 338058
rect 233325 337922 233391 337925
rect 236407 337922 236473 337925
rect 238523 337924 238589 337925
rect 238518 337922 238524 337924
rect 233325 337920 236473 337922
rect 233325 337864 233330 337920
rect 233386 337864 236412 337920
rect 236468 337864 236473 337920
rect 233325 337862 236473 337864
rect 238432 337862 238524 337922
rect 233325 337859 233391 337862
rect 236407 337859 236473 337862
rect 238518 337860 238524 337862
rect 238588 337860 238594 337924
rect 239254 337860 239260 337924
rect 239324 337922 239330 337924
rect 239443 337922 239509 337925
rect 239324 337920 239509 337922
rect 239324 337864 239448 337920
rect 239504 337864 239509 337920
rect 239324 337862 239509 337864
rect 239324 337860 239330 337862
rect 238523 337859 238589 337860
rect 239443 337859 239509 337862
rect 239627 337920 239693 337925
rect 239627 337864 239632 337920
rect 239688 337864 239693 337920
rect 239627 337859 239693 337864
rect 239811 337920 239877 337925
rect 239811 337864 239816 337920
rect 239872 337864 239877 337920
rect 239811 337859 239877 337864
rect 241148 337920 241257 337925
rect 241148 337864 241196 337920
rect 241252 337864 241257 337920
rect 242203 337920 242269 337925
rect 241148 337862 241257 337864
rect 241191 337859 241257 337862
rect 242019 337886 242085 337891
rect 235533 337786 235599 337789
rect 239630 337786 239690 337859
rect 235533 337784 239690 337786
rect 235533 337728 235538 337784
rect 235594 337728 239690 337784
rect 235533 337726 239690 337728
rect 239814 337789 239874 337859
rect 242019 337830 242024 337886
rect 242080 337830 242085 337886
rect 242203 337864 242208 337920
rect 242264 337864 242269 337920
rect 242203 337859 242269 337864
rect 242939 337920 243005 337925
rect 242939 337864 242944 337920
rect 243000 337864 243005 337920
rect 242939 337859 243005 337864
rect 242019 337825 242085 337830
rect 239814 337784 239923 337789
rect 239814 337728 239862 337784
rect 239918 337728 239923 337784
rect 239814 337726 239923 337728
rect 235533 337723 235599 337726
rect 239857 337723 239923 337726
rect 238518 337588 238524 337652
rect 238588 337650 238594 337652
rect 239489 337650 239555 337653
rect 238588 337648 239555 337650
rect 238588 337592 239494 337648
rect 239550 337592 239555 337648
rect 238588 337590 239555 337592
rect 238588 337588 238594 337590
rect 239489 337587 239555 337590
rect 240961 337650 241027 337653
rect 241145 337650 241211 337653
rect 240961 337648 241211 337650
rect 240961 337592 240966 337648
rect 241022 337592 241150 337648
rect 241206 337592 241211 337648
rect 240961 337590 241211 337592
rect 240961 337587 241027 337590
rect 241145 337587 241211 337590
rect 241881 337514 241947 337517
rect 242022 337514 242082 337825
rect 242206 337789 242266 337859
rect 242942 337789 243002 337859
rect 242206 337784 242315 337789
rect 242206 337728 242254 337784
rect 242310 337728 242315 337784
rect 242206 337726 242315 337728
rect 242249 337723 242315 337726
rect 242893 337784 243002 337789
rect 242893 337728 242898 337784
rect 242954 337728 243002 337784
rect 242893 337726 243002 337728
rect 243169 337786 243235 337789
rect 243862 337786 243922 337998
rect 246254 337925 246314 337998
rect 279006 337959 279066 338134
rect 287605 338131 287671 338134
rect 249931 337954 249997 337959
rect 244871 337922 244937 337925
rect 245699 337924 245765 337925
rect 245694 337922 245700 337924
rect 244414 337920 244937 337922
rect 244043 337886 244109 337891
rect 244043 337830 244048 337886
rect 244104 337830 244109 337886
rect 244043 337825 244109 337830
rect 244414 337864 244876 337920
rect 244932 337864 244937 337920
rect 244414 337862 244937 337864
rect 245608 337862 245700 337922
rect 243169 337784 243922 337786
rect 243169 337728 243174 337784
rect 243230 337728 243922 337784
rect 243169 337726 243922 337728
rect 242893 337723 242959 337726
rect 243169 337723 243235 337726
rect 244046 337653 244106 337825
rect 244046 337648 244155 337653
rect 244046 337592 244094 337648
rect 244150 337592 244155 337648
rect 244046 337590 244155 337592
rect 244089 337587 244155 337590
rect 241881 337512 242082 337514
rect 241881 337456 241886 337512
rect 241942 337456 242082 337512
rect 241881 337454 242082 337456
rect 243721 337514 243787 337517
rect 244414 337514 244474 337862
rect 244871 337859 244937 337862
rect 245694 337860 245700 337862
rect 245764 337860 245770 337924
rect 246067 337920 246133 337925
rect 246067 337864 246072 337920
rect 246128 337864 246133 337920
rect 245699 337859 245765 337860
rect 246067 337859 246133 337864
rect 246251 337920 246317 337925
rect 246251 337864 246256 337920
rect 246312 337864 246317 337920
rect 247723 337920 247789 337925
rect 246251 337859 246317 337864
rect 247355 337886 247421 337891
rect 244549 337786 244615 337789
rect 246070 337786 246130 337859
rect 247355 337830 247360 337886
rect 247416 337830 247421 337886
rect 247723 337864 247728 337920
rect 247784 337864 247789 337920
rect 249379 337920 249445 337925
rect 247723 337859 247789 337864
rect 247907 337886 247973 337891
rect 247355 337825 247421 337830
rect 244549 337784 246130 337786
rect 244549 337728 244554 337784
rect 244610 337728 246130 337784
rect 244549 337726 246130 337728
rect 246987 337784 247053 337789
rect 246987 337728 246992 337784
rect 247048 337728 247053 337784
rect 244549 337723 244615 337726
rect 246987 337723 247053 337728
rect 245653 337652 245719 337653
rect 245653 337648 245700 337652
rect 245764 337650 245770 337652
rect 245929 337650 245995 337653
rect 246990 337650 247050 337723
rect 245653 337592 245658 337648
rect 245653 337588 245700 337592
rect 245764 337590 245810 337650
rect 245929 337648 247050 337650
rect 245929 337592 245934 337648
rect 245990 337592 247050 337648
rect 245929 337590 247050 337592
rect 245764 337588 245770 337590
rect 245653 337587 245719 337588
rect 245929 337587 245995 337590
rect 243721 337512 244474 337514
rect 243721 337456 243726 337512
rect 243782 337456 244474 337512
rect 243721 337454 244474 337456
rect 247358 337517 247418 337825
rect 247358 337512 247467 337517
rect 247358 337456 247406 337512
rect 247462 337456 247467 337512
rect 247358 337454 247467 337456
rect 241881 337451 241947 337454
rect 243721 337451 243787 337454
rect 247401 337451 247467 337454
rect 247585 337514 247651 337517
rect 247726 337514 247786 337859
rect 247907 337830 247912 337886
rect 247968 337830 247973 337886
rect 249379 337864 249384 337920
rect 249440 337864 249445 337920
rect 249931 337898 249936 337954
rect 249992 337898 249997 337954
rect 249931 337893 249997 337898
rect 251035 337954 251101 337959
rect 251035 337898 251040 337954
rect 251096 337898 251101 337954
rect 251035 337893 251101 337898
rect 252875 337954 252941 337959
rect 252875 337898 252880 337954
rect 252936 337898 252941 337954
rect 252875 337893 252941 337898
rect 254899 337954 254965 337959
rect 254899 337898 254904 337954
rect 254960 337898 254965 337954
rect 254899 337893 254965 337898
rect 255267 337954 255333 337959
rect 255267 337898 255272 337954
rect 255328 337898 255333 337954
rect 255267 337893 255333 337898
rect 255451 337954 255517 337959
rect 255451 337898 255456 337954
rect 255512 337898 255517 337954
rect 255451 337893 255517 337898
rect 255819 337954 255885 337959
rect 255819 337898 255824 337954
rect 255880 337898 255885 337954
rect 255819 337893 255885 337898
rect 256923 337954 256989 337959
rect 256923 337898 256928 337954
rect 256984 337898 256989 337954
rect 256923 337893 256989 337898
rect 257659 337954 257725 337959
rect 257659 337898 257664 337954
rect 257720 337898 257725 337954
rect 257659 337893 257725 337898
rect 258211 337954 258277 337959
rect 258211 337898 258216 337954
rect 258272 337898 258277 337954
rect 258211 337893 258277 337898
rect 258395 337954 258461 337959
rect 258395 337898 258400 337954
rect 258456 337898 258461 337954
rect 258395 337893 258461 337898
rect 258579 337954 258645 337959
rect 258579 337898 258584 337954
rect 258640 337898 258645 337954
rect 258579 337893 258645 337898
rect 258947 337954 259013 337959
rect 258947 337898 258952 337954
rect 259008 337898 259013 337954
rect 258947 337893 259013 337898
rect 259131 337954 259197 337959
rect 259131 337898 259136 337954
rect 259192 337898 259197 337954
rect 259131 337893 259197 337898
rect 259315 337954 259381 337959
rect 259315 337898 259320 337954
rect 259376 337898 259381 337954
rect 259315 337893 259381 337898
rect 259499 337954 259565 337959
rect 259499 337898 259504 337954
rect 259560 337898 259565 337954
rect 264283 337954 264349 337959
rect 259499 337893 259565 337898
rect 263547 337920 263613 337925
rect 249379 337859 249445 337864
rect 247907 337825 247973 337830
rect 247910 337653 247970 337825
rect 249382 337789 249442 337859
rect 249934 337789 249994 337893
rect 249382 337784 249491 337789
rect 249382 337728 249430 337784
rect 249486 337728 249491 337784
rect 249382 337726 249491 337728
rect 249425 337723 249491 337726
rect 249885 337784 249994 337789
rect 249885 337728 249890 337784
rect 249946 337728 249994 337784
rect 249885 337726 249994 337728
rect 251038 337789 251098 337893
rect 251038 337784 251147 337789
rect 251038 337728 251086 337784
rect 251142 337728 251147 337784
rect 251038 337726 251147 337728
rect 249885 337723 249951 337726
rect 251081 337723 251147 337726
rect 252878 337653 252938 337893
rect 254902 337789 254962 337893
rect 254531 337784 254597 337789
rect 254531 337728 254536 337784
rect 254592 337728 254597 337784
rect 254531 337723 254597 337728
rect 254853 337784 254962 337789
rect 254853 337728 254858 337784
rect 254914 337728 254962 337784
rect 254853 337726 254962 337728
rect 255270 337789 255330 337893
rect 255454 337789 255514 337893
rect 255822 337789 255882 337893
rect 256926 337789 256986 337893
rect 257662 337789 257722 337893
rect 255270 337784 255379 337789
rect 255270 337728 255318 337784
rect 255374 337728 255379 337784
rect 255270 337726 255379 337728
rect 255454 337784 255563 337789
rect 255454 337728 255502 337784
rect 255558 337728 255563 337784
rect 255454 337726 255563 337728
rect 255822 337784 255931 337789
rect 255822 337728 255870 337784
rect 255926 337728 255931 337784
rect 255822 337726 255931 337728
rect 256926 337784 257035 337789
rect 256926 337728 256974 337784
rect 257030 337728 257035 337784
rect 256926 337726 257035 337728
rect 254853 337723 254919 337726
rect 255313 337723 255379 337726
rect 255497 337723 255563 337726
rect 255865 337723 255931 337726
rect 256969 337723 257035 337726
rect 257659 337784 257725 337789
rect 257659 337728 257664 337784
rect 257720 337728 257725 337784
rect 257659 337723 257725 337728
rect 254534 337653 254594 337723
rect 247910 337648 248019 337653
rect 247910 337592 247958 337648
rect 248014 337592 248019 337648
rect 247910 337590 248019 337592
rect 252878 337648 252987 337653
rect 252878 337592 252926 337648
rect 252982 337592 252987 337648
rect 252878 337590 252987 337592
rect 247953 337587 248019 337590
rect 252921 337587 252987 337590
rect 254485 337648 254594 337653
rect 254485 337592 254490 337648
rect 254546 337592 254594 337648
rect 254485 337590 254594 337592
rect 254485 337587 254551 337590
rect 247585 337512 247786 337514
rect 247585 337456 247590 337512
rect 247646 337456 247786 337512
rect 247585 337454 247786 337456
rect 247585 337451 247651 337454
rect 258214 337378 258274 337893
rect 258398 337789 258458 337893
rect 258398 337784 258507 337789
rect 258398 337728 258446 337784
rect 258502 337728 258507 337784
rect 258398 337726 258507 337728
rect 258582 337786 258642 337893
rect 258809 337786 258875 337789
rect 258582 337784 258875 337786
rect 258582 337728 258814 337784
rect 258870 337728 258875 337784
rect 258582 337726 258875 337728
rect 258441 337723 258507 337726
rect 258809 337723 258875 337726
rect 258950 337653 259010 337893
rect 258950 337648 259059 337653
rect 258950 337592 258998 337648
rect 259054 337592 259059 337648
rect 258950 337590 259059 337592
rect 258993 337587 259059 337590
rect 259134 337517 259194 337893
rect 259318 337789 259378 337893
rect 259502 337789 259562 337893
rect 263547 337864 263552 337920
rect 263608 337864 263613 337920
rect 264283 337898 264288 337954
rect 264344 337898 264349 337954
rect 264283 337893 264349 337898
rect 264651 337954 264717 337959
rect 264651 337898 264656 337954
rect 264712 337898 264717 337954
rect 264651 337893 264717 337898
rect 264835 337954 264901 337959
rect 264835 337898 264840 337954
rect 264896 337922 264901 337954
rect 268699 337956 268765 337959
rect 268699 337954 268822 337956
rect 268699 337924 268704 337954
rect 268760 337924 268822 337954
rect 272931 337954 272997 337959
rect 264896 337898 264990 337922
rect 264835 337893 264990 337898
rect 263547 337859 263613 337864
rect 259318 337784 259427 337789
rect 259318 337728 259366 337784
rect 259422 337728 259427 337784
rect 259318 337726 259427 337728
rect 259502 337784 259611 337789
rect 259502 337728 259550 337784
rect 259606 337728 259611 337784
rect 259502 337726 259611 337728
rect 263550 337786 263610 337859
rect 263685 337786 263751 337789
rect 263550 337784 263751 337786
rect 263550 337728 263690 337784
rect 263746 337728 263751 337784
rect 263550 337726 263751 337728
rect 259361 337723 259427 337726
rect 259545 337723 259611 337726
rect 263685 337723 263751 337726
rect 259085 337512 259194 337517
rect 259085 337456 259090 337512
rect 259146 337456 259194 337512
rect 259085 337454 259194 337456
rect 264286 337514 264346 337893
rect 264654 337786 264714 337893
rect 264838 337862 264990 337893
rect 264930 337789 264990 337862
rect 266123 337886 266189 337891
rect 266123 337830 266128 337886
rect 266184 337830 266189 337886
rect 268694 337860 268700 337924
rect 268764 337896 268822 337924
rect 268883 337920 268949 337925
rect 268764 337860 268770 337896
rect 268883 337864 268888 337920
rect 268944 337864 268949 337920
rect 268883 337859 268949 337864
rect 269251 337920 269317 337925
rect 269251 337864 269256 337920
rect 269312 337864 269317 337920
rect 269251 337859 269317 337864
rect 269619 337920 269685 337925
rect 269619 337864 269624 337920
rect 269680 337864 269685 337920
rect 269619 337859 269685 337864
rect 270355 337920 270421 337925
rect 270355 337864 270360 337920
rect 270416 337864 270421 337920
rect 270355 337859 270421 337864
rect 270723 337920 270789 337925
rect 270723 337864 270728 337920
rect 270784 337864 270789 337920
rect 270723 337859 270789 337864
rect 271183 337922 271249 337925
rect 272103 337922 272169 337925
rect 272558 337922 272564 337924
rect 271183 337920 271522 337922
rect 271183 337864 271188 337920
rect 271244 337864 271522 337920
rect 271183 337862 271522 337864
rect 271183 337859 271249 337862
rect 266123 337825 266189 337830
rect 264789 337786 264855 337789
rect 264654 337784 264855 337786
rect 264654 337728 264794 337784
rect 264850 337728 264855 337784
rect 264654 337726 264855 337728
rect 264930 337784 265039 337789
rect 264930 337728 264978 337784
rect 265034 337728 265039 337784
rect 264930 337726 265039 337728
rect 264789 337723 264855 337726
rect 264973 337723 265039 337726
rect 266126 337653 266186 337825
rect 268886 337786 268946 337859
rect 269021 337786 269087 337789
rect 268886 337784 269087 337786
rect 268886 337728 269026 337784
rect 269082 337728 269087 337784
rect 268886 337726 269087 337728
rect 269021 337723 269087 337726
rect 266077 337648 266186 337653
rect 266077 337592 266082 337648
rect 266138 337592 266186 337648
rect 266077 337590 266186 337592
rect 266077 337587 266143 337590
rect 268561 337514 268627 337517
rect 264286 337512 268627 337514
rect 264286 337456 268566 337512
rect 268622 337456 268627 337512
rect 264286 337454 268627 337456
rect 269254 337514 269314 337859
rect 269622 337653 269682 337859
rect 270358 337789 270418 337859
rect 270358 337784 270467 337789
rect 270358 337728 270406 337784
rect 270462 337728 270467 337784
rect 270358 337726 270467 337728
rect 270401 337723 270467 337726
rect 269622 337648 269731 337653
rect 269622 337592 269670 337648
rect 269726 337592 269731 337648
rect 269622 337590 269731 337592
rect 269665 337587 269731 337590
rect 270726 337517 270786 337859
rect 271462 337789 271522 337862
rect 272103 337920 272564 337922
rect 272103 337864 272108 337920
rect 272164 337864 272564 337920
rect 272103 337862 272564 337864
rect 272103 337859 272169 337862
rect 272558 337860 272564 337862
rect 272628 337860 272634 337924
rect 272931 337898 272936 337954
rect 272992 337898 272997 337954
rect 274955 337954 275021 337959
rect 272931 337893 272997 337898
rect 274495 337920 274561 337925
rect 272934 337789 272994 337893
rect 273115 337886 273181 337891
rect 273115 337830 273120 337886
rect 273176 337830 273181 337886
rect 274495 337864 274500 337920
rect 274556 337864 274561 337920
rect 274955 337898 274960 337954
rect 275016 337898 275021 337954
rect 274955 337893 275021 337898
rect 275875 337954 275941 337959
rect 275875 337898 275880 337954
rect 275936 337898 275941 337954
rect 275875 337893 275941 337898
rect 276059 337954 276125 337959
rect 276059 337898 276064 337954
rect 276120 337898 276125 337954
rect 276059 337893 276125 337898
rect 276243 337954 276309 337959
rect 276243 337898 276248 337954
rect 276304 337898 276309 337954
rect 276243 337893 276309 337898
rect 276703 337956 276769 337959
rect 276703 337954 276812 337956
rect 276703 337898 276708 337954
rect 276764 337898 276812 337954
rect 276703 337893 276812 337898
rect 276979 337954 277045 337959
rect 276979 337898 276984 337954
rect 277040 337898 277045 337954
rect 278451 337954 278517 337959
rect 276979 337893 277045 337898
rect 277899 337920 277965 337925
rect 278267 337924 278333 337925
rect 278262 337922 278268 337924
rect 274495 337859 274561 337864
rect 273115 337825 273181 337830
rect 271462 337784 271571 337789
rect 271462 337728 271510 337784
rect 271566 337728 271571 337784
rect 271462 337726 271571 337728
rect 271505 337723 271571 337726
rect 272885 337784 272994 337789
rect 272885 337728 272890 337784
rect 272946 337728 272994 337784
rect 272885 337726 272994 337728
rect 272885 337723 272951 337726
rect 273118 337653 273178 337825
rect 273069 337648 273178 337653
rect 273069 337592 273074 337648
rect 273130 337592 273178 337648
rect 273069 337590 273178 337592
rect 273069 337587 273135 337590
rect 270125 337514 270191 337517
rect 269254 337512 270191 337514
rect 269254 337456 270130 337512
rect 270186 337456 270191 337512
rect 269254 337454 270191 337456
rect 270726 337512 270835 337517
rect 270726 337456 270774 337512
rect 270830 337456 270835 337512
rect 270726 337454 270835 337456
rect 274498 337514 274558 337859
rect 274633 337514 274699 337517
rect 274498 337512 274699 337514
rect 274498 337456 274638 337512
rect 274694 337456 274699 337512
rect 274498 337454 274699 337456
rect 274958 337514 275018 337893
rect 275878 337789 275938 337893
rect 275878 337784 275987 337789
rect 275878 337728 275926 337784
rect 275982 337728 275987 337784
rect 275878 337726 275987 337728
rect 275921 337723 275987 337726
rect 276062 337650 276122 337893
rect 276246 337789 276306 337893
rect 276197 337784 276306 337789
rect 276197 337728 276202 337784
rect 276258 337728 276306 337784
rect 276197 337726 276306 337728
rect 276197 337723 276263 337726
rect 276289 337650 276355 337653
rect 276062 337648 276355 337650
rect 276062 337592 276294 337648
rect 276350 337592 276355 337648
rect 276062 337590 276355 337592
rect 276289 337587 276355 337590
rect 275829 337514 275895 337517
rect 274958 337512 275895 337514
rect 274958 337456 275834 337512
rect 275890 337456 275895 337512
rect 274958 337454 275895 337456
rect 259085 337451 259151 337454
rect 268561 337451 268627 337454
rect 270125 337451 270191 337454
rect 270769 337451 270835 337454
rect 274633 337451 274699 337454
rect 275829 337451 275895 337454
rect 259177 337378 259243 337381
rect 258214 337376 259243 337378
rect 258214 337320 259182 337376
rect 259238 337320 259243 337376
rect 258214 337318 259243 337320
rect 276752 337378 276812 337893
rect 276982 337786 277042 337893
rect 277899 337864 277904 337920
rect 277960 337864 277965 337920
rect 277899 337859 277965 337864
rect 278176 337862 278268 337922
rect 278262 337860 278268 337862
rect 278332 337860 278338 337924
rect 278451 337898 278456 337954
rect 278512 337898 278517 337954
rect 278451 337893 278517 337898
rect 278819 337954 278885 337959
rect 278819 337898 278824 337954
rect 278880 337898 278885 337954
rect 278819 337893 278885 337898
rect 279003 337954 279069 337959
rect 279003 337898 279008 337954
rect 279064 337898 279069 337954
rect 280383 337954 280449 337959
rect 279831 337922 279897 337925
rect 279003 337893 279069 337898
rect 279558 337920 279897 337922
rect 278267 337859 278333 337860
rect 277902 337789 277962 337859
rect 277117 337786 277183 337789
rect 276982 337784 277183 337786
rect 276982 337728 277122 337784
rect 277178 337728 277183 337784
rect 276982 337726 277183 337728
rect 277902 337784 278011 337789
rect 277902 337728 277950 337784
rect 278006 337728 278011 337784
rect 277902 337726 278011 337728
rect 277117 337723 277183 337726
rect 277945 337723 278011 337726
rect 277853 337650 277919 337653
rect 278454 337650 278514 337893
rect 277853 337648 278514 337650
rect 277853 337592 277858 337648
rect 277914 337592 278514 337648
rect 277853 337590 278514 337592
rect 278822 337650 278882 337893
rect 279558 337864 279836 337920
rect 279892 337864 279897 337920
rect 280383 337898 280388 337954
rect 280444 337898 280449 337954
rect 282591 337956 282657 337959
rect 282591 337954 282700 337956
rect 280383 337893 280449 337898
rect 282315 337920 282381 337925
rect 282591 337922 282596 337954
rect 279558 337862 279897 337864
rect 278957 337650 279023 337653
rect 278822 337648 279023 337650
rect 278822 337592 278962 337648
rect 279018 337592 279023 337648
rect 278822 337590 279023 337592
rect 277853 337587 277919 337590
rect 278957 337587 279023 337590
rect 279417 337650 279483 337653
rect 279558 337650 279618 337862
rect 279831 337859 279897 337862
rect 280386 337786 280446 337893
rect 280659 337886 280725 337891
rect 280659 337830 280664 337886
rect 280720 337830 280725 337886
rect 280659 337825 280725 337830
rect 281395 337886 281461 337891
rect 281395 337830 281400 337886
rect 281456 337830 281461 337886
rect 282315 337864 282320 337920
rect 282376 337864 282381 337920
rect 282315 337859 282381 337864
rect 282502 337898 282596 337922
rect 282652 337898 282700 337954
rect 282502 337862 282700 337898
rect 283235 337954 283301 337959
rect 283235 337898 283240 337954
rect 283296 337898 283301 337954
rect 284155 337954 284221 337959
rect 283235 337893 283301 337898
rect 283419 337920 283485 337925
rect 281395 337825 281461 337830
rect 279417 337648 279618 337650
rect 279417 337592 279422 337648
rect 279478 337592 279618 337648
rect 279417 337590 279618 337592
rect 280294 337726 280446 337786
rect 279417 337587 279483 337590
rect 277117 337378 277183 337381
rect 276752 337376 277183 337378
rect 276752 337320 277122 337376
rect 277178 337320 277183 337376
rect 276752 337318 277183 337320
rect 280294 337378 280354 337726
rect 280429 337650 280495 337653
rect 280662 337650 280722 337825
rect 280429 337648 280722 337650
rect 280429 337592 280434 337648
rect 280490 337592 280722 337648
rect 280429 337590 280722 337592
rect 281257 337650 281323 337653
rect 281398 337650 281458 337825
rect 281257 337648 281458 337650
rect 281257 337592 281262 337648
rect 281318 337592 281458 337648
rect 281257 337590 281458 337592
rect 280429 337587 280495 337590
rect 281257 337587 281323 337590
rect 282318 337517 282378 337859
rect 282502 337789 282562 337862
rect 282502 337784 282611 337789
rect 282502 337728 282550 337784
rect 282606 337728 282611 337784
rect 282502 337726 282611 337728
rect 282545 337723 282611 337726
rect 282269 337512 282378 337517
rect 282269 337456 282274 337512
rect 282330 337456 282378 337512
rect 282269 337454 282378 337456
rect 283238 337514 283298 337893
rect 283419 337864 283424 337920
rect 283480 337864 283485 337920
rect 284155 337898 284160 337954
rect 284216 337898 284221 337954
rect 284155 337893 284221 337898
rect 284615 337922 284681 337925
rect 285489 337922 285555 337925
rect 284615 337920 285555 337922
rect 283419 337859 283485 337864
rect 283971 337886 284037 337891
rect 283422 337653 283482 337859
rect 283971 337830 283976 337886
rect 284032 337830 284037 337886
rect 283971 337825 284037 337830
rect 283974 337653 284034 337825
rect 284158 337789 284218 337893
rect 284615 337864 284620 337920
rect 284676 337864 285494 337920
rect 285550 337864 285555 337920
rect 284615 337862 285555 337864
rect 284615 337859 284681 337862
rect 285489 337859 285555 337862
rect 284109 337784 284218 337789
rect 284109 337728 284114 337784
rect 284170 337728 284218 337784
rect 284109 337726 284218 337728
rect 284109 337723 284175 337726
rect 283373 337648 283482 337653
rect 283373 337592 283378 337648
rect 283434 337592 283482 337648
rect 283373 337590 283482 337592
rect 283925 337648 284034 337653
rect 283925 337592 283930 337648
rect 283986 337592 284034 337648
rect 283925 337590 284034 337592
rect 283373 337587 283439 337590
rect 283925 337587 283991 337590
rect 287329 337514 287395 337517
rect 283238 337512 287395 337514
rect 283238 337456 287334 337512
rect 287390 337456 287395 337512
rect 283238 337454 287395 337456
rect 282269 337451 282335 337454
rect 287329 337451 287395 337454
rect 286869 337378 286935 337381
rect 280294 337376 286935 337378
rect 280294 337320 286874 337376
rect 286930 337320 286935 337376
rect 280294 337318 286935 337320
rect 259177 337315 259243 337318
rect 277117 337315 277183 337318
rect 286869 337315 286935 337318
rect 50981 336698 51047 336701
rect 238753 336698 238819 336701
rect 50981 336696 238819 336698
rect 50981 336640 50986 336696
rect 51042 336640 238758 336696
rect 238814 336640 238819 336696
rect 50981 336638 238819 336640
rect 50981 336635 51047 336638
rect 238753 336635 238819 336638
rect 282361 336698 282427 336701
rect 304257 336698 304323 336701
rect 282361 336696 304323 336698
rect 282361 336640 282366 336696
rect 282422 336640 304262 336696
rect 304318 336640 304323 336696
rect 282361 336638 304323 336640
rect 282361 336635 282427 336638
rect 304257 336635 304323 336638
rect 38561 336562 38627 336565
rect 238017 336562 238083 336565
rect 38561 336560 238083 336562
rect 38561 336504 38566 336560
rect 38622 336504 238022 336560
rect 238078 336504 238083 336560
rect 38561 336502 238083 336504
rect 38561 336499 38627 336502
rect 238017 336499 238083 336502
rect 269021 336562 269087 336565
rect 282913 336562 282979 336565
rect 304441 336562 304507 336565
rect 269021 336560 278146 336562
rect 269021 336504 269026 336560
rect 269082 336504 278146 336560
rect 269021 336502 278146 336504
rect 269021 336499 269087 336502
rect 33041 336426 33107 336429
rect 237649 336426 237715 336429
rect 33041 336424 237715 336426
rect 33041 336368 33046 336424
rect 33102 336368 237654 336424
rect 237710 336368 237715 336424
rect 33041 336366 237715 336368
rect 33041 336363 33107 336366
rect 237649 336363 237715 336366
rect 273161 336426 273227 336429
rect 277485 336426 277551 336429
rect 273161 336424 277551 336426
rect 273161 336368 273166 336424
rect 273222 336368 277490 336424
rect 277546 336368 277551 336424
rect 273161 336366 277551 336368
rect 278086 336426 278146 336502
rect 282913 336560 304507 336562
rect 282913 336504 282918 336560
rect 282974 336504 304446 336560
rect 304502 336504 304507 336560
rect 282913 336502 304507 336504
rect 282913 336499 282979 336502
rect 304441 336499 304507 336502
rect 398097 336426 398163 336429
rect 278086 336424 398163 336426
rect 278086 336368 398102 336424
rect 398158 336368 398163 336424
rect 278086 336366 398163 336368
rect 273161 336363 273227 336366
rect 277485 336363 277551 336366
rect 398097 336363 398163 336366
rect 31661 336290 31727 336293
rect 234981 336290 235047 336293
rect 31661 336288 235047 336290
rect 31661 336232 31666 336288
rect 31722 336232 234986 336288
rect 235042 336232 235047 336288
rect 31661 336230 235047 336232
rect 31661 336227 31727 336230
rect 234981 336227 235047 336230
rect 269849 336290 269915 336293
rect 416037 336290 416103 336293
rect 269849 336288 416103 336290
rect 269849 336232 269854 336288
rect 269910 336232 416042 336288
rect 416098 336232 416103 336288
rect 269849 336230 416103 336232
rect 269849 336227 269915 336230
rect 416037 336227 416103 336230
rect 234613 336154 234679 336157
rect 242801 336154 242867 336157
rect 234613 336152 242867 336154
rect 234613 336096 234618 336152
rect 234674 336096 242806 336152
rect 242862 336096 242867 336152
rect 234613 336094 242867 336096
rect 234613 336091 234679 336094
rect 242801 336091 242867 336094
rect 270401 336154 270467 336157
rect 420177 336154 420243 336157
rect 270401 336152 420243 336154
rect 270401 336096 270406 336152
rect 270462 336096 420182 336152
rect 420238 336096 420243 336152
rect 270401 336094 420243 336096
rect 270401 336091 270467 336094
rect 420177 336091 420243 336094
rect 15101 336018 15167 336021
rect 236085 336018 236151 336021
rect 15101 336016 236151 336018
rect 15101 335960 15106 336016
rect 15162 335960 236090 336016
rect 236146 335960 236151 336016
rect 15101 335958 236151 335960
rect 15101 335955 15167 335958
rect 236085 335955 236151 335958
rect 236729 336018 236795 336021
rect 241237 336018 241303 336021
rect 236729 336016 241303 336018
rect 236729 335960 236734 336016
rect 236790 335960 241242 336016
rect 241298 335960 241303 336016
rect 236729 335958 241303 335960
rect 236729 335955 236795 335958
rect 241237 335955 241303 335958
rect 270585 336018 270651 336021
rect 422937 336018 423003 336021
rect 270585 336016 423003 336018
rect 270585 335960 270590 336016
rect 270646 335960 422942 336016
rect 422998 335960 423003 336016
rect 270585 335958 423003 335960
rect 270585 335955 270651 335958
rect 422937 335955 423003 335958
rect 57881 335882 57947 335885
rect 235533 335882 235599 335885
rect 57881 335880 235599 335882
rect 57881 335824 57886 335880
rect 57942 335824 235538 335880
rect 235594 335824 235599 335880
rect 57881 335822 235599 335824
rect 57881 335819 57947 335822
rect 235533 335819 235599 335822
rect 277485 335882 277551 335885
rect 286317 335882 286383 335885
rect 277485 335880 286383 335882
rect 277485 335824 277490 335880
rect 277546 335824 286322 335880
rect 286378 335824 286383 335880
rect 277485 335822 286383 335824
rect 277485 335819 277551 335822
rect 286317 335819 286383 335822
rect 236177 335746 236243 335749
rect 256141 335746 256207 335749
rect 236177 335744 256207 335746
rect 236177 335688 236182 335744
rect 236238 335688 256146 335744
rect 256202 335688 256207 335744
rect 236177 335686 256207 335688
rect 236177 335683 236243 335686
rect 256141 335683 256207 335686
rect 274817 335746 274883 335749
rect 280889 335746 280955 335749
rect 274817 335744 280955 335746
rect 274817 335688 274822 335744
rect 274878 335688 280894 335744
rect 280950 335688 280955 335744
rect 274817 335686 280955 335688
rect 274817 335683 274883 335686
rect 280889 335683 280955 335686
rect 15193 335610 15259 335613
rect 236361 335610 236427 335613
rect 254577 335610 254643 335613
rect 15193 335608 254643 335610
rect 15193 335552 15198 335608
rect 15254 335552 236366 335608
rect 236422 335552 254582 335608
rect 254638 335552 254643 335608
rect 15193 335550 254643 335552
rect 15193 335547 15259 335550
rect 236361 335547 236427 335550
rect 254577 335547 254643 335550
rect 272558 335548 272564 335612
rect 272628 335610 272634 335612
rect 284385 335610 284451 335613
rect 272628 335608 284451 335610
rect 272628 335552 284390 335608
rect 284446 335552 284451 335608
rect 272628 335550 284451 335552
rect 272628 335548 272634 335550
rect 284385 335547 284451 335550
rect 24853 335474 24919 335477
rect 236821 335474 236887 335477
rect 24853 335472 236887 335474
rect 24853 335416 24858 335472
rect 24914 335416 236826 335472
rect 236882 335416 236887 335472
rect 24853 335414 236887 335416
rect 24853 335411 24919 335414
rect 236821 335411 236887 335414
rect 237005 335474 237071 335477
rect 237373 335474 237439 335477
rect 237005 335472 237439 335474
rect 237005 335416 237010 335472
rect 237066 335416 237378 335472
rect 237434 335416 237439 335472
rect 237005 335414 237439 335416
rect 237005 335411 237071 335414
rect 237373 335411 237439 335414
rect 282269 335474 282335 335477
rect 286777 335474 286843 335477
rect 282269 335472 286843 335474
rect 282269 335416 282274 335472
rect 282330 335416 286782 335472
rect 286838 335416 286843 335472
rect 282269 335414 286843 335416
rect 282269 335411 282335 335414
rect 286777 335411 286843 335414
rect 158621 335338 158687 335341
rect 240133 335338 240199 335341
rect 158621 335336 240199 335338
rect 158621 335280 158626 335336
rect 158682 335280 240138 335336
rect 240194 335280 240199 335336
rect 158621 335278 240199 335280
rect 158621 335275 158687 335278
rect 240133 335275 240199 335278
rect 279877 335338 279943 335341
rect 547965 335338 548031 335341
rect 279877 335336 548031 335338
rect 279877 335280 279882 335336
rect 279938 335280 547970 335336
rect 548026 335280 548031 335336
rect 279877 335278 548031 335280
rect 279877 335275 279943 335278
rect 547965 335275 548031 335278
rect 140681 335202 140747 335205
rect 246389 335202 246455 335205
rect 140681 335200 246455 335202
rect 140681 335144 140686 335200
rect 140742 335144 246394 335200
rect 246450 335144 246455 335200
rect 140681 335142 246455 335144
rect 140681 335139 140747 335142
rect 246389 335139 246455 335142
rect 273437 335202 273503 335205
rect 274357 335202 274423 335205
rect 273437 335200 274423 335202
rect 273437 335144 273442 335200
rect 273498 335144 274362 335200
rect 274418 335144 274423 335200
rect 273437 335142 274423 335144
rect 273437 335139 273503 335142
rect 274357 335139 274423 335142
rect 280061 335202 280127 335205
rect 550633 335202 550699 335205
rect 280061 335200 550699 335202
rect 280061 335144 280066 335200
rect 280122 335144 550638 335200
rect 550694 335144 550699 335200
rect 280061 335142 550699 335144
rect 280061 335139 280127 335142
rect 550633 335139 550699 335142
rect 136449 335066 136515 335069
rect 244549 335066 244615 335069
rect 136449 335064 244615 335066
rect 136449 335008 136454 335064
rect 136510 335008 244554 335064
rect 244610 335008 244615 335064
rect 136449 335006 244615 335008
rect 136449 335003 136515 335006
rect 244549 335003 244615 335006
rect 281165 335066 281231 335069
rect 564433 335066 564499 335069
rect 281165 335064 564499 335066
rect 281165 335008 281170 335064
rect 281226 335008 564438 335064
rect 564494 335008 564499 335064
rect 281165 335006 564499 335008
rect 281165 335003 281231 335006
rect 564433 335003 564499 335006
rect 129641 334930 129707 334933
rect 245469 334930 245535 334933
rect 129641 334928 245535 334930
rect 129641 334872 129646 334928
rect 129702 334872 245474 334928
rect 245530 334872 245535 334928
rect 129641 334870 245535 334872
rect 129641 334867 129707 334870
rect 245469 334867 245535 334870
rect 281441 334930 281507 334933
rect 568573 334930 568639 334933
rect 281441 334928 568639 334930
rect 281441 334872 281446 334928
rect 281502 334872 568578 334928
rect 568634 334872 568639 334928
rect 281441 334870 568639 334872
rect 281441 334867 281507 334870
rect 568573 334867 568639 334870
rect 55121 334794 55187 334797
rect 239254 334794 239260 334796
rect 55121 334792 239260 334794
rect 55121 334736 55126 334792
rect 55182 334736 239260 334792
rect 55121 334734 239260 334736
rect 55121 334731 55187 334734
rect 239254 334732 239260 334734
rect 239324 334732 239330 334796
rect 277945 334792 278011 334797
rect 277945 334736 277950 334792
rect 278006 334736 278011 334792
rect 277945 334731 278011 334736
rect 281901 334794 281967 334797
rect 572713 334794 572779 334797
rect 281901 334792 572779 334794
rect 281901 334736 281906 334792
rect 281962 334736 572718 334792
rect 572774 334736 572779 334792
rect 281901 334734 572779 334736
rect 281901 334731 281967 334734
rect 572713 334731 572779 334734
rect 16573 334658 16639 334661
rect 236177 334658 236243 334661
rect 16573 334656 236243 334658
rect 16573 334600 16578 334656
rect 16634 334600 236182 334656
rect 236238 334600 236243 334656
rect 16573 334598 236243 334600
rect 16573 334595 16639 334598
rect 236177 334595 236243 334598
rect 277948 334386 278008 334731
rect 282177 334658 282243 334661
rect 575473 334658 575539 334661
rect 282177 334656 575539 334658
rect 282177 334600 282182 334656
rect 282238 334600 575478 334656
rect 575534 334600 575539 334656
rect 282177 334598 575539 334600
rect 282177 334595 282243 334598
rect 575473 334595 575539 334598
rect 278262 334460 278268 334524
rect 278332 334522 278338 334524
rect 427077 334522 427143 334525
rect 278332 334520 427143 334522
rect 278332 334464 427082 334520
rect 427138 334464 427143 334520
rect 278332 334462 427143 334464
rect 278332 334460 278338 334462
rect 427077 334459 427143 334462
rect 290457 334386 290523 334389
rect 277948 334384 290523 334386
rect 277948 334328 290462 334384
rect 290518 334328 290523 334384
rect 277948 334326 290523 334328
rect 290457 334323 290523 334326
rect 283005 334250 283071 334253
rect 285581 334250 285647 334253
rect 283005 334248 285647 334250
rect 283005 334192 283010 334248
rect 283066 334192 285586 334248
rect 285642 334192 285647 334248
rect 283005 334190 285647 334192
rect 283005 334187 283071 334190
rect 285581 334187 285647 334190
rect 231301 334114 231367 334117
rect 236729 334114 236795 334117
rect 231301 334112 236795 334114
rect 231301 334056 231306 334112
rect 231362 334056 236734 334112
rect 236790 334056 236795 334112
rect 231301 334054 236795 334056
rect 231301 334051 231367 334054
rect 236729 334051 236795 334054
rect 237833 334114 237899 334117
rect 248597 334114 248663 334117
rect 237833 334112 248663 334114
rect 237833 334056 237838 334112
rect 237894 334056 248602 334112
rect 248658 334056 248663 334112
rect 237833 334054 248663 334056
rect 237833 334051 237899 334054
rect 248597 334051 248663 334054
rect 282637 334114 282703 334117
rect 282913 334114 282979 334117
rect 282637 334112 282979 334114
rect 282637 334056 282642 334112
rect 282698 334056 282918 334112
rect 282974 334056 282979 334112
rect 282637 334054 282979 334056
rect 282637 334051 282703 334054
rect 282913 334051 282979 334054
rect 128261 333978 128327 333981
rect 245193 333978 245259 333981
rect 128261 333976 245259 333978
rect 128261 333920 128266 333976
rect 128322 333920 245198 333976
rect 245254 333920 245259 333976
rect 128261 333918 245259 333920
rect 128261 333915 128327 333918
rect 245193 333915 245259 333918
rect 268694 333916 268700 333980
rect 268764 333978 268770 333980
rect 412633 333978 412699 333981
rect 268764 333976 412699 333978
rect 268764 333920 412638 333976
rect 412694 333920 412699 333976
rect 268764 333918 412699 333920
rect 268764 333916 268770 333918
rect 412633 333915 412699 333918
rect 81341 333842 81407 333845
rect 236361 333842 236427 333845
rect 81341 333840 236427 333842
rect 81341 333784 81346 333840
rect 81402 333784 236366 333840
rect 236422 333784 236427 333840
rect 81341 333782 236427 333784
rect 81341 333779 81407 333782
rect 236361 333779 236427 333782
rect 236637 333842 236703 333845
rect 243353 333842 243419 333845
rect 236637 333840 243419 333842
rect 236637 333784 236642 333840
rect 236698 333784 243358 333840
rect 243414 333784 243419 333840
rect 236637 333782 243419 333784
rect 236637 333779 236703 333782
rect 243353 333779 243419 333782
rect 270125 333842 270191 333845
rect 418797 333842 418863 333845
rect 270125 333840 418863 333842
rect 270125 333784 270130 333840
rect 270186 333784 418802 333840
rect 418858 333784 418863 333840
rect 270125 333782 418863 333784
rect 270125 333779 270191 333782
rect 418797 333779 418863 333782
rect 48221 333706 48287 333709
rect 238201 333706 238267 333709
rect 48221 333704 238267 333706
rect 48221 333648 48226 333704
rect 48282 333648 238206 333704
rect 238262 333648 238267 333704
rect 48221 333646 238267 333648
rect 48221 333643 48287 333646
rect 238201 333643 238267 333646
rect 270309 333706 270375 333709
rect 423673 333706 423739 333709
rect 270309 333704 423739 333706
rect 270309 333648 270314 333704
rect 270370 333648 423678 333704
rect 423734 333648 423739 333704
rect 270309 333646 423739 333648
rect 270309 333643 270375 333646
rect 423673 333643 423739 333646
rect 40677 333570 40743 333573
rect 234613 333570 234679 333573
rect 40677 333568 234679 333570
rect 40677 333512 40682 333568
rect 40738 333512 234618 333568
rect 234674 333512 234679 333568
rect 40677 333510 234679 333512
rect 40677 333507 40743 333510
rect 234613 333507 234679 333510
rect 236361 333570 236427 333573
rect 237925 333570 237991 333573
rect 236361 333568 237991 333570
rect 236361 333512 236366 333568
rect 236422 333512 237930 333568
rect 237986 333512 237991 333568
rect 236361 333510 237991 333512
rect 236361 333507 236427 333510
rect 237925 333507 237991 333510
rect 270769 333570 270835 333573
rect 432597 333570 432663 333573
rect 270769 333568 432663 333570
rect 270769 333512 270774 333568
rect 270830 333512 432602 333568
rect 432658 333512 432663 333568
rect 270769 333510 432663 333512
rect 270769 333507 270835 333510
rect 432597 333507 432663 333510
rect 32397 333434 32463 333437
rect 234797 333434 234863 333437
rect 32397 333432 234863 333434
rect 32397 333376 32402 333432
rect 32458 333376 234802 333432
rect 234858 333376 234863 333432
rect 32397 333374 234863 333376
rect 32397 333371 32463 333374
rect 234797 333371 234863 333374
rect 237465 333434 237531 333437
rect 238293 333434 238359 333437
rect 237465 333432 238359 333434
rect 237465 333376 237470 333432
rect 237526 333376 238298 333432
rect 238354 333376 238359 333432
rect 237465 333374 238359 333376
rect 237465 333371 237531 333374
rect 238293 333371 238359 333374
rect 272425 333434 272491 333437
rect 438209 333434 438275 333437
rect 272425 333432 438275 333434
rect 272425 333376 272430 333432
rect 272486 333376 438214 333432
rect 438270 333376 438275 333432
rect 272425 333374 438275 333376
rect 272425 333371 272491 333374
rect 438209 333371 438275 333374
rect 28993 333298 29059 333301
rect 237005 333298 237071 333301
rect 249241 333298 249307 333301
rect 28993 333296 237071 333298
rect 28993 333240 28998 333296
rect 29054 333240 237010 333296
rect 237066 333240 237071 333296
rect 28993 333238 237071 333240
rect 28993 333235 29059 333238
rect 237005 333235 237071 333238
rect 244230 333296 249307 333298
rect 244230 333240 249246 333296
rect 249302 333240 249307 333296
rect 244230 333238 249307 333240
rect 236913 333162 236979 333165
rect 244230 333162 244290 333238
rect 249241 333235 249307 333238
rect 271781 333298 271847 333301
rect 439497 333298 439563 333301
rect 271781 333296 439563 333298
rect 271781 333240 271786 333296
rect 271842 333240 439502 333296
rect 439558 333240 439563 333296
rect 271781 333238 439563 333240
rect 271781 333235 271847 333238
rect 439497 333235 439563 333238
rect 236913 333160 244290 333162
rect 236913 333104 236918 333160
rect 236974 333104 244290 333160
rect 236913 333102 244290 333104
rect 236913 333099 236979 333102
rect 238293 332618 238359 332621
rect 245469 332618 245535 332621
rect 238293 332616 245535 332618
rect 238293 332560 238298 332616
rect 238354 332560 245474 332616
rect 245530 332560 245535 332616
rect 238293 332558 245535 332560
rect 238293 332555 238359 332558
rect 245469 332555 245535 332558
rect 280429 332482 280495 332485
rect 551277 332482 551343 332485
rect 280429 332480 551343 332482
rect -960 332196 480 332436
rect 280429 332424 280434 332480
rect 280490 332424 551282 332480
rect 551338 332424 551343 332480
rect 280429 332422 551343 332424
rect 280429 332419 280495 332422
rect 551277 332419 551343 332422
rect 66161 332346 66227 332349
rect 240409 332346 240475 332349
rect 66161 332344 240475 332346
rect 66161 332288 66166 332344
rect 66222 332288 240414 332344
rect 240470 332288 240475 332344
rect 66161 332286 240475 332288
rect 66161 332283 66227 332286
rect 240409 332283 240475 332286
rect 280705 332346 280771 332349
rect 558177 332346 558243 332349
rect 280705 332344 558243 332346
rect 280705 332288 280710 332344
rect 280766 332288 558182 332344
rect 558238 332288 558243 332344
rect 280705 332286 558243 332288
rect 280705 332283 280771 332286
rect 558177 332283 558243 332286
rect 53097 332210 53163 332213
rect 239213 332210 239279 332213
rect 53097 332208 239279 332210
rect 53097 332152 53102 332208
rect 53158 332152 239218 332208
rect 239274 332152 239279 332208
rect 53097 332150 239279 332152
rect 53097 332147 53163 332150
rect 239213 332147 239279 332150
rect 281349 332210 281415 332213
rect 562317 332210 562383 332213
rect 281349 332208 562383 332210
rect 281349 332152 281354 332208
rect 281410 332152 562322 332208
rect 562378 332152 562383 332208
rect 281349 332150 562383 332152
rect 281349 332147 281415 332150
rect 562317 332147 562383 332150
rect 43437 332074 43503 332077
rect 235441 332074 235507 332077
rect 43437 332072 235507 332074
rect 43437 332016 43442 332072
rect 43498 332016 235446 332072
rect 235502 332016 235507 332072
rect 43437 332014 235507 332016
rect 43437 332011 43503 332014
rect 235441 332011 235507 332014
rect 281625 332074 281691 332077
rect 569217 332074 569283 332077
rect 281625 332072 569283 332074
rect 281625 332016 281630 332072
rect 281686 332016 569222 332072
rect 569278 332016 569283 332072
rect 281625 332014 569283 332016
rect 281625 332011 281691 332014
rect 569217 332011 569283 332014
rect 39297 331938 39363 331941
rect 235165 331938 235231 331941
rect 39297 331936 235231 331938
rect 39297 331880 39302 331936
rect 39358 331880 235170 331936
rect 235226 331880 235231 331936
rect 39297 331878 235231 331880
rect 39297 331875 39363 331878
rect 235165 331875 235231 331878
rect 281993 331938 282059 331941
rect 572805 331938 572871 331941
rect 281993 331936 572871 331938
rect 281993 331880 281998 331936
rect 282054 331880 572810 331936
rect 572866 331880 572871 331936
rect 281993 331878 572871 331880
rect 281993 331875 282059 331878
rect 572805 331875 572871 331878
rect 36537 331802 36603 331805
rect 235073 331802 235139 331805
rect 36537 331800 235139 331802
rect 36537 331744 36542 331800
rect 36598 331744 235078 331800
rect 235134 331744 235139 331800
rect 36537 331742 235139 331744
rect 36537 331739 36603 331742
rect 235073 331739 235139 331742
rect 282361 331802 282427 331805
rect 574737 331802 574803 331805
rect 282361 331800 574803 331802
rect 282361 331744 282366 331800
rect 282422 331744 574742 331800
rect 574798 331744 574803 331800
rect 282361 331742 574803 331744
rect 282361 331739 282427 331742
rect 574737 331739 574803 331742
rect 70301 330850 70367 330853
rect 241145 330850 241211 330853
rect 70301 330848 241211 330850
rect 70301 330792 70306 330848
rect 70362 330792 241150 330848
rect 241206 330792 241211 330848
rect 70301 330790 241211 330792
rect 70301 330787 70367 330790
rect 241145 330787 241211 330790
rect 270401 330850 270467 330853
rect 427813 330850 427879 330853
rect 270401 330848 427879 330850
rect 270401 330792 270406 330848
rect 270462 330792 427818 330848
rect 427874 330792 427879 330848
rect 270401 330790 427879 330792
rect 270401 330787 270467 330790
rect 427813 330787 427879 330790
rect 62021 330714 62087 330717
rect 239949 330714 240015 330717
rect 62021 330712 240015 330714
rect 62021 330656 62026 330712
rect 62082 330656 239954 330712
rect 240010 330656 240015 330712
rect 62021 330654 240015 330656
rect 62021 330651 62087 330654
rect 239949 330651 240015 330654
rect 270585 330714 270651 330717
rect 438853 330714 438919 330717
rect 270585 330712 438919 330714
rect 270585 330656 270590 330712
rect 270646 330656 438858 330712
rect 438914 330656 438919 330712
rect 270585 330654 438919 330656
rect 270585 330651 270651 330654
rect 438853 330651 438919 330654
rect 61377 330578 61443 330581
rect 239765 330578 239831 330581
rect 61377 330576 239831 330578
rect 61377 330520 61382 330576
rect 61438 330520 239770 330576
rect 239826 330520 239831 330576
rect 61377 330518 239831 330520
rect 61377 330515 61443 330518
rect 239765 330515 239831 330518
rect 279233 330578 279299 330581
rect 537017 330578 537083 330581
rect 279233 330576 537083 330578
rect 279233 330520 279238 330576
rect 279294 330520 537022 330576
rect 537078 330520 537083 330576
rect 279233 330518 537083 330520
rect 279233 330515 279299 330518
rect 537017 330515 537083 330518
rect 25497 330442 25563 330445
rect 233325 330442 233391 330445
rect 25497 330440 233391 330442
rect 25497 330384 25502 330440
rect 25558 330384 233330 330440
rect 233386 330384 233391 330440
rect 25497 330382 233391 330384
rect 25497 330379 25563 330382
rect 233325 330379 233391 330382
rect 256141 330442 256207 330445
rect 519537 330442 519603 330445
rect 256141 330440 519603 330442
rect 256141 330384 256146 330440
rect 256202 330384 519542 330440
rect 519598 330384 519603 330440
rect 256141 330382 519603 330384
rect 256141 330379 256207 330382
rect 519537 330379 519603 330382
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 467833 322554 467899 322557
rect 469397 322556 469463 322557
rect 474549 322556 474615 322557
rect 468150 322554 468156 322556
rect 467833 322552 468156 322554
rect 467833 322496 467838 322552
rect 467894 322496 468156 322552
rect 467833 322494 468156 322496
rect 467833 322491 467899 322494
rect 468150 322492 468156 322494
rect 468220 322492 468226 322556
rect 469397 322552 469444 322556
rect 469508 322554 469514 322556
rect 469397 322496 469402 322552
rect 469397 322492 469444 322496
rect 469508 322494 469554 322554
rect 474549 322552 474596 322556
rect 474660 322554 474666 322556
rect 476573 322554 476639 322557
rect 479149 322556 479215 322557
rect 476798 322554 476804 322556
rect 474549 322496 474554 322552
rect 469508 322492 469514 322494
rect 474549 322492 474596 322496
rect 474660 322494 474706 322554
rect 476573 322552 476804 322554
rect 476573 322496 476578 322552
rect 476634 322496 476804 322552
rect 476573 322494 476804 322496
rect 474660 322492 474666 322494
rect 469397 322491 469463 322492
rect 474549 322491 474615 322492
rect 476573 322491 476639 322494
rect 476798 322492 476804 322494
rect 476868 322492 476874 322556
rect 479149 322552 479196 322556
rect 479260 322554 479266 322556
rect 481633 322554 481699 322557
rect 481950 322554 481956 322556
rect 479149 322496 479154 322552
rect 479149 322492 479196 322496
rect 479260 322494 479306 322554
rect 481633 322552 481956 322554
rect 481633 322496 481638 322552
rect 481694 322496 481956 322552
rect 481633 322494 481956 322496
rect 479260 322492 479266 322494
rect 479149 322491 479215 322492
rect 481633 322491 481699 322494
rect 481950 322492 481956 322494
rect 482020 322492 482026 322556
rect 483013 322554 483079 322557
rect 483238 322554 483244 322556
rect 483013 322552 483244 322554
rect 483013 322496 483018 322552
rect 483074 322496 483244 322552
rect 483013 322494 483244 322496
rect 483013 322491 483079 322494
rect 483238 322492 483244 322494
rect 483308 322492 483314 322556
rect 484853 322554 484919 322557
rect 485446 322554 485452 322556
rect 484853 322552 485452 322554
rect 484853 322496 484858 322552
rect 484914 322496 485452 322552
rect 484853 322494 485452 322496
rect 484853 322491 484919 322494
rect 485446 322492 485452 322494
rect 485516 322492 485522 322556
rect 488533 322554 488599 322557
rect 490557 322556 490623 322557
rect 489494 322554 489500 322556
rect 488533 322552 489500 322554
rect 488533 322496 488538 322552
rect 488594 322496 489500 322552
rect 488533 322494 489500 322496
rect 488533 322491 488599 322494
rect 489494 322492 489500 322494
rect 489564 322492 489570 322556
rect 490557 322552 490604 322556
rect 490668 322554 490674 322556
rect 492673 322554 492739 322557
rect 492990 322554 492996 322556
rect 490557 322496 490562 322552
rect 490557 322492 490604 322496
rect 490668 322494 490714 322554
rect 492673 322552 492996 322554
rect 492673 322496 492678 322552
rect 492734 322496 492996 322552
rect 492673 322494 492996 322496
rect 490668 322492 490674 322494
rect 490557 322491 490623 322492
rect 492673 322491 492739 322494
rect 492990 322492 492996 322494
rect 493060 322492 493066 322556
rect 519537 322420 519603 322421
rect 519486 322356 519492 322420
rect 519556 322418 519603 322420
rect 519556 322416 519648 322418
rect 519598 322360 519648 322416
rect 519556 322358 519648 322360
rect 519556 322356 519603 322358
rect 519537 322355 519603 322356
rect 485773 322010 485839 322013
rect 486918 322010 486924 322012
rect 485773 322008 486924 322010
rect 485773 321952 485778 322008
rect 485834 321952 486924 322008
rect 485773 321950 486924 321952
rect 485773 321947 485839 321950
rect 486918 321948 486924 321950
rect 486988 321948 486994 322012
rect 470685 321604 470751 321605
rect 471973 321604 472039 321605
rect 470685 321600 470732 321604
rect 470796 321602 470802 321604
rect 470685 321544 470690 321600
rect 470685 321540 470732 321544
rect 470796 321542 470842 321602
rect 471973 321600 472020 321604
rect 472084 321602 472090 321604
rect 472249 321602 472315 321605
rect 473118 321602 473124 321604
rect 471973 321544 471978 321600
rect 470796 321540 470802 321542
rect 471973 321540 472020 321544
rect 472084 321542 472130 321602
rect 472249 321600 473124 321602
rect 472249 321544 472254 321600
rect 472310 321544 473124 321600
rect 472249 321542 473124 321544
rect 472084 321540 472090 321542
rect 470685 321539 470751 321540
rect 471973 321539 472039 321540
rect 472249 321539 472315 321542
rect 473118 321540 473124 321542
rect 473188 321540 473194 321604
rect 475469 321602 475535 321605
rect 478229 321604 478295 321605
rect 480621 321604 480687 321605
rect 484393 321604 484459 321605
rect 475694 321602 475700 321604
rect 475469 321600 475700 321602
rect 475469 321544 475474 321600
rect 475530 321544 475700 321600
rect 475469 321542 475700 321544
rect 475469 321539 475535 321542
rect 475694 321540 475700 321542
rect 475764 321540 475770 321604
rect 478229 321600 478276 321604
rect 478340 321602 478346 321604
rect 478229 321544 478234 321600
rect 478229 321540 478276 321544
rect 478340 321542 478386 321602
rect 480621 321600 480668 321604
rect 480732 321602 480738 321604
rect 484342 321602 484348 321604
rect 480621 321544 480626 321600
rect 478340 321540 478346 321542
rect 480621 321540 480668 321544
rect 480732 321542 480778 321602
rect 484302 321542 484348 321602
rect 484412 321600 484459 321604
rect 484454 321544 484459 321600
rect 480732 321540 480738 321542
rect 484342 321540 484348 321542
rect 484412 321540 484459 321544
rect 478229 321539 478295 321540
rect 480621 321539 480687 321540
rect 484393 321539 484459 321540
rect 488165 321602 488231 321605
rect 492213 321604 492279 321605
rect 494237 321604 494303 321605
rect 488165 321600 488274 321602
rect 488165 321544 488170 321600
rect 488226 321544 488274 321600
rect 488165 321539 488274 321544
rect 492213 321600 492260 321604
rect 492324 321602 492330 321604
rect 492213 321544 492218 321600
rect 492213 321540 492260 321544
rect 492324 321542 492370 321602
rect 494237 321600 494284 321604
rect 494348 321602 494354 321604
rect 495525 321602 495591 321605
rect 496813 321604 496879 321605
rect 498193 321604 498259 321605
rect 494237 321544 494242 321600
rect 492324 321540 492330 321542
rect 494237 321540 494284 321544
rect 494348 321542 494394 321602
rect 495525 321600 495634 321602
rect 495525 321544 495530 321600
rect 495586 321544 495634 321600
rect 494348 321540 494354 321542
rect 492213 321539 492279 321540
rect 494237 321539 494303 321540
rect 495525 321539 495634 321544
rect 496813 321600 496860 321604
rect 496924 321602 496930 321604
rect 498142 321602 498148 321604
rect 496813 321544 496818 321600
rect 496813 321540 496860 321544
rect 496924 321542 496970 321602
rect 498102 321542 498148 321602
rect 498212 321600 498259 321604
rect 498254 321544 498259 321600
rect 496924 321540 496930 321542
rect 498142 321540 498148 321542
rect 498212 321540 498259 321544
rect 496813 321539 496879 321540
rect 498193 321539 498259 321540
rect 498653 321602 498719 321605
rect 500677 321604 500743 321605
rect 498653 321600 499314 321602
rect 498653 321544 498658 321600
rect 498714 321544 499314 321600
rect 498653 321542 499314 321544
rect 498653 321539 498719 321542
rect 488214 321332 488274 321539
rect 495574 321332 495634 321539
rect 499254 321332 499314 321542
rect 500677 321600 500724 321604
rect 500788 321602 500794 321604
rect 501045 321602 501111 321605
rect 503253 321604 503319 321605
rect 504173 321604 504239 321605
rect 505461 321604 505527 321605
rect 506933 321604 506999 321605
rect 530025 321604 530091 321605
rect 501822 321602 501828 321604
rect 500677 321544 500682 321600
rect 500677 321540 500724 321544
rect 500788 321542 500834 321602
rect 501045 321600 501828 321602
rect 501045 321544 501050 321600
rect 501106 321544 501828 321600
rect 501045 321542 501828 321544
rect 500788 321540 500794 321542
rect 500677 321539 500743 321540
rect 501045 321539 501111 321542
rect 501822 321540 501828 321542
rect 501892 321540 501898 321604
rect 503253 321600 503300 321604
rect 503364 321602 503370 321604
rect 503253 321544 503258 321600
rect 503253 321540 503300 321544
rect 503364 321542 503410 321602
rect 504173 321600 504220 321604
rect 504284 321602 504290 321604
rect 504173 321544 504178 321600
rect 503364 321540 503370 321542
rect 504173 321540 504220 321544
rect 504284 321542 504330 321602
rect 505461 321600 505508 321604
rect 505572 321602 505578 321604
rect 505461 321544 505466 321600
rect 504284 321540 504290 321542
rect 505461 321540 505508 321544
rect 505572 321542 505618 321602
rect 506933 321600 506980 321604
rect 507044 321602 507050 321604
rect 529974 321602 529980 321604
rect 506933 321544 506938 321600
rect 505572 321540 505578 321542
rect 506933 321540 506980 321544
rect 507044 321542 507090 321602
rect 529934 321542 529980 321602
rect 530044 321600 530091 321604
rect 530086 321544 530091 321600
rect 507044 321540 507050 321542
rect 529974 321540 529980 321542
rect 530044 321540 530091 321544
rect 503253 321539 503319 321540
rect 504173 321539 504239 321540
rect 505461 321539 505527 321540
rect 506933 321539 506999 321540
rect 530025 321539 530091 321540
rect 488206 321268 488212 321332
rect 488276 321268 488282 321332
rect 495566 321268 495572 321332
rect 495636 321268 495642 321332
rect 499246 321268 499252 321332
rect 499316 321268 499322 321332
rect -960 319290 480 319380
rect 3509 319290 3575 319293
rect -960 319288 3575 319290
rect -960 319232 3514 319288
rect 3570 319232 3575 319288
rect -960 319230 3575 319232
rect -960 319140 480 319230
rect 3509 319227 3575 319230
rect 538305 316570 538371 316573
rect 536422 316568 538371 316570
rect 536422 316512 538310 316568
rect 538366 316512 538371 316568
rect 536422 316510 538371 316512
rect 536422 316500 536482 316510
rect 538305 316507 538371 316510
rect 535900 316440 536482 316500
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3049 293178 3115 293181
rect -960 293176 3115 293178
rect -960 293120 3054 293176
rect 3110 293120 3115 293176
rect -960 293118 3115 293120
rect -960 293028 480 293118
rect 3049 293115 3115 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 437473 274274 437539 274277
rect 438761 274274 438827 274277
rect 437473 274272 439882 274274
rect 437473 274216 437478 274272
rect 437534 274216 438766 274272
rect 438822 274216 439882 274272
rect 437473 274214 439882 274216
rect 437473 274211 437539 274214
rect 438761 274211 438827 274214
rect 439822 274204 439882 274214
rect 439822 274144 440032 274204
rect 439822 272920 440032 272980
rect 436645 272914 436711 272917
rect 437381 272914 437447 272917
rect 439822 272914 439882 272920
rect 436645 272912 439882 272914
rect 436645 272856 436650 272912
rect 436706 272856 437386 272912
rect 437442 272856 439882 272912
rect 436645 272854 439882 272856
rect 436645 272851 436711 272854
rect 437381 272851 437447 272854
rect 579981 272234 580047 272237
rect 583520 272234 584960 272324
rect 579981 272232 584960 272234
rect 579981 272176 579986 272232
rect 580042 272176 584960 272232
rect 579981 272174 584960 272176
rect 579981 272171 580047 272174
rect 583520 272084 584960 272174
rect 436829 271282 436895 271285
rect 438669 271282 438735 271285
rect 436829 271280 439882 271282
rect 436829 271224 436834 271280
rect 436890 271224 438674 271280
rect 438730 271224 439882 271280
rect 436829 271222 439882 271224
rect 436829 271219 436895 271222
rect 438669 271219 438735 271222
rect 439822 271212 439882 271222
rect 439822 271152 440032 271212
rect 436829 270194 436895 270197
rect 438577 270194 438643 270197
rect 436829 270192 439882 270194
rect 436829 270136 436834 270192
rect 436890 270136 438582 270192
rect 438638 270136 439882 270192
rect 436829 270134 439882 270136
rect 436829 270131 436895 270134
rect 438577 270131 438643 270134
rect 439822 270124 439882 270134
rect 439822 270064 440032 270124
rect 439822 268432 440032 268492
rect 437289 268426 437355 268429
rect 439822 268426 439882 268432
rect 437289 268424 439882 268426
rect 437289 268368 437294 268424
rect 437350 268368 439882 268424
rect 437289 268366 439882 268368
rect 437289 268363 437355 268366
rect 439454 267480 440032 267540
rect 436093 267474 436159 267477
rect 439454 267474 439514 267480
rect 436093 267472 439514 267474
rect 436093 267416 436098 267472
rect 436154 267416 439514 267472
rect 436093 267414 439514 267416
rect 436093 267411 436159 267414
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 439822 265712 440032 265772
rect 437197 265706 437263 265709
rect 439822 265706 439882 265712
rect 437197 265704 439882 265706
rect 437197 265648 437202 265704
rect 437258 265648 439882 265704
rect 437197 265646 439882 265648
rect 437197 265643 437263 265646
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 535900 256600 536482 256660
rect 536422 256594 536482 256600
rect 538305 256594 538371 256597
rect 536422 256592 538371 256594
rect 536422 256536 538310 256592
rect 538366 256536 538371 256592
rect 536422 256534 538371 256536
rect 538305 256531 538371 256534
rect 535900 254968 536482 255028
rect 536422 254962 536482 254968
rect 538489 254962 538555 254965
rect 536422 254960 538555 254962
rect 536422 254904 538494 254960
rect 538550 254904 538555 254960
rect 536422 254902 538555 254904
rect 538489 254899 538555 254902
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 535900 253608 536482 253668
rect 536422 253602 536482 253608
rect 538397 253602 538463 253605
rect 536422 253600 538463 253602
rect 536422 253544 538402 253600
rect 538458 253544 538463 253600
rect 536422 253542 538463 253544
rect 538397 253539 538463 253542
rect 436093 247346 436159 247349
rect 436093 247344 439514 247346
rect 436093 247288 436098 247344
rect 436154 247288 439514 247344
rect 436093 247286 439514 247288
rect 436093 247283 436159 247286
rect 439454 247276 439514 247286
rect 439454 247216 440032 247276
rect 439454 245584 440032 245644
rect 436737 245578 436803 245581
rect 439454 245578 439514 245584
rect 436737 245576 439514 245578
rect 436737 245520 436742 245576
rect 436798 245520 439514 245576
rect 436737 245518 439514 245520
rect 580809 245578 580875 245581
rect 583520 245578 584960 245668
rect 580809 245576 584960 245578
rect 580809 245520 580814 245576
rect 580870 245520 584960 245576
rect 580809 245518 584960 245520
rect 436737 245515 436803 245518
rect 580809 245515 580875 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 272701 239866 272767 239869
rect 445569 239866 445635 239869
rect 445845 239868 445911 239869
rect 445845 239866 445854 239868
rect 272701 239864 445635 239866
rect 272701 239808 272706 239864
rect 272762 239808 445574 239864
rect 445630 239808 445635 239864
rect 272701 239806 445635 239808
rect 445762 239864 445854 239866
rect 445762 239808 445850 239864
rect 445762 239806 445854 239808
rect 272701 239803 272767 239806
rect 445569 239803 445635 239806
rect 445845 239804 445854 239806
rect 445918 239804 445924 239868
rect 451089 239866 451155 239869
rect 452745 239866 452811 239869
rect 451089 239864 452811 239866
rect 451089 239808 451094 239864
rect 451150 239808 452750 239864
rect 452806 239808 452811 239864
rect 451089 239806 452811 239808
rect 445845 239803 445911 239804
rect 451089 239803 451155 239806
rect 452745 239803 452811 239806
rect 460933 239866 460999 239869
rect 522665 239868 522731 239869
rect 469240 239866 469246 239868
rect 460933 239864 469246 239866
rect 460933 239808 460938 239864
rect 460994 239808 469246 239864
rect 460933 239806 469246 239808
rect 460933 239803 460999 239806
rect 469240 239804 469246 239806
rect 469310 239804 469316 239868
rect 522665 239866 522694 239868
rect 522602 239864 522694 239866
rect 522602 239808 522670 239864
rect 522602 239806 522694 239808
rect 522665 239804 522694 239806
rect 522758 239804 522764 239868
rect 522960 239804 522966 239868
rect 523030 239866 523036 239868
rect 523125 239866 523191 239869
rect 523030 239864 523191 239866
rect 523030 239808 523130 239864
rect 523186 239808 523191 239864
rect 523030 239806 523191 239808
rect 523030 239804 523036 239806
rect 522665 239803 522731 239804
rect 523125 239803 523191 239806
rect 275185 239730 275251 239733
rect 462405 239730 462471 239733
rect 473169 239732 473235 239733
rect 475653 239732 475719 239733
rect 523125 239732 523191 239733
rect 473169 239730 473190 239732
rect 275185 239728 462471 239730
rect 275185 239672 275190 239728
rect 275246 239672 462410 239728
rect 462466 239672 462471 239728
rect 275185 239670 462471 239672
rect 473098 239728 473190 239730
rect 473098 239672 473174 239728
rect 473098 239670 473190 239672
rect 275185 239667 275251 239670
rect 462405 239667 462471 239670
rect 473169 239668 473190 239670
rect 473254 239668 473260 239732
rect 475632 239668 475638 239732
rect 475702 239730 475719 239732
rect 475702 239728 475794 239730
rect 475714 239672 475794 239728
rect 475702 239670 475794 239672
rect 475702 239668 475719 239670
rect 523096 239668 523102 239732
rect 523166 239730 523191 239732
rect 523166 239728 523258 239730
rect 523186 239672 523258 239728
rect 523166 239670 523258 239672
rect 523166 239668 523191 239670
rect 473169 239667 473235 239668
rect 475653 239667 475719 239668
rect 523125 239667 523191 239668
rect 276381 239594 276447 239597
rect 465257 239594 465323 239597
rect 471973 239596 472039 239597
rect 479333 239596 479399 239597
rect 487889 239596 487955 239597
rect 495617 239596 495683 239597
rect 496813 239596 496879 239597
rect 500493 239596 500559 239597
rect 501873 239596 501939 239597
rect 503069 239596 503135 239597
rect 505553 239596 505619 239597
rect 506749 239596 506815 239597
rect 276381 239592 465323 239594
rect 276381 239536 276386 239592
rect 276442 239536 465262 239592
rect 465318 239536 465323 239592
rect 276381 239534 465323 239536
rect 276381 239531 276447 239534
rect 465257 239531 465323 239534
rect 471960 239532 471966 239596
rect 472030 239594 472039 239596
rect 472030 239592 472122 239594
rect 472034 239536 472122 239592
rect 472030 239534 472122 239536
rect 472030 239532 472039 239534
rect 473302 239532 473308 239596
rect 473372 239594 473378 239596
rect 474408 239594 474414 239596
rect 473372 239534 474414 239594
rect 473372 239532 473378 239534
rect 474408 239532 474414 239534
rect 474478 239532 474484 239596
rect 479304 239532 479310 239596
rect 479374 239594 479399 239596
rect 479374 239592 479466 239594
rect 479394 239536 479466 239592
rect 479374 239534 479466 239536
rect 479374 239532 479399 239534
rect 487872 239532 487878 239596
rect 487942 239594 487955 239596
rect 487942 239592 488034 239594
rect 487950 239536 488034 239592
rect 487942 239534 488034 239536
rect 487942 239532 487955 239534
rect 492990 239532 492996 239596
rect 493060 239594 493066 239596
rect 493992 239594 493998 239596
rect 493060 239534 493998 239594
rect 493060 239532 493066 239534
rect 493992 239532 493998 239534
rect 494062 239532 494068 239596
rect 495617 239594 495630 239596
rect 495538 239592 495630 239594
rect 495538 239536 495622 239592
rect 495538 239534 495630 239536
rect 495617 239532 495630 239534
rect 495694 239532 495700 239596
rect 496813 239594 496854 239596
rect 496762 239592 496854 239594
rect 496762 239536 496818 239592
rect 496762 239534 496854 239536
rect 496813 239532 496854 239534
rect 496918 239532 496924 239596
rect 500493 239594 500526 239596
rect 500434 239592 500526 239594
rect 500434 239536 500498 239592
rect 500434 239534 500526 239536
rect 500493 239532 500526 239534
rect 500590 239532 500596 239596
rect 501873 239594 501886 239596
rect 501794 239592 501886 239594
rect 501794 239536 501878 239592
rect 501794 239534 501886 239536
rect 501873 239532 501886 239534
rect 501950 239532 501956 239596
rect 503069 239594 503110 239596
rect 503018 239592 503110 239594
rect 503018 239536 503074 239592
rect 503018 239534 503110 239536
rect 503069 239532 503110 239534
rect 503174 239532 503180 239596
rect 505552 239594 505558 239596
rect 505466 239534 505558 239594
rect 505552 239532 505558 239534
rect 505622 239532 505628 239596
rect 506749 239594 506782 239596
rect 506690 239592 506782 239594
rect 506690 239536 506754 239592
rect 506690 239534 506782 239536
rect 506749 239532 506782 239534
rect 506846 239532 506852 239596
rect 471973 239531 472039 239532
rect 479333 239531 479399 239532
rect 487889 239531 487955 239532
rect 495617 239531 495683 239532
rect 496813 239531 496879 239532
rect 500493 239531 500559 239532
rect 501873 239531 501939 239532
rect 503069 239531 503135 239532
rect 505553 239531 505619 239532
rect 506749 239531 506815 239532
rect 273713 239458 273779 239461
rect 468477 239458 468543 239461
rect 273713 239456 468543 239458
rect 273713 239400 273718 239456
rect 273774 239400 468482 239456
rect 468538 239400 468543 239456
rect 273713 239398 468543 239400
rect 273713 239395 273779 239398
rect 468477 239395 468543 239398
rect 445661 239322 445727 239325
rect 451089 239322 451155 239325
rect 445661 239320 451155 239322
rect 445661 239264 445666 239320
rect 445722 239264 451094 239320
rect 451150 239264 451155 239320
rect 445661 239262 451155 239264
rect 445661 239259 445727 239262
rect 451089 239259 451155 239262
rect 452561 239322 452627 239325
rect 461025 239322 461091 239325
rect 452561 239320 461091 239322
rect 452561 239264 452566 239320
rect 452622 239264 461030 239320
rect 461086 239264 461091 239320
rect 452561 239262 461091 239264
rect 452561 239259 452627 239262
rect 461025 239259 461091 239262
rect 445569 239186 445635 239189
rect 452653 239186 452719 239189
rect 445569 239184 452719 239186
rect 445569 239128 445574 239184
rect 445630 239128 452658 239184
rect 452714 239128 452719 239184
rect 445569 239126 452719 239128
rect 445569 239123 445635 239126
rect 452653 239123 452719 239126
rect 455454 239124 455460 239188
rect 455524 239186 455530 239188
rect 537109 239186 537175 239189
rect 455524 239184 537175 239186
rect 455524 239128 537114 239184
rect 537170 239128 537175 239184
rect 455524 239126 537175 239128
rect 455524 239124 455530 239126
rect 537109 239123 537175 239126
rect 254669 239050 254735 239053
rect 457846 239050 457852 239052
rect 254669 239048 457852 239050
rect 254669 238992 254674 239048
rect 254730 238992 457852 239048
rect 254669 238990 457852 238992
rect 254669 238987 254735 238990
rect 457846 238988 457852 238990
rect 457916 238988 457922 239052
rect 235349 238914 235415 238917
rect 456742 238914 456748 238916
rect 235349 238912 456748 238914
rect 235349 238856 235354 238912
rect 235410 238856 456748 238912
rect 235349 238854 456748 238856
rect 235349 238851 235415 238854
rect 456742 238852 456748 238854
rect 456812 238852 456818 238916
rect 236729 238778 236795 238781
rect 459134 238778 459140 238780
rect 236729 238776 459140 238778
rect 236729 238720 236734 238776
rect 236790 238720 459140 238776
rect 236729 238718 459140 238720
rect 236729 238715 236795 238718
rect 459134 238716 459140 238718
rect 459204 238716 459210 238780
rect 477358 238718 477970 238778
rect 234153 238642 234219 238645
rect 477358 238642 477418 238718
rect 477677 238644 477743 238645
rect 477677 238642 477724 238644
rect 234153 238640 477418 238642
rect 234153 238584 234158 238640
rect 234214 238584 477418 238640
rect 234153 238582 477418 238584
rect 477632 238640 477724 238642
rect 477632 238584 477682 238640
rect 477632 238582 477724 238584
rect 234153 238579 234219 238582
rect 477677 238580 477724 238582
rect 477788 238580 477794 238644
rect 477910 238642 477970 238718
rect 483381 238644 483447 238645
rect 484393 238644 484459 238645
rect 481398 238642 481404 238644
rect 477910 238582 481404 238642
rect 481398 238580 481404 238582
rect 481468 238580 481474 238644
rect 483381 238642 483428 238644
rect 483336 238640 483428 238642
rect 483336 238584 483386 238640
rect 483336 238582 483428 238584
rect 483381 238580 483428 238582
rect 483492 238580 483498 238644
rect 484342 238580 484348 238644
rect 484412 238642 484459 238644
rect 485405 238644 485471 238645
rect 485405 238642 485452 238644
rect 484412 238640 484504 238642
rect 484454 238584 484504 238640
rect 484412 238582 484504 238584
rect 485360 238640 485452 238642
rect 485360 238584 485410 238640
rect 485360 238582 485452 238584
rect 484412 238580 484459 238582
rect 477677 238579 477743 238580
rect 483381 238579 483447 238580
rect 484393 238579 484459 238580
rect 485405 238580 485452 238582
rect 485516 238580 485522 238644
rect 485405 238579 485471 238580
rect 234061 238506 234127 238509
rect 482277 238508 482343 238509
rect 484853 238508 484919 238509
rect 478822 238506 478828 238508
rect 234061 238504 478828 238506
rect 234061 238448 234066 238504
rect 234122 238448 478828 238504
rect 234061 238446 478828 238448
rect 234061 238443 234127 238446
rect 478822 238444 478828 238446
rect 478892 238444 478898 238508
rect 482277 238506 482324 238508
rect 482232 238504 482324 238506
rect 482232 238448 482282 238504
rect 482232 238446 482324 238448
rect 482277 238444 482324 238446
rect 482388 238444 482394 238508
rect 484853 238506 484900 238508
rect 484808 238504 484900 238506
rect 484808 238448 484858 238504
rect 484808 238446 484900 238448
rect 484853 238444 484900 238446
rect 484964 238444 484970 238508
rect 482277 238443 482343 238444
rect 484853 238443 484919 238444
rect 233877 238370 233943 238373
rect 476573 238372 476639 238373
rect 480621 238372 480687 238373
rect 481725 238372 481791 238373
rect 485957 238372 486023 238373
rect 488165 238372 488231 238373
rect 474038 238370 474044 238372
rect 233877 238368 474044 238370
rect 233877 238312 233882 238368
rect 233938 238312 474044 238368
rect 233877 238310 474044 238312
rect 233877 238307 233943 238310
rect 474038 238308 474044 238310
rect 474108 238308 474114 238372
rect 476573 238370 476620 238372
rect 476528 238368 476620 238370
rect 476528 238312 476578 238368
rect 476528 238310 476620 238312
rect 476573 238308 476620 238310
rect 476684 238308 476690 238372
rect 480621 238370 480668 238372
rect 480576 238368 480668 238370
rect 480576 238312 480626 238368
rect 480576 238310 480668 238312
rect 480621 238308 480668 238310
rect 480732 238308 480738 238372
rect 481725 238370 481772 238372
rect 481680 238368 481772 238370
rect 481680 238312 481730 238368
rect 481680 238310 481772 238312
rect 481725 238308 481772 238310
rect 481836 238308 481842 238372
rect 485957 238370 486004 238372
rect 485912 238368 486004 238370
rect 485912 238312 485962 238368
rect 485912 238310 486004 238312
rect 485957 238308 486004 238310
rect 486068 238308 486074 238372
rect 488165 238370 488212 238372
rect 488120 238368 488212 238370
rect 488120 238312 488170 238368
rect 488120 238310 488212 238312
rect 488165 238308 488212 238310
rect 488276 238308 488282 238372
rect 476573 238307 476639 238308
rect 480621 238307 480687 238308
rect 481725 238307 481791 238308
rect 485957 238307 486023 238308
rect 488165 238307 488231 238308
rect 293217 238234 293283 238237
rect 491661 238236 491727 238237
rect 492765 238236 492831 238237
rect 495157 238236 495223 238237
rect 490782 238234 490788 238236
rect 293217 238232 490788 238234
rect 293217 238176 293222 238232
rect 293278 238176 490788 238232
rect 293217 238174 490788 238176
rect 293217 238171 293283 238174
rect 490782 238172 490788 238174
rect 490852 238172 490858 238236
rect 491661 238234 491708 238236
rect 491616 238232 491708 238234
rect 491616 238176 491666 238232
rect 491616 238174 491708 238176
rect 491661 238172 491708 238174
rect 491772 238172 491778 238236
rect 492765 238234 492812 238236
rect 492720 238232 492812 238234
rect 492720 238176 492770 238232
rect 492720 238174 492812 238176
rect 492765 238172 492812 238174
rect 492876 238172 492882 238236
rect 495157 238234 495204 238236
rect 495112 238232 495204 238234
rect 495112 238176 495162 238232
rect 495112 238174 495204 238176
rect 495157 238172 495204 238174
rect 495268 238172 495274 238236
rect 491661 238171 491727 238172
rect 492765 238171 492831 238172
rect 495157 238171 495223 238172
rect 437289 238098 437355 238101
rect 538397 238098 538463 238101
rect 437289 238096 538463 238098
rect 437289 238040 437294 238096
rect 437350 238040 538402 238096
rect 538458 238040 538463 238096
rect 437289 238038 538463 238040
rect 437289 238035 437355 238038
rect 538397 238035 538463 238038
rect 437197 237962 437263 237965
rect 538305 237962 538371 237965
rect 437197 237960 538371 237962
rect 437197 237904 437202 237960
rect 437258 237904 538310 237960
rect 538366 237904 538371 237960
rect 437197 237902 538371 237904
rect 437197 237899 437263 237902
rect 538305 237899 538371 237902
rect 439681 237826 439747 237829
rect 497590 237826 497596 237828
rect 439681 237824 497596 237826
rect 439681 237768 439686 237824
rect 439742 237768 497596 237824
rect 439681 237766 497596 237768
rect 439681 237763 439747 237766
rect 497590 237764 497596 237766
rect 497660 237764 497666 237828
rect 467189 237692 467255 237693
rect 467833 237692 467899 237693
rect 467189 237690 467236 237692
rect 467144 237688 467236 237690
rect 467144 237632 467194 237688
rect 467144 237630 467236 237632
rect 467189 237628 467236 237630
rect 467300 237628 467306 237692
rect 467782 237628 467788 237692
rect 467852 237690 467899 237692
rect 467852 237688 467944 237690
rect 467894 237632 467944 237688
rect 467852 237630 467944 237632
rect 467852 237628 467899 237630
rect 467189 237627 467255 237628
rect 467833 237627 467899 237628
rect 462313 237282 462379 237285
rect 463693 237284 463759 237285
rect 462630 237282 462636 237284
rect 462313 237280 462636 237282
rect 462313 237224 462318 237280
rect 462374 237224 462636 237280
rect 462313 237222 462636 237224
rect 462313 237219 462379 237222
rect 462630 237220 462636 237222
rect 462700 237220 462706 237284
rect 463693 237282 463740 237284
rect 463648 237280 463740 237282
rect 463648 237224 463698 237280
rect 463648 237222 463740 237224
rect 463693 237220 463740 237222
rect 463804 237220 463810 237284
rect 465073 237282 465139 237285
rect 466126 237282 466132 237284
rect 465073 237280 466132 237282
rect 465073 237224 465078 237280
rect 465134 237224 466132 237280
rect 465073 237222 466132 237224
rect 463693 237219 463759 237220
rect 465073 237219 465139 237222
rect 466126 237220 466132 237222
rect 466196 237220 466202 237284
rect 467833 237282 467899 237285
rect 468334 237282 468340 237284
rect 467833 237280 468340 237282
rect 467833 237224 467838 237280
rect 467894 237224 468340 237280
rect 467833 237222 468340 237224
rect 467833 237219 467899 237222
rect 468334 237220 468340 237222
rect 468404 237220 468410 237284
rect 469213 237282 469279 237285
rect 469622 237282 469628 237284
rect 469213 237280 469628 237282
rect 469213 237224 469218 237280
rect 469274 237224 469628 237280
rect 469213 237222 469628 237224
rect 469213 237219 469279 237222
rect 469622 237220 469628 237222
rect 469692 237220 469698 237284
rect 470593 237282 470659 237285
rect 470726 237282 470732 237284
rect 470593 237280 470732 237282
rect 470593 237224 470598 237280
rect 470654 237224 470732 237280
rect 470593 237222 470732 237224
rect 470593 237219 470659 237222
rect 470726 237220 470732 237222
rect 470796 237220 470802 237284
rect 485773 237282 485839 237285
rect 487102 237282 487108 237284
rect 485773 237280 487108 237282
rect 485773 237224 485778 237280
rect 485834 237224 487108 237280
rect 485773 237222 487108 237224
rect 485773 237219 485839 237222
rect 487102 237220 487108 237222
rect 487172 237220 487178 237284
rect 498193 237282 498259 237285
rect 498694 237282 498700 237284
rect 498193 237280 498700 237282
rect 498193 237224 498198 237280
rect 498254 237224 498700 237280
rect 498193 237222 498700 237224
rect 498193 237219 498259 237222
rect 498694 237220 498700 237222
rect 498764 237220 498770 237284
rect 503713 237282 503779 237285
rect 504214 237282 504220 237284
rect 503713 237280 504220 237282
rect 503713 237224 503718 237280
rect 503774 237224 504220 237280
rect 503713 237222 504220 237224
rect 503713 237219 503779 237222
rect 504214 237220 504220 237222
rect 504284 237220 504290 237284
rect 521653 237282 521719 237285
rect 522798 237282 522804 237284
rect 521653 237280 522804 237282
rect 521653 237224 521658 237280
rect 521714 237224 522804 237280
rect 521653 237222 522804 237224
rect 521653 237219 521719 237222
rect 522798 237220 522804 237222
rect 522868 237220 522874 237284
rect 233969 237146 234035 237149
rect 483054 237146 483060 237148
rect 233969 237144 483060 237146
rect 233969 237088 233974 237144
rect 234030 237088 483060 237144
rect 233969 237086 483060 237088
rect 233969 237083 234035 237086
rect 483054 237084 483060 237086
rect 483124 237084 483130 237148
rect 490281 237146 490347 237149
rect 490598 237146 490604 237148
rect 490281 237144 490604 237146
rect 490281 237088 490286 237144
rect 490342 237088 490604 237144
rect 490281 237086 490604 237088
rect 490281 237083 490347 237086
rect 490598 237084 490604 237086
rect 490668 237084 490674 237148
rect 492673 237146 492739 237149
rect 493174 237146 493180 237148
rect 492673 237144 493180 237146
rect 492673 237088 492678 237144
rect 492734 237088 493180 237144
rect 492673 237086 493180 237088
rect 492673 237083 492739 237086
rect 493174 237084 493180 237086
rect 493244 237084 493250 237148
rect 494053 237146 494119 237149
rect 494278 237146 494284 237148
rect 494053 237144 494284 237146
rect 494053 237088 494058 237144
rect 494114 237088 494284 237144
rect 494053 237086 494284 237088
rect 494053 237083 494119 237086
rect 494278 237084 494284 237086
rect 494348 237084 494354 237148
rect 234245 237010 234311 237013
rect 491293 237012 491359 237013
rect 480294 237010 480300 237012
rect 234245 237008 480300 237010
rect 234245 236952 234250 237008
rect 234306 236952 480300 237008
rect 234245 236950 480300 236952
rect 234245 236947 234311 236950
rect 480294 236948 480300 236950
rect 480364 236948 480370 237012
rect 491293 237010 491340 237012
rect 491248 237008 491340 237010
rect 491248 236952 491298 237008
rect 491248 236950 491340 236952
rect 491293 236948 491340 236950
rect 491404 236948 491410 237012
rect 491293 236947 491359 236948
rect 249241 236874 249307 236877
rect 460054 236874 460060 236876
rect 249241 236872 460060 236874
rect 249241 236816 249246 236872
rect 249302 236816 460060 236872
rect 249241 236814 460060 236816
rect 249241 236811 249307 236814
rect 460054 236812 460060 236814
rect 460124 236812 460130 236876
rect 461117 236874 461183 236877
rect 465073 236876 465139 236877
rect 461342 236874 461348 236876
rect 461117 236872 461348 236874
rect 461117 236816 461122 236872
rect 461178 236816 461348 236872
rect 461117 236814 461348 236816
rect 461117 236811 461183 236814
rect 461342 236812 461348 236814
rect 461412 236812 461418 236876
rect 465022 236812 465028 236876
rect 465092 236874 465139 236876
rect 471973 236874 472039 236877
rect 473353 236876 473419 236877
rect 472934 236874 472940 236876
rect 465092 236872 465184 236874
rect 465134 236816 465184 236872
rect 465092 236814 465184 236816
rect 471973 236872 472940 236874
rect 471973 236816 471978 236872
rect 472034 236816 472940 236872
rect 471973 236814 472940 236816
rect 465092 236812 465139 236814
rect 465073 236811 465139 236812
rect 471973 236811 472039 236814
rect 472934 236812 472940 236814
rect 473004 236812 473010 236876
rect 473302 236812 473308 236876
rect 473372 236874 473419 236876
rect 474733 236874 474799 236877
rect 475326 236874 475332 236876
rect 473372 236872 473464 236874
rect 473414 236816 473464 236872
rect 473372 236814 473464 236816
rect 474733 236872 475332 236874
rect 474733 236816 474738 236872
rect 474794 236816 475332 236872
rect 474733 236814 475332 236816
rect 473372 236812 473419 236814
rect 473353 236811 473419 236812
rect 474733 236811 474799 236814
rect 475326 236812 475332 236814
rect 475396 236812 475402 236876
rect 476113 236874 476179 236877
rect 476798 236874 476804 236876
rect 476113 236872 476804 236874
rect 476113 236816 476118 236872
rect 476174 236816 476804 236872
rect 476113 236814 476804 236816
rect 476113 236811 476179 236814
rect 476798 236812 476804 236814
rect 476868 236812 476874 236876
rect 485773 236874 485839 236877
rect 486550 236874 486556 236876
rect 485773 236872 486556 236874
rect 485773 236816 485778 236872
rect 485834 236816 486556 236872
rect 485773 236814 486556 236816
rect 485773 236811 485839 236814
rect 486550 236812 486556 236814
rect 486620 236812 486626 236876
rect 488533 236874 488599 236877
rect 489310 236874 489316 236876
rect 488533 236872 489316 236874
rect 488533 236816 488538 236872
rect 488594 236816 489316 236872
rect 488533 236814 489316 236816
rect 488533 236811 488599 236814
rect 489310 236812 489316 236814
rect 489380 236812 489386 236876
rect 293309 236738 293375 236741
rect 492990 236738 492996 236740
rect 293309 236736 492996 236738
rect 293309 236680 293314 236736
rect 293370 236680 492996 236736
rect 293309 236678 492996 236680
rect 293309 236675 293375 236678
rect 492990 236676 492996 236678
rect 493060 236676 493066 236740
rect 297633 236602 297699 236605
rect 497774 236602 497780 236604
rect 297633 236600 497780 236602
rect 297633 236544 297638 236600
rect 297694 236544 497780 236600
rect 297633 236542 497780 236544
rect 297633 236539 297699 236542
rect 497774 236540 497780 236542
rect 497844 236540 497850 236604
rect 234337 236466 234403 236469
rect 489126 236466 489132 236468
rect 234337 236464 489132 236466
rect 234337 236408 234342 236464
rect 234398 236408 489132 236464
rect 234337 236406 489132 236408
rect 234337 236403 234403 236406
rect 489126 236404 489132 236406
rect 489196 236404 489202 236468
rect 470869 236330 470935 236333
rect 471830 236330 471836 236332
rect 470869 236328 471836 236330
rect 470869 236272 470874 236328
rect 470930 236272 471836 236328
rect 470869 236270 471836 236272
rect 470869 236267 470935 236270
rect 471830 236268 471836 236270
rect 471900 236268 471906 236332
rect 469213 236196 469279 236197
rect 469213 236194 469260 236196
rect 469168 236192 469260 236194
rect 469168 236136 469218 236192
rect 469168 236134 469260 236136
rect 469213 236132 469260 236134
rect 469324 236132 469330 236196
rect 477493 236194 477559 236197
rect 478086 236194 478092 236196
rect 477493 236192 478092 236194
rect 477493 236136 477498 236192
rect 477554 236136 478092 236192
rect 477493 236134 478092 236136
rect 469213 236131 469279 236132
rect 477493 236131 477559 236134
rect 478086 236132 478092 236134
rect 478156 236132 478162 236196
rect 495433 236194 495499 236197
rect 496486 236194 496492 236196
rect 495433 236192 496492 236194
rect 495433 236136 495438 236192
rect 495494 236136 496492 236192
rect 495433 236134 496492 236136
rect 495433 236131 495499 236134
rect 496486 236132 496492 236134
rect 496556 236132 496562 236196
rect 580901 232386 580967 232389
rect 583520 232386 584960 232476
rect 580901 232384 584960 232386
rect 580901 232328 580906 232384
rect 580962 232328 584960 232384
rect 580901 232326 584960 232328
rect 580901 232323 580967 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580625 205730 580691 205733
rect 583520 205730 584960 205820
rect 580625 205728 584960 205730
rect 580625 205672 580630 205728
rect 580686 205672 584960 205728
rect 580625 205670 584960 205672
rect 580625 205667 580691 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 580717 192538 580783 192541
rect 583520 192538 584960 192628
rect 580717 192536 584960 192538
rect 580717 192480 580722 192536
rect 580778 192480 584960 192536
rect 580717 192478 584960 192480
rect 580717 192475 580783 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 579613 179210 579679 179213
rect 583520 179210 584960 179300
rect 579613 179208 584960 179210
rect 579613 179152 579618 179208
rect 579674 179152 584960 179208
rect 579613 179150 584960 179152
rect 579613 179147 579679 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580533 165882 580599 165885
rect 583520 165882 584960 165972
rect 580533 165880 584960 165882
rect 580533 165824 580538 165880
rect 580594 165824 584960 165880
rect 580533 165822 584960 165824
rect 580533 165819 580599 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 580441 152690 580507 152693
rect 583520 152690 584960 152780
rect 580441 152688 584960 152690
rect 580441 152632 580446 152688
rect 580502 152632 584960 152688
rect 580441 152630 584960 152632
rect 580441 152627 580507 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 580349 126034 580415 126037
rect 583520 126034 584960 126124
rect 580349 126032 584960 126034
rect 580349 125976 580354 126032
rect 580410 125976 584960 126032
rect 580349 125974 584960 125976
rect 580349 125971 580415 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580257 112842 580323 112845
rect 583520 112842 584960 112932
rect 580257 112840 584960 112842
rect 580257 112784 580262 112840
rect 580318 112784 584960 112840
rect 580257 112782 584960 112784
rect 580257 112779 580323 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 2773 71634 2839 71637
rect -960 71632 2839 71634
rect -960 71576 2778 71632
rect 2834 71576 2839 71632
rect -960 71574 2839 71576
rect -960 71484 480 71574
rect 2773 71571 2839 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 277577 4858 277643 4861
rect 533705 4858 533771 4861
rect 277577 4856 533771 4858
rect 277577 4800 277582 4856
rect 277638 4800 533710 4856
rect 533766 4800 533771 4856
rect 277577 4798 533771 4800
rect 277577 4795 277643 4798
rect 533705 4795 533771 4798
rect 427077 3906 427143 3909
rect 530117 3906 530183 3909
rect 427077 3904 530183 3906
rect 427077 3848 427082 3904
rect 427138 3848 530122 3904
rect 530178 3848 530183 3904
rect 427077 3846 530183 3848
rect 427077 3843 427143 3846
rect 530117 3843 530183 3846
rect 289169 3770 289235 3773
rect 515949 3770 516015 3773
rect 289169 3768 516015 3770
rect 289169 3712 289174 3768
rect 289230 3712 515954 3768
rect 516010 3712 516015 3768
rect 289169 3710 516015 3712
rect 289169 3707 289235 3710
rect 515949 3707 516015 3710
rect 290641 3634 290707 3637
rect 519537 3634 519603 3637
rect 290641 3632 519603 3634
rect 290641 3576 290646 3632
rect 290702 3576 519542 3632
rect 519598 3576 519603 3632
rect 290641 3574 519603 3576
rect 290641 3571 290707 3574
rect 519537 3571 519603 3574
rect 290457 3498 290523 3501
rect 523033 3498 523099 3501
rect 290457 3496 523099 3498
rect 290457 3440 290462 3496
rect 290518 3440 523038 3496
rect 523094 3440 523099 3496
rect 290457 3438 523099 3440
rect 290457 3435 290523 3438
rect 523033 3435 523099 3438
rect 279325 3362 279391 3365
rect 526621 3362 526687 3365
rect 279325 3360 526687 3362
rect 279325 3304 279330 3360
rect 279386 3304 526626 3360
rect 526682 3304 526687 3360
rect 279325 3302 526687 3304
rect 279325 3299 279391 3302
rect 526621 3299 526687 3302
<< via3 >>
rect 238524 337920 238588 337924
rect 238524 337864 238528 337920
rect 238528 337864 238584 337920
rect 238584 337864 238588 337920
rect 238524 337860 238588 337864
rect 239260 337860 239324 337924
rect 238524 337588 238588 337652
rect 245700 337920 245764 337924
rect 245700 337864 245704 337920
rect 245704 337864 245760 337920
rect 245760 337864 245764 337920
rect 245700 337860 245764 337864
rect 245700 337648 245764 337652
rect 245700 337592 245714 337648
rect 245714 337592 245764 337648
rect 245700 337588 245764 337592
rect 268700 337898 268704 337924
rect 268704 337898 268760 337924
rect 268760 337898 268764 337924
rect 268700 337860 268764 337898
rect 272564 337860 272628 337924
rect 278268 337920 278332 337924
rect 278268 337864 278272 337920
rect 278272 337864 278328 337920
rect 278328 337864 278332 337920
rect 278268 337860 278332 337864
rect 272564 335548 272628 335612
rect 239260 334732 239324 334796
rect 278268 334460 278332 334524
rect 268700 333916 268764 333980
rect 468156 322492 468220 322556
rect 469444 322552 469508 322556
rect 469444 322496 469458 322552
rect 469458 322496 469508 322552
rect 469444 322492 469508 322496
rect 474596 322552 474660 322556
rect 474596 322496 474610 322552
rect 474610 322496 474660 322552
rect 474596 322492 474660 322496
rect 476804 322492 476868 322556
rect 479196 322552 479260 322556
rect 479196 322496 479210 322552
rect 479210 322496 479260 322552
rect 479196 322492 479260 322496
rect 481956 322492 482020 322556
rect 483244 322492 483308 322556
rect 485452 322492 485516 322556
rect 489500 322492 489564 322556
rect 490604 322552 490668 322556
rect 490604 322496 490618 322552
rect 490618 322496 490668 322552
rect 490604 322492 490668 322496
rect 492996 322492 493060 322556
rect 519492 322416 519556 322420
rect 519492 322360 519542 322416
rect 519542 322360 519556 322416
rect 519492 322356 519556 322360
rect 486924 321948 486988 322012
rect 470732 321600 470796 321604
rect 470732 321544 470746 321600
rect 470746 321544 470796 321600
rect 470732 321540 470796 321544
rect 472020 321600 472084 321604
rect 472020 321544 472034 321600
rect 472034 321544 472084 321600
rect 472020 321540 472084 321544
rect 473124 321540 473188 321604
rect 475700 321540 475764 321604
rect 478276 321600 478340 321604
rect 478276 321544 478290 321600
rect 478290 321544 478340 321600
rect 478276 321540 478340 321544
rect 480668 321600 480732 321604
rect 480668 321544 480682 321600
rect 480682 321544 480732 321600
rect 480668 321540 480732 321544
rect 484348 321600 484412 321604
rect 484348 321544 484398 321600
rect 484398 321544 484412 321600
rect 484348 321540 484412 321544
rect 492260 321600 492324 321604
rect 492260 321544 492274 321600
rect 492274 321544 492324 321600
rect 492260 321540 492324 321544
rect 494284 321600 494348 321604
rect 494284 321544 494298 321600
rect 494298 321544 494348 321600
rect 494284 321540 494348 321544
rect 496860 321600 496924 321604
rect 496860 321544 496874 321600
rect 496874 321544 496924 321600
rect 496860 321540 496924 321544
rect 498148 321600 498212 321604
rect 498148 321544 498198 321600
rect 498198 321544 498212 321600
rect 498148 321540 498212 321544
rect 500724 321600 500788 321604
rect 500724 321544 500738 321600
rect 500738 321544 500788 321600
rect 500724 321540 500788 321544
rect 501828 321540 501892 321604
rect 503300 321600 503364 321604
rect 503300 321544 503314 321600
rect 503314 321544 503364 321600
rect 503300 321540 503364 321544
rect 504220 321600 504284 321604
rect 504220 321544 504234 321600
rect 504234 321544 504284 321600
rect 504220 321540 504284 321544
rect 505508 321600 505572 321604
rect 505508 321544 505522 321600
rect 505522 321544 505572 321600
rect 505508 321540 505572 321544
rect 506980 321600 507044 321604
rect 506980 321544 506994 321600
rect 506994 321544 507044 321600
rect 506980 321540 507044 321544
rect 529980 321600 530044 321604
rect 529980 321544 530030 321600
rect 530030 321544 530044 321600
rect 529980 321540 530044 321544
rect 488212 321268 488276 321332
rect 495572 321268 495636 321332
rect 499252 321268 499316 321332
rect 445854 239864 445918 239868
rect 445854 239808 445906 239864
rect 445906 239808 445918 239864
rect 445854 239804 445918 239808
rect 469246 239804 469310 239868
rect 522694 239864 522758 239868
rect 522694 239808 522726 239864
rect 522726 239808 522758 239864
rect 522694 239804 522758 239808
rect 522966 239804 523030 239868
rect 473190 239728 473254 239732
rect 473190 239672 473230 239728
rect 473230 239672 473254 239728
rect 473190 239668 473254 239672
rect 475638 239728 475702 239732
rect 475638 239672 475658 239728
rect 475658 239672 475702 239728
rect 475638 239668 475702 239672
rect 523102 239728 523166 239732
rect 523102 239672 523130 239728
rect 523130 239672 523166 239728
rect 523102 239668 523166 239672
rect 471966 239592 472030 239596
rect 471966 239536 471978 239592
rect 471978 239536 472030 239592
rect 471966 239532 472030 239536
rect 473308 239532 473372 239596
rect 474414 239532 474478 239596
rect 479310 239592 479374 239596
rect 479310 239536 479338 239592
rect 479338 239536 479374 239592
rect 479310 239532 479374 239536
rect 487878 239592 487942 239596
rect 487878 239536 487894 239592
rect 487894 239536 487942 239592
rect 487878 239532 487942 239536
rect 492996 239532 493060 239596
rect 493998 239532 494062 239596
rect 495630 239592 495694 239596
rect 495630 239536 495678 239592
rect 495678 239536 495694 239592
rect 495630 239532 495694 239536
rect 496854 239592 496918 239596
rect 496854 239536 496874 239592
rect 496874 239536 496918 239592
rect 496854 239532 496918 239536
rect 500526 239592 500590 239596
rect 500526 239536 500554 239592
rect 500554 239536 500590 239592
rect 500526 239532 500590 239536
rect 501886 239592 501950 239596
rect 501886 239536 501934 239592
rect 501934 239536 501950 239592
rect 501886 239532 501950 239536
rect 503110 239592 503174 239596
rect 503110 239536 503130 239592
rect 503130 239536 503174 239592
rect 503110 239532 503174 239536
rect 505558 239592 505622 239596
rect 505558 239536 505614 239592
rect 505614 239536 505622 239592
rect 505558 239532 505622 239536
rect 506782 239592 506846 239596
rect 506782 239536 506810 239592
rect 506810 239536 506846 239592
rect 506782 239532 506846 239536
rect 455460 239124 455524 239188
rect 457852 238988 457916 239052
rect 456748 238852 456812 238916
rect 459140 238716 459204 238780
rect 477724 238640 477788 238644
rect 477724 238584 477738 238640
rect 477738 238584 477788 238640
rect 477724 238580 477788 238584
rect 481404 238580 481468 238644
rect 483428 238640 483492 238644
rect 483428 238584 483442 238640
rect 483442 238584 483492 238640
rect 483428 238580 483492 238584
rect 484348 238640 484412 238644
rect 484348 238584 484398 238640
rect 484398 238584 484412 238640
rect 484348 238580 484412 238584
rect 485452 238640 485516 238644
rect 485452 238584 485466 238640
rect 485466 238584 485516 238640
rect 485452 238580 485516 238584
rect 478828 238444 478892 238508
rect 482324 238504 482388 238508
rect 482324 238448 482338 238504
rect 482338 238448 482388 238504
rect 482324 238444 482388 238448
rect 484900 238504 484964 238508
rect 484900 238448 484914 238504
rect 484914 238448 484964 238504
rect 484900 238444 484964 238448
rect 474044 238308 474108 238372
rect 476620 238368 476684 238372
rect 476620 238312 476634 238368
rect 476634 238312 476684 238368
rect 476620 238308 476684 238312
rect 480668 238368 480732 238372
rect 480668 238312 480682 238368
rect 480682 238312 480732 238368
rect 480668 238308 480732 238312
rect 481772 238368 481836 238372
rect 481772 238312 481786 238368
rect 481786 238312 481836 238368
rect 481772 238308 481836 238312
rect 486004 238368 486068 238372
rect 486004 238312 486018 238368
rect 486018 238312 486068 238368
rect 486004 238308 486068 238312
rect 488212 238368 488276 238372
rect 488212 238312 488226 238368
rect 488226 238312 488276 238368
rect 488212 238308 488276 238312
rect 490788 238172 490852 238236
rect 491708 238232 491772 238236
rect 491708 238176 491722 238232
rect 491722 238176 491772 238232
rect 491708 238172 491772 238176
rect 492812 238232 492876 238236
rect 492812 238176 492826 238232
rect 492826 238176 492876 238232
rect 492812 238172 492876 238176
rect 495204 238232 495268 238236
rect 495204 238176 495218 238232
rect 495218 238176 495268 238232
rect 495204 238172 495268 238176
rect 497596 237764 497660 237828
rect 467236 237688 467300 237692
rect 467236 237632 467250 237688
rect 467250 237632 467300 237688
rect 467236 237628 467300 237632
rect 467788 237688 467852 237692
rect 467788 237632 467838 237688
rect 467838 237632 467852 237688
rect 467788 237628 467852 237632
rect 462636 237220 462700 237284
rect 463740 237280 463804 237284
rect 463740 237224 463754 237280
rect 463754 237224 463804 237280
rect 463740 237220 463804 237224
rect 466132 237220 466196 237284
rect 468340 237220 468404 237284
rect 469628 237220 469692 237284
rect 470732 237220 470796 237284
rect 487108 237220 487172 237284
rect 498700 237220 498764 237284
rect 504220 237220 504284 237284
rect 522804 237220 522868 237284
rect 483060 237084 483124 237148
rect 490604 237084 490668 237148
rect 493180 237084 493244 237148
rect 494284 237084 494348 237148
rect 480300 236948 480364 237012
rect 491340 237008 491404 237012
rect 491340 236952 491354 237008
rect 491354 236952 491404 237008
rect 491340 236948 491404 236952
rect 460060 236812 460124 236876
rect 461348 236812 461412 236876
rect 465028 236872 465092 236876
rect 465028 236816 465078 236872
rect 465078 236816 465092 236872
rect 465028 236812 465092 236816
rect 472940 236812 473004 236876
rect 473308 236872 473372 236876
rect 473308 236816 473358 236872
rect 473358 236816 473372 236872
rect 473308 236812 473372 236816
rect 475332 236812 475396 236876
rect 476804 236812 476868 236876
rect 486556 236812 486620 236876
rect 489316 236812 489380 236876
rect 492996 236676 493060 236740
rect 497780 236540 497844 236604
rect 489132 236404 489196 236468
rect 471836 236268 471900 236332
rect 469260 236192 469324 236196
rect 469260 236136 469274 236192
rect 469274 236136 469324 236192
rect 469260 236132 469324 236136
rect 478092 236132 478156 236196
rect 496492 236132 496556 236196
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 390000 236414 416898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 390000 240134 420618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 390000 243854 424338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 390000 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 390000 254414 398898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 390000 258134 402618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 390000 261854 406338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 390000 265574 410058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 390000 272414 416898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 390000 276134 420618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 390000 279854 424338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 390000 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 254568 381454 254888 381486
rect 254568 381218 254610 381454
rect 254846 381218 254888 381454
rect 254568 381134 254888 381218
rect 254568 380898 254610 381134
rect 254846 380898 254888 381134
rect 254568 380866 254888 380898
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 239208 363454 239528 363486
rect 239208 363218 239250 363454
rect 239486 363218 239528 363454
rect 239208 363134 239528 363218
rect 239208 362898 239250 363134
rect 239486 362898 239528 363134
rect 239208 362866 239528 362898
rect 269928 363454 270248 363486
rect 269928 363218 269970 363454
rect 270206 363218 270248 363454
rect 269928 363134 270248 363218
rect 269928 362898 269970 363134
rect 270206 362898 270248 363134
rect 269928 362866 270248 362898
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 254568 345454 254888 345486
rect 254568 345218 254610 345454
rect 254846 345218 254888 345454
rect 254568 345134 254888 345218
rect 254568 344898 254610 345134
rect 254846 344898 254888 345134
rect 254568 344866 254888 344898
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 238523 337924 238589 337925
rect 238523 337860 238524 337924
rect 238588 337860 238589 337924
rect 238523 337859 238589 337860
rect 239259 337924 239325 337925
rect 239259 337860 239260 337924
rect 239324 337860 239325 337924
rect 239259 337859 239325 337860
rect 245699 337924 245765 337925
rect 245699 337860 245700 337924
rect 245764 337860 245765 337924
rect 245699 337859 245765 337860
rect 268699 337924 268765 337925
rect 268699 337860 268700 337924
rect 268764 337860 268765 337924
rect 268699 337859 268765 337860
rect 272563 337924 272629 337925
rect 272563 337860 272564 337924
rect 272628 337860 272629 337924
rect 272563 337859 272629 337860
rect 278267 337924 278333 337925
rect 278267 337860 278268 337924
rect 278332 337860 278333 337924
rect 278267 337859 278333 337860
rect 238526 337653 238586 337859
rect 238523 337652 238589 337653
rect 238523 337588 238524 337652
rect 238588 337588 238589 337652
rect 238523 337587 238589 337588
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 309454 236414 336000
rect 239262 334797 239322 337859
rect 245702 337653 245762 337859
rect 245699 337652 245765 337653
rect 245699 337588 245700 337652
rect 245764 337588 245765 337652
rect 245699 337587 245765 337588
rect 239259 334796 239325 334797
rect 239259 334732 239260 334796
rect 239324 334732 239325 334796
rect 239259 334731 239325 334732
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 313174 240134 336000
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 277174 240134 312618
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 316894 243854 336000
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 320614 247574 336000
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 327454 254414 336000
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 331174 258134 336000
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 334894 261854 336000
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 302614 265574 336000
rect 268702 333981 268762 337859
rect 268699 333980 268765 333981
rect 268699 333916 268700 333980
rect 268764 333916 268765 333980
rect 268699 333915 268765 333916
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 309454 272414 336000
rect 272566 335613 272626 337859
rect 272563 335612 272629 335613
rect 272563 335548 272564 335612
rect 272628 335548 272629 335612
rect 272563 335547 272629 335548
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 313174 276134 336000
rect 278270 334525 278330 337859
rect 278267 334524 278333 334525
rect 278267 334460 278268 334524
rect 278332 334460 278333 334524
rect 278267 334459 278333 334460
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 316894 279854 336000
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 320614 283574 336000
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 321500 438134 330618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 321500 441854 334338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 321500 445574 338058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 321500 452414 344898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 321500 456134 348618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 321500 459854 352338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 321500 463574 356058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 468155 322556 468221 322557
rect 468155 322492 468156 322556
rect 468220 322492 468221 322556
rect 468155 322491 468221 322492
rect 469443 322556 469509 322557
rect 469443 322492 469444 322556
rect 469508 322492 469509 322556
rect 469443 322491 469509 322492
rect 468158 319970 468218 322491
rect 469446 319970 469506 322491
rect 469794 321500 470414 326898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 470731 321604 470797 321605
rect 470731 321540 470732 321604
rect 470796 321540 470797 321604
rect 470731 321539 470797 321540
rect 472019 321604 472085 321605
rect 472019 321540 472020 321604
rect 472084 321540 472085 321604
rect 472019 321539 472085 321540
rect 473123 321604 473189 321605
rect 473123 321540 473124 321604
rect 473188 321540 473189 321604
rect 473123 321539 473189 321540
rect 470734 319970 470794 321539
rect 472022 319970 472082 321539
rect 468158 319910 468220 319970
rect 469446 319910 469580 319970
rect 468160 319394 468220 319910
rect 469520 319394 469580 319910
rect 470608 319910 470794 319970
rect 471968 319910 472082 319970
rect 473126 319970 473186 321539
rect 473514 321500 474134 330618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 474595 322556 474661 322557
rect 474595 322492 474596 322556
rect 474660 322492 474661 322556
rect 474595 322491 474661 322492
rect 476803 322556 476869 322557
rect 476803 322492 476804 322556
rect 476868 322492 476869 322556
rect 476803 322491 476869 322492
rect 474598 319970 474658 322491
rect 475699 321604 475765 321605
rect 475699 321540 475700 321604
rect 475764 321540 475765 321604
rect 475699 321539 475765 321540
rect 473126 319910 473252 319970
rect 470608 319394 470668 319910
rect 471968 319394 472028 319910
rect 473192 319394 473252 319910
rect 474552 319910 474658 319970
rect 475702 319970 475762 321539
rect 476806 319970 476866 322491
rect 477234 321500 477854 334338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 479195 322556 479261 322557
rect 479195 322492 479196 322556
rect 479260 322492 479261 322556
rect 479195 322491 479261 322492
rect 478275 321604 478341 321605
rect 478275 321540 478276 321604
rect 478340 321540 478341 321604
rect 478275 321539 478341 321540
rect 478278 319970 478338 321539
rect 475702 319910 475836 319970
rect 476806 319910 476924 319970
rect 474552 319394 474612 319910
rect 475776 319394 475836 319910
rect 476864 319394 476924 319910
rect 478224 319910 478338 319970
rect 479198 319970 479258 322491
rect 480667 321604 480733 321605
rect 480667 321540 480668 321604
rect 480732 321540 480733 321604
rect 480667 321539 480733 321540
rect 480670 319970 480730 321539
rect 480954 321500 481574 338058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 481955 322556 482021 322557
rect 481955 322492 481956 322556
rect 482020 322492 482021 322556
rect 481955 322491 482021 322492
rect 483243 322556 483309 322557
rect 483243 322492 483244 322556
rect 483308 322492 483309 322556
rect 483243 322491 483309 322492
rect 485451 322556 485517 322557
rect 485451 322492 485452 322556
rect 485516 322492 485517 322556
rect 485451 322491 485517 322492
rect 481958 319970 482018 322491
rect 479198 319910 479372 319970
rect 480670 319910 480732 319970
rect 478224 319394 478284 319910
rect 479312 319394 479372 319910
rect 480672 319394 480732 319910
rect 481896 319910 482018 319970
rect 483246 319970 483306 322491
rect 484347 321604 484413 321605
rect 484347 321540 484348 321604
rect 484412 321540 484413 321604
rect 484347 321539 484413 321540
rect 484350 319970 484410 321539
rect 483246 319910 483316 319970
rect 481896 319394 481956 319910
rect 483256 319394 483316 319910
rect 484344 319910 484410 319970
rect 485454 319970 485514 322491
rect 486923 322012 486989 322013
rect 486923 321948 486924 322012
rect 486988 321948 486989 322012
rect 486923 321947 486989 321948
rect 486926 319970 486986 321947
rect 487794 321500 488414 344898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 489499 322556 489565 322557
rect 489499 322492 489500 322556
rect 489564 322492 489565 322556
rect 489499 322491 489565 322492
rect 490603 322556 490669 322557
rect 490603 322492 490604 322556
rect 490668 322492 490669 322556
rect 490603 322491 490669 322492
rect 488211 321332 488277 321333
rect 488211 321268 488212 321332
rect 488276 321268 488277 321332
rect 488211 321267 488277 321268
rect 488214 319970 488274 321267
rect 485454 319910 485628 319970
rect 486926 319910 486988 319970
rect 484344 319394 484404 319910
rect 485568 319394 485628 319910
rect 486928 319394 486988 319910
rect 488152 319910 488274 319970
rect 489502 319970 489562 322491
rect 490606 319970 490666 322491
rect 491514 321500 492134 348618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 492995 322556 493061 322557
rect 492995 322492 492996 322556
rect 493060 322492 493061 322556
rect 492995 322491 493061 322492
rect 492259 321604 492325 321605
rect 492259 321540 492260 321604
rect 492324 321540 492325 321604
rect 492259 321539 492325 321540
rect 492262 319970 492322 321539
rect 489502 319910 489572 319970
rect 488152 319394 488212 319910
rect 489512 319394 489572 319910
rect 490600 319910 490666 319970
rect 491960 319910 492322 319970
rect 492998 319970 493058 322491
rect 494283 321604 494349 321605
rect 494283 321540 494284 321604
rect 494348 321540 494349 321604
rect 494283 321539 494349 321540
rect 494286 319970 494346 321539
rect 495234 321500 495854 352338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 496859 321604 496925 321605
rect 496859 321540 496860 321604
rect 496924 321540 496925 321604
rect 496859 321539 496925 321540
rect 498147 321604 498213 321605
rect 498147 321540 498148 321604
rect 498212 321540 498213 321604
rect 498147 321539 498213 321540
rect 495571 321332 495637 321333
rect 495571 321268 495572 321332
rect 495636 321268 495637 321332
rect 495571 321267 495637 321268
rect 492998 319910 493108 319970
rect 490600 319394 490660 319910
rect 491960 319394 492020 319910
rect 493048 319394 493108 319910
rect 494272 319910 494346 319970
rect 495574 319970 495634 321267
rect 496862 319970 496922 321539
rect 495574 319910 495692 319970
rect 494272 319394 494332 319910
rect 495632 319394 495692 319910
rect 496856 319910 496922 319970
rect 498150 319970 498210 321539
rect 498954 321500 499574 356058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 500723 321604 500789 321605
rect 500723 321540 500724 321604
rect 500788 321540 500789 321604
rect 500723 321539 500789 321540
rect 501827 321604 501893 321605
rect 501827 321540 501828 321604
rect 501892 321540 501893 321604
rect 501827 321539 501893 321540
rect 503299 321604 503365 321605
rect 503299 321540 503300 321604
rect 503364 321540 503365 321604
rect 503299 321539 503365 321540
rect 504219 321604 504285 321605
rect 504219 321540 504220 321604
rect 504284 321540 504285 321604
rect 504219 321539 504285 321540
rect 505507 321604 505573 321605
rect 505507 321540 505508 321604
rect 505572 321540 505573 321604
rect 505507 321539 505573 321540
rect 499251 321332 499317 321333
rect 499251 321268 499252 321332
rect 499316 321268 499317 321332
rect 499251 321267 499317 321268
rect 499254 319970 499314 321267
rect 500726 319970 500786 321539
rect 498150 319910 498276 319970
rect 499254 319910 499364 319970
rect 496856 319394 496916 319910
rect 498216 319394 498276 319910
rect 499304 319394 499364 319910
rect 500664 319910 500786 319970
rect 501830 319970 501890 321539
rect 503302 319970 503362 321539
rect 501830 319910 501948 319970
rect 500664 319394 500724 319910
rect 501888 319394 501948 319910
rect 503248 319910 503362 319970
rect 504222 319970 504282 321539
rect 505510 319970 505570 321539
rect 505794 321500 506414 326898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 506979 321604 507045 321605
rect 506979 321540 506980 321604
rect 507044 321540 507045 321604
rect 506979 321539 507045 321540
rect 506982 319970 507042 321539
rect 509514 321500 510134 330618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 321500 513854 334338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 321500 517574 338058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 519491 322420 519557 322421
rect 519491 322356 519492 322420
rect 519556 322356 519557 322420
rect 519491 322355 519557 322356
rect 519494 319970 519554 322355
rect 523794 321500 524414 344898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 321500 528134 348618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 529979 321604 530045 321605
rect 529979 321540 529980 321604
rect 530044 321540 530045 321604
rect 529979 321539 530045 321540
rect 504222 319910 504396 319970
rect 505510 319910 505620 319970
rect 503248 319394 503308 319910
rect 504336 319394 504396 319910
rect 505560 319394 505620 319910
rect 506920 319910 507042 319970
rect 519432 319910 519554 319970
rect 529982 319970 530042 321539
rect 531234 321500 531854 352338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 321500 535574 356058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 529982 319910 530100 319970
rect 506920 319394 506980 319910
rect 519432 319394 519492 319910
rect 530040 319394 530100 319910
rect 440272 309454 440620 309486
rect 440272 309218 440328 309454
rect 440564 309218 440620 309454
rect 440272 309134 440620 309218
rect 440272 308898 440328 309134
rect 440564 308898 440620 309134
rect 440272 308866 440620 308898
rect 535336 309454 535684 309486
rect 535336 309218 535392 309454
rect 535628 309218 535684 309454
rect 535336 309134 535684 309218
rect 535336 308898 535392 309134
rect 535628 308898 535684 309134
rect 535336 308866 535684 308898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 440952 291454 441300 291486
rect 440952 291218 441008 291454
rect 441244 291218 441300 291454
rect 440952 291134 441300 291218
rect 440952 290898 441008 291134
rect 441244 290898 441300 291134
rect 440952 290866 441300 290898
rect 534656 291454 535004 291486
rect 534656 291218 534712 291454
rect 534948 291218 535004 291454
rect 534656 291134 535004 291218
rect 534656 290898 534712 291134
rect 534948 290898 535004 291134
rect 534656 290866 535004 290898
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 440272 273454 440620 273486
rect 440272 273218 440328 273454
rect 440564 273218 440620 273454
rect 440272 273134 440620 273218
rect 440272 272898 440328 273134
rect 440564 272898 440620 273134
rect 440272 272866 440620 272898
rect 535336 273454 535684 273486
rect 535336 273218 535392 273454
rect 535628 273218 535684 273454
rect 535336 273134 535684 273218
rect 535336 272898 535392 273134
rect 535628 272898 535684 273134
rect 535336 272866 535684 272898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 440952 255454 441300 255486
rect 440952 255218 441008 255454
rect 441244 255218 441300 255454
rect 440952 255134 441300 255218
rect 440952 254898 441008 255134
rect 441244 254898 441300 255134
rect 440952 254866 441300 254898
rect 534656 255454 535004 255486
rect 534656 255218 534712 255454
rect 534948 255218 535004 255454
rect 534656 255134 535004 255218
rect 534656 254898 534712 255134
rect 534948 254898 535004 255134
rect 534656 254866 535004 254898
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 445856 239869 445916 240040
rect 445853 239868 445919 239869
rect 445853 239804 445854 239868
rect 445918 239804 445919 239868
rect 445853 239803 445919 239804
rect 455512 239730 455572 240040
rect 455462 239670 455572 239730
rect 456736 239730 456796 240040
rect 457824 239730 457884 240040
rect 459184 239730 459244 240040
rect 460136 239730 460196 240040
rect 461360 239730 461420 240040
rect 456736 239670 456810 239730
rect 457824 239670 457914 239730
rect 455462 239189 455522 239670
rect 455459 239188 455525 239189
rect 455459 239124 455460 239188
rect 455524 239124 455525 239188
rect 455459 239123 455525 239124
rect 456750 238917 456810 239670
rect 457854 239053 457914 239670
rect 459142 239670 459244 239730
rect 460062 239670 460196 239730
rect 461350 239670 461420 239730
rect 462584 239730 462644 240040
rect 463672 239730 463732 240040
rect 465032 239730 465092 240040
rect 462584 239670 462698 239730
rect 463672 239670 463802 239730
rect 457851 239052 457917 239053
rect 457851 238988 457852 239052
rect 457916 238988 457917 239052
rect 457851 238987 457917 238988
rect 456747 238916 456813 238917
rect 456747 238852 456748 238916
rect 456812 238852 456813 238916
rect 456747 238851 456813 238852
rect 459142 238781 459202 239670
rect 459139 238780 459205 238781
rect 459139 238716 459140 238780
rect 459204 238716 459205 238780
rect 459139 238715 459205 238716
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 223174 438134 238000
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 226894 441854 238000
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 230614 445574 238000
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 237454 452414 238000
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 205174 456134 238000
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 208894 459854 238000
rect 460062 236877 460122 239670
rect 461350 236877 461410 239670
rect 462638 237285 462698 239670
rect 462635 237284 462701 237285
rect 462635 237220 462636 237284
rect 462700 237220 462701 237284
rect 462635 237219 462701 237220
rect 460059 236876 460125 236877
rect 460059 236812 460060 236876
rect 460124 236812 460125 236876
rect 460059 236811 460125 236812
rect 461347 236876 461413 236877
rect 461347 236812 461348 236876
rect 461412 236812 461413 236876
rect 461347 236811 461413 236812
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 212614 463574 238000
rect 463742 237285 463802 239670
rect 465030 239670 465092 239730
rect 466120 239730 466180 240040
rect 467208 239730 467268 240040
rect 467888 239730 467948 240040
rect 466120 239670 466194 239730
rect 467208 239670 467298 239730
rect 463739 237284 463805 237285
rect 463739 237220 463740 237284
rect 463804 237220 463805 237284
rect 463739 237219 463805 237220
rect 465030 236877 465090 239670
rect 466134 237285 466194 239670
rect 467238 237693 467298 239670
rect 467790 239670 467948 239730
rect 468296 239730 468356 240040
rect 469248 239869 469308 240040
rect 469245 239868 469311 239869
rect 469245 239804 469246 239868
rect 469310 239804 469311 239868
rect 469245 239803 469311 239804
rect 469656 239730 469716 240040
rect 470336 239730 470396 240040
rect 470744 239730 470804 240040
rect 468296 239670 468402 239730
rect 467790 237693 467850 239670
rect 467235 237692 467301 237693
rect 467235 237628 467236 237692
rect 467300 237628 467301 237692
rect 467235 237627 467301 237628
rect 467787 237692 467853 237693
rect 467787 237628 467788 237692
rect 467852 237628 467853 237692
rect 467787 237627 467853 237628
rect 468342 237285 468402 239670
rect 469262 239670 469716 239730
rect 469814 239670 470396 239730
rect 470734 239670 470804 239730
rect 471832 239730 471892 240040
rect 471832 239670 471898 239730
rect 466131 237284 466197 237285
rect 466131 237220 466132 237284
rect 466196 237220 466197 237284
rect 466131 237219 466197 237220
rect 468339 237284 468405 237285
rect 468339 237220 468340 237284
rect 468404 237220 468405 237284
rect 468339 237219 468405 237220
rect 465027 236876 465093 236877
rect 465027 236812 465028 236876
rect 465092 236812 465093 236876
rect 465027 236811 465093 236812
rect 469262 236197 469322 239670
rect 469814 238370 469874 239670
rect 469630 238310 469874 238370
rect 469630 237285 469690 238310
rect 469627 237284 469693 237285
rect 469627 237220 469628 237284
rect 469692 237220 469693 237284
rect 469627 237219 469693 237220
rect 469259 236196 469325 236197
rect 469259 236132 469260 236196
rect 469324 236132 469325 236196
rect 469259 236131 469325 236132
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 219454 470414 238000
rect 470734 237285 470794 239670
rect 470731 237284 470797 237285
rect 470731 237220 470732 237284
rect 470796 237220 470797 237284
rect 470731 237219 470797 237220
rect 471838 236333 471898 239670
rect 471968 239597 472028 240040
rect 473056 239730 473116 240040
rect 473192 239733 473252 240040
rect 472942 239670 473116 239730
rect 473189 239732 473255 239733
rect 471965 239596 472031 239597
rect 471965 239532 471966 239596
rect 472030 239532 472031 239596
rect 471965 239531 472031 239532
rect 472942 236877 473002 239670
rect 473189 239668 473190 239732
rect 473254 239668 473255 239732
rect 474144 239730 474204 240040
rect 473189 239667 473255 239668
rect 474046 239670 474204 239730
rect 473307 239596 473373 239597
rect 473307 239532 473308 239596
rect 473372 239532 473373 239596
rect 473307 239531 473373 239532
rect 473310 236877 473370 239531
rect 474046 238373 474106 239670
rect 474416 239597 474476 240040
rect 475504 239730 475564 240040
rect 475640 239733 475700 240040
rect 475334 239670 475564 239730
rect 475637 239732 475703 239733
rect 474413 239596 474479 239597
rect 474413 239532 474414 239596
rect 474478 239532 474479 239596
rect 474413 239531 474479 239532
rect 474043 238372 474109 238373
rect 474043 238308 474044 238372
rect 474108 238308 474109 238372
rect 474043 238307 474109 238308
rect 472939 236876 473005 236877
rect 472939 236812 472940 236876
rect 473004 236812 473005 236876
rect 472939 236811 473005 236812
rect 473307 236876 473373 236877
rect 473307 236812 473308 236876
rect 473372 236812 473373 236876
rect 473307 236811 473373 236812
rect 471835 236332 471901 236333
rect 471835 236268 471836 236332
rect 471900 236268 471901 236332
rect 471835 236267 471901 236268
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 223174 474134 238000
rect 475334 236877 475394 239670
rect 475637 239668 475638 239732
rect 475702 239668 475703 239732
rect 476592 239730 476652 240040
rect 476864 239730 476924 240040
rect 476592 239670 476682 239730
rect 475637 239667 475703 239668
rect 476622 238373 476682 239670
rect 476806 239670 476924 239730
rect 476619 238372 476685 238373
rect 476619 238308 476620 238372
rect 476684 238308 476685 238372
rect 476619 238307 476685 238308
rect 476806 236877 476866 239670
rect 477680 239050 477740 240040
rect 477816 239730 477876 240040
rect 478904 239730 478964 240040
rect 477816 239670 478154 239730
rect 477680 238990 477786 239050
rect 477726 238645 477786 238990
rect 477723 238644 477789 238645
rect 477723 238580 477724 238644
rect 477788 238580 477789 238644
rect 477723 238579 477789 238580
rect 475331 236876 475397 236877
rect 475331 236812 475332 236876
rect 475396 236812 475397 236876
rect 475331 236811 475397 236812
rect 476803 236876 476869 236877
rect 476803 236812 476804 236876
rect 476868 236812 476869 236876
rect 476803 236811 476869 236812
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 226894 477854 238000
rect 478094 236197 478154 239670
rect 478830 239670 478964 239730
rect 478830 238509 478890 239670
rect 479312 239597 479372 240040
rect 480264 239730 480324 240040
rect 480672 239730 480732 240040
rect 480264 239670 480362 239730
rect 479309 239596 479375 239597
rect 479309 239532 479310 239596
rect 479374 239532 479375 239596
rect 479309 239531 479375 239532
rect 478827 238508 478893 238509
rect 478827 238444 478828 238508
rect 478892 238444 478893 238508
rect 478827 238443 478893 238444
rect 480302 237013 480362 239670
rect 480670 239670 480732 239730
rect 481352 239730 481412 240040
rect 481896 239730 481956 240040
rect 482440 239730 482500 240040
rect 483120 239730 483180 240040
rect 483528 239730 483588 240040
rect 481352 239670 481466 239730
rect 480670 238373 480730 239670
rect 481406 238645 481466 239670
rect 481774 239670 481956 239730
rect 482326 239670 482500 239730
rect 483062 239670 483180 239730
rect 483430 239670 483588 239730
rect 484344 239730 484404 240040
rect 484888 239730 484948 240040
rect 485568 239730 485628 240040
rect 484344 239670 484410 239730
rect 484888 239670 484962 239730
rect 481403 238644 481469 238645
rect 481403 238580 481404 238644
rect 481468 238580 481469 238644
rect 481403 238579 481469 238580
rect 481774 238373 481834 239670
rect 482326 238509 482386 239670
rect 482323 238508 482389 238509
rect 482323 238444 482324 238508
rect 482388 238444 482389 238508
rect 482323 238443 482389 238444
rect 480667 238372 480733 238373
rect 480667 238308 480668 238372
rect 480732 238308 480733 238372
rect 480667 238307 480733 238308
rect 481771 238372 481837 238373
rect 481771 238308 481772 238372
rect 481836 238308 481837 238372
rect 481771 238307 481837 238308
rect 480299 237012 480365 237013
rect 480299 236948 480300 237012
rect 480364 236948 480365 237012
rect 480299 236947 480365 236948
rect 478091 236196 478157 236197
rect 478091 236132 478092 236196
rect 478156 236132 478157 236196
rect 478091 236131 478157 236132
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 230614 481574 238000
rect 483062 237149 483122 239670
rect 483430 238645 483490 239670
rect 484350 238645 484410 239670
rect 483427 238644 483493 238645
rect 483427 238580 483428 238644
rect 483492 238580 483493 238644
rect 483427 238579 483493 238580
rect 484347 238644 484413 238645
rect 484347 238580 484348 238644
rect 484412 238580 484413 238644
rect 484347 238579 484413 238580
rect 484902 238509 484962 239670
rect 485454 239670 485628 239730
rect 485976 239730 486036 240040
rect 486656 239730 486716 240040
rect 485976 239670 486066 239730
rect 485454 238645 485514 239670
rect 485451 238644 485517 238645
rect 485451 238580 485452 238644
rect 485516 238580 485517 238644
rect 485451 238579 485517 238580
rect 484899 238508 484965 238509
rect 484899 238444 484900 238508
rect 484964 238444 484965 238508
rect 484899 238443 484965 238444
rect 486006 238373 486066 239670
rect 486558 239670 486716 239730
rect 487064 239730 487124 240040
rect 487064 239670 487170 239730
rect 486003 238372 486069 238373
rect 486003 238308 486004 238372
rect 486068 238308 486069 238372
rect 486003 238307 486069 238308
rect 483059 237148 483125 237149
rect 483059 237084 483060 237148
rect 483124 237084 483125 237148
rect 483059 237083 483125 237084
rect 486558 236877 486618 239670
rect 487110 237285 487170 239670
rect 487880 239597 487940 240040
rect 488288 239730 488348 240040
rect 488214 239670 488348 239730
rect 489104 239730 489164 240040
rect 489376 239730 489436 240040
rect 489104 239670 489194 239730
rect 487877 239596 487943 239597
rect 487877 239532 487878 239596
rect 487942 239532 487943 239596
rect 487877 239531 487943 239532
rect 488214 238373 488274 239670
rect 488211 238372 488277 238373
rect 488211 238308 488212 238372
rect 488276 238308 488277 238372
rect 488211 238307 488277 238308
rect 487794 237454 488414 238000
rect 487107 237284 487173 237285
rect 487107 237220 487108 237284
rect 487172 237220 487173 237284
rect 487107 237219 487173 237220
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 486555 236876 486621 236877
rect 486555 236812 486556 236876
rect 486620 236812 486621 236876
rect 486555 236811 486621 236812
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 201454 488414 236898
rect 489134 236469 489194 239670
rect 489318 239670 489436 239730
rect 490600 239730 490660 240040
rect 490736 239730 490796 240040
rect 491416 239730 491476 240040
rect 491824 239730 491884 240040
rect 492912 239730 492972 240040
rect 493184 239730 493244 240040
rect 490600 239670 490666 239730
rect 490736 239670 490850 239730
rect 489318 236877 489378 239670
rect 490606 237149 490666 239670
rect 490790 238237 490850 239670
rect 491342 239670 491476 239730
rect 491710 239670 491884 239730
rect 492814 239670 492972 239730
rect 493182 239670 493244 239730
rect 490787 238236 490853 238237
rect 490787 238172 490788 238236
rect 490852 238172 490853 238236
rect 490787 238171 490853 238172
rect 490603 237148 490669 237149
rect 490603 237084 490604 237148
rect 490668 237084 490669 237148
rect 490603 237083 490669 237084
rect 491342 237013 491402 239670
rect 491710 238237 491770 239670
rect 492814 238237 492874 239670
rect 492995 239596 493061 239597
rect 492995 239532 492996 239596
rect 493060 239532 493061 239596
rect 492995 239531 493061 239532
rect 491707 238236 491773 238237
rect 491707 238172 491708 238236
rect 491772 238172 491773 238236
rect 491707 238171 491773 238172
rect 492811 238236 492877 238237
rect 492811 238172 492812 238236
rect 492876 238172 492877 238236
rect 492811 238171 492877 238172
rect 491339 237012 491405 237013
rect 491339 236948 491340 237012
rect 491404 236948 491405 237012
rect 491339 236947 491405 236948
rect 489315 236876 489381 236877
rect 489315 236812 489316 236876
rect 489380 236812 489381 236876
rect 489315 236811 489381 236812
rect 489131 236468 489197 236469
rect 489131 236404 489132 236468
rect 489196 236404 489197 236468
rect 489131 236403 489197 236404
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 205174 492134 238000
rect 492998 236741 493058 239531
rect 493182 237149 493242 239670
rect 494000 239597 494060 240040
rect 494408 239730 494468 240040
rect 495224 239730 495284 240040
rect 494286 239670 494468 239730
rect 495206 239670 495284 239730
rect 493997 239596 494063 239597
rect 493997 239532 493998 239596
rect 494062 239532 494063 239596
rect 493997 239531 494063 239532
rect 494286 237149 494346 239670
rect 495206 238237 495266 239670
rect 495632 239597 495692 240040
rect 496584 239730 496644 240040
rect 496494 239670 496644 239730
rect 495629 239596 495695 239597
rect 495629 239532 495630 239596
rect 495694 239532 495695 239596
rect 495629 239531 495695 239532
rect 495203 238236 495269 238237
rect 495203 238172 495204 238236
rect 495268 238172 495269 238236
rect 495203 238171 495269 238172
rect 493179 237148 493245 237149
rect 493179 237084 493180 237148
rect 493244 237084 493245 237148
rect 493179 237083 493245 237084
rect 494283 237148 494349 237149
rect 494283 237084 494284 237148
rect 494348 237084 494349 237148
rect 494283 237083 494349 237084
rect 492995 236740 493061 236741
rect 492995 236676 492996 236740
rect 493060 236676 493061 236740
rect 492995 236675 493061 236676
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 208894 495854 238000
rect 496494 236197 496554 239670
rect 496856 239597 496916 240040
rect 497672 239730 497732 240040
rect 497598 239670 497732 239730
rect 496853 239596 496919 239597
rect 496853 239532 496854 239596
rect 496918 239532 496919 239596
rect 496853 239531 496919 239532
rect 497598 237829 497658 239670
rect 497808 239050 497868 240040
rect 499304 239730 499364 240040
rect 497782 238990 497868 239050
rect 498702 239670 499364 239730
rect 497595 237828 497661 237829
rect 497595 237764 497596 237828
rect 497660 237764 497661 237828
rect 497595 237763 497661 237764
rect 497782 236605 497842 238990
rect 498702 237285 498762 239670
rect 500528 239597 500588 240040
rect 501888 239597 501948 240040
rect 503112 239597 503172 240040
rect 504336 239730 504396 240040
rect 504222 239670 504396 239730
rect 500525 239596 500591 239597
rect 500525 239532 500526 239596
rect 500590 239532 500591 239596
rect 500525 239531 500591 239532
rect 501885 239596 501951 239597
rect 501885 239532 501886 239596
rect 501950 239532 501951 239596
rect 501885 239531 501951 239532
rect 503109 239596 503175 239597
rect 503109 239532 503110 239596
rect 503174 239532 503175 239596
rect 503109 239531 503175 239532
rect 498699 237284 498765 237285
rect 498699 237220 498700 237284
rect 498764 237220 498765 237284
rect 498699 237219 498765 237220
rect 497779 236604 497845 236605
rect 497779 236540 497780 236604
rect 497844 236540 497845 236604
rect 497779 236539 497845 236540
rect 496491 236196 496557 236197
rect 496491 236132 496492 236196
rect 496556 236132 496557 236196
rect 496491 236131 496557 236132
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 212614 499574 238000
rect 504222 237285 504282 239670
rect 505560 239597 505620 240040
rect 506784 239597 506844 240040
rect 522696 239869 522756 240040
rect 522693 239868 522759 239869
rect 522693 239804 522694 239868
rect 522758 239804 522759 239868
rect 522693 239803 522759 239804
rect 522832 239730 522892 240040
rect 522968 239869 523028 240040
rect 522965 239868 523031 239869
rect 522965 239804 522966 239868
rect 523030 239804 523031 239868
rect 522965 239803 523031 239804
rect 523104 239733 523164 240040
rect 522806 239670 522892 239730
rect 523101 239732 523167 239733
rect 505557 239596 505623 239597
rect 505557 239532 505558 239596
rect 505622 239532 505623 239596
rect 505557 239531 505623 239532
rect 506781 239596 506847 239597
rect 506781 239532 506782 239596
rect 506846 239532 506847 239596
rect 506781 239531 506847 239532
rect 504219 237284 504285 237285
rect 504219 237220 504220 237284
rect 504284 237220 504285 237284
rect 504219 237219 504285 237220
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 219454 506414 238000
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 223174 510134 238000
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 226894 513854 238000
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 230614 517574 238000
rect 522806 237285 522866 239670
rect 523101 239668 523102 239732
rect 523166 239668 523167 239732
rect 523101 239667 523167 239668
rect 523794 237454 524414 238000
rect 522803 237284 522869 237285
rect 522803 237220 522804 237284
rect 522868 237220 522869 237284
rect 522803 237219 522869 237220
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 205174 528134 238000
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 208894 531854 238000
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 212614 535574 238000
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 254610 381218 254846 381454
rect 254610 380898 254846 381134
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 239250 363218 239486 363454
rect 239250 362898 239486 363134
rect 269970 363218 270206 363454
rect 269970 362898 270206 363134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 254610 345218 254846 345454
rect 254610 344898 254846 345134
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 440328 309218 440564 309454
rect 440328 308898 440564 309134
rect 535392 309218 535628 309454
rect 535392 308898 535628 309134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 441008 291218 441244 291454
rect 441008 290898 441244 291134
rect 534712 291218 534948 291454
rect 534712 290898 534948 291134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 440328 273218 440564 273454
rect 440328 272898 440564 273134
rect 535392 273218 535628 273454
rect 535392 272898 535628 273134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 441008 255218 441244 255454
rect 441008 254898 441244 255134
rect 534712 255218 534948 255454
rect 534712 254898 534948 255134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 254610 381454
rect 254846 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 254610 381134
rect 254846 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 239250 363454
rect 239486 363218 269970 363454
rect 270206 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 239250 363134
rect 239486 362898 269970 363134
rect 270206 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 254610 345454
rect 254846 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 254610 345134
rect 254846 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 440328 309454
rect 440564 309218 535392 309454
rect 535628 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 440328 309134
rect 440564 308898 535392 309134
rect 535628 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 441008 291454
rect 441244 291218 534712 291454
rect 534948 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 441008 291134
rect 441244 290898 534712 291134
rect 534948 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 440328 273454
rect 440564 273218 535392 273454
rect 535628 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 440328 273134
rect 440564 272898 535392 273134
rect 535628 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 441008 255454
rect 441244 255218 534712 255454
rect 534948 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 441008 255134
rect 441244 254898 534712 255134
rect 534948 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 1636669832
transform 1 0 235000 0 1 338000
box 0 0 50000 50000
use sky130_sram_1kbyte_1rw1r_32x256_8  SRAM0
timestamp 1636669832
transform 1 0 440000 0 1 240000
box 0 0 95956 79500
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 336000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 390000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 321500 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 321500 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 336000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 390000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 321500 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 321500 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 321500 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 336000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 390000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 321500 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 321500 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 321500 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 336000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 390000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 321500 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 321500 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 321500 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 336000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 336000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 390000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 390000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 321500 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 321500 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 321500 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 336000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 336000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 390000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 390000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 321500 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 321500 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 321500 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 336000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 336000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 390000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 390000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 321500 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 321500 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 321500 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 336000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 336000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 390000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 390000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 321500 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 321500 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 321500 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
