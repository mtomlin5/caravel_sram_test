magic
tech sky130A
magscale 1 2
timestamp 1636725598
<< locali >>
rect 257905 390303 257939 390609
rect 247417 390235 247451 390269
rect 247417 390201 248337 390235
rect 249107 388161 249625 388195
rect 236745 386427 236779 387821
rect 240885 386563 240919 387889
rect 235089 336515 235123 337977
rect 236653 336651 236687 337841
rect 237849 336991 237883 337841
rect 236595 336617 236687 336651
rect 235273 336515 235307 336617
rect 233801 336175 233835 336345
rect 235641 335563 235675 336073
rect 236653 336039 236687 336617
rect 238677 336039 238711 336073
rect 238527 336005 238711 336039
rect 238769 335971 238803 337909
rect 239079 336685 239321 336719
rect 235031 335529 235675 335563
rect 238677 335937 238803 335971
rect 235181 335359 235215 335461
rect 238677 333251 238711 335937
rect 239229 335767 239263 336617
rect 239321 335699 239355 336345
rect 239505 335495 239539 335733
rect 238769 334271 238803 335393
rect 238953 334475 238987 334645
rect 238861 334271 238895 334441
rect 240425 333523 240459 337909
rect 240701 337535 240735 337841
rect 240885 331959 240919 337705
rect 240977 333251 241011 337773
rect 241345 336447 241379 337025
rect 241195 336345 241437 336379
rect 241897 336277 241989 336311
rect 241897 336107 241931 336277
rect 241655 336073 241931 336107
rect 242357 336039 242391 337909
rect 242633 336243 242667 337773
rect 242817 337603 242851 337909
rect 242909 336447 242943 336753
rect 242449 335427 242483 336005
rect 242817 335563 242851 335937
rect 243277 335767 243311 337909
rect 243369 336515 243403 337773
rect 242081 335393 242483 335427
rect 243461 335427 243495 337909
rect 242081 335359 242115 335393
rect 243737 333319 243771 337909
rect 244013 335903 244047 336277
rect 244105 334475 244139 336277
rect 244933 333795 244967 337841
rect 245025 336175 245059 337909
rect 245209 337603 245243 337909
rect 245301 336379 245335 337909
rect 245485 336651 245519 337773
rect 245577 332231 245611 337773
rect 245853 333251 245887 337773
rect 245945 333931 245979 337909
rect 247233 334611 247267 337841
rect 247601 333047 247635 337773
rect 248061 333183 248095 337841
rect 248981 335495 249015 336821
rect 249165 335427 249199 336753
rect 249717 333999 249751 337909
rect 249901 332435 249935 337909
rect 250085 334815 250119 337705
rect 250361 334883 250395 337841
rect 250545 333183 250579 337977
rect 251281 335699 251315 337705
rect 251557 337535 251591 337909
rect 251741 333183 251775 337841
rect 252201 332843 252235 337909
rect 252753 336107 252787 337841
rect 253029 336447 253063 337841
rect 253489 332775 253523 337773
rect 254225 335767 254259 337909
rect 255513 337467 255547 337841
rect 255605 337535 255639 337841
rect 257169 337603 257203 337909
rect 257537 337671 257571 337909
rect 257629 335971 257663 337773
rect 257721 336175 257755 337909
rect 258089 333455 258123 337841
rect 259285 335291 259319 337909
rect 260481 336379 260515 337841
rect 260573 333999 260607 337909
rect 261861 332775 261895 337909
rect 262229 334475 262263 336073
rect 262873 335835 262907 335937
rect 262965 335903 262999 337773
rect 262781 335699 262815 335801
rect 263241 335767 263275 337841
rect 262873 332367 262907 335529
rect 263333 332435 263367 337909
rect 263425 336107 263459 337841
rect 263517 335359 263551 336413
rect 263885 333183 263919 337773
rect 266093 335699 266127 336821
rect 266645 336243 266679 337909
rect 267105 333047 267139 337841
rect 267381 336311 267415 337909
rect 267473 335631 267507 335733
rect 267657 333931 267691 337841
rect 267749 333319 267783 337705
rect 267933 333319 267967 337841
rect 268117 337399 268151 337909
rect 269163 336617 269347 336651
rect 269313 336175 269347 336617
rect 268945 335155 268979 335529
rect 269865 335291 269899 335733
rect 269957 335223 269991 335597
rect 270049 335155 270083 337909
rect 270267 336005 270359 336039
rect 270325 335359 270359 336005
rect 270417 333591 270451 337909
rect 270785 336515 270819 336685
rect 270785 336481 270969 336515
rect 270693 335563 270727 335801
rect 270877 332299 270911 336141
rect 271061 333523 271095 337909
rect 271429 333455 271463 337909
rect 272199 337841 272291 337875
rect 271705 333387 271739 335665
rect 271797 333319 271831 337773
rect 271981 335495 272015 337841
rect 272073 335563 272107 336753
rect 272165 336243 272199 336753
rect 271463 333149 272199 333183
rect 272165 332911 272199 333149
rect 272257 330259 272291 337841
rect 272625 330191 272659 337773
rect 272809 337535 272843 337909
rect 273361 337263 273395 337841
rect 272901 336651 272935 336957
rect 272993 336583 273027 337025
rect 273085 335971 273119 336549
rect 273361 336175 273395 337025
rect 273453 336243 273487 336957
rect 273027 335937 273119 335971
rect 273177 335767 273211 335937
rect 273119 335733 273211 335767
rect 273729 334543 273763 334645
rect 273821 334611 273855 334781
rect 273913 334645 274005 334679
rect 273913 334543 273947 334645
rect 274097 334611 274131 337909
rect 274373 337603 274407 337773
rect 274557 336719 274591 337977
rect 274741 335971 274775 336753
rect 275293 335291 275327 337841
rect 276397 337535 276431 337909
rect 275845 334815 275879 336073
rect 275937 335971 275971 336209
rect 276949 335359 276983 336073
rect 277225 335767 277259 337909
rect 277317 335223 277351 335869
rect 277409 335223 277443 337161
rect 277501 335903 277535 337841
rect 277593 336175 277627 336209
rect 277593 336141 278421 336175
rect 277777 336073 278605 336107
rect 277777 335971 277811 336073
rect 278697 335971 278731 336889
rect 278789 334951 278823 337909
rect 279433 335155 279467 337909
rect 279617 337671 279651 338045
rect 279893 337399 279927 337909
rect 279433 335121 279525 335155
rect 280445 334815 280479 335869
rect 280537 335699 280571 337841
rect 280445 334781 280537 334815
rect 280721 334747 280755 337909
rect 273729 334509 273947 334543
rect 280111 332265 280445 332299
rect 281181 330599 281215 337841
rect 281825 330531 281859 337773
rect 282009 334611 282043 337841
rect 282469 336107 282503 338113
rect 282561 336719 282595 336957
rect 282377 334339 282411 335257
rect 282469 334951 282503 335121
rect 282561 334475 282595 334917
rect 282653 334339 282687 338045
rect 282745 335427 282779 335597
rect 282837 335427 282871 337093
rect 282929 335937 283147 335971
rect 282929 335631 282963 335937
rect 283021 335359 283055 335869
rect 283113 335835 283147 335937
rect 284769 335563 284803 335665
rect 284343 335393 285413 335427
rect 282963 335325 283055 335359
rect 285597 335359 285631 336957
rect 286517 335631 286551 335801
rect 287345 335563 287379 335869
rect 284861 331279 284895 331653
rect 240701 321079 240735 326417
rect 441445 239853 441537 239887
rect 441445 239343 441479 239853
rect 441387 239309 441479 239343
rect 441537 239275 441571 239309
rect 441295 239241 441571 239275
rect 456717 236079 456751 239649
rect 298109 5457 298293 5491
rect 298109 5423 298143 5457
rect 281733 5049 282285 5083
rect 281733 4879 281767 5049
rect 282135 4981 282377 5015
rect 293083 4709 293785 4743
rect 128369 2907 128403 3009
rect 233893 2839 233927 4097
rect 239137 3383 239171 3689
rect 296085 3655 296119 3961
rect 296085 3621 296269 3655
<< viali >>
rect 257905 390609 257939 390643
rect 247417 390269 247451 390303
rect 257905 390269 257939 390303
rect 248337 390201 248371 390235
rect 249073 388161 249107 388195
rect 249625 388161 249659 388195
rect 240885 387889 240919 387923
rect 236745 387821 236779 387855
rect 240885 386529 240919 386563
rect 236745 386393 236779 386427
rect 282469 338113 282503 338147
rect 279617 338045 279651 338079
rect 235089 337977 235123 338011
rect 250545 337977 250579 338011
rect 238769 337909 238803 337943
rect 236653 337841 236687 337875
rect 237849 337841 237883 337875
rect 237849 336957 237883 336991
rect 235089 336481 235123 336515
rect 235273 336617 235307 336651
rect 236561 336617 236595 336651
rect 235273 336481 235307 336515
rect 233801 336345 233835 336379
rect 233801 336141 233835 336175
rect 235641 336073 235675 336107
rect 238677 336073 238711 336107
rect 236653 336005 236687 336039
rect 238493 336005 238527 336039
rect 240425 337909 240459 337943
rect 239045 336685 239079 336719
rect 239321 336685 239355 336719
rect 234997 335529 235031 335563
rect 239229 336617 239263 336651
rect 235181 335461 235215 335495
rect 235181 335325 235215 335359
rect 239229 335733 239263 335767
rect 239321 336345 239355 336379
rect 239321 335665 239355 335699
rect 239505 335733 239539 335767
rect 239505 335461 239539 335495
rect 238769 335393 238803 335427
rect 238953 334645 238987 334679
rect 238769 334237 238803 334271
rect 238861 334441 238895 334475
rect 238953 334441 238987 334475
rect 238861 334237 238895 334271
rect 242357 337909 242391 337943
rect 240701 337841 240735 337875
rect 240977 337773 241011 337807
rect 240701 337501 240735 337535
rect 240885 337705 240919 337739
rect 240425 333489 240459 333523
rect 238677 333217 238711 333251
rect 241345 337025 241379 337059
rect 241345 336413 241379 336447
rect 241161 336345 241195 336379
rect 241437 336345 241471 336379
rect 241989 336277 242023 336311
rect 241621 336073 241655 336107
rect 242817 337909 242851 337943
rect 242633 337773 242667 337807
rect 242817 337569 242851 337603
rect 243277 337909 243311 337943
rect 242909 336753 242943 336787
rect 242909 336413 242943 336447
rect 242633 336209 242667 336243
rect 242357 336005 242391 336039
rect 242449 336005 242483 336039
rect 242817 335937 242851 335971
rect 243461 337909 243495 337943
rect 243369 337773 243403 337807
rect 243369 336481 243403 336515
rect 243277 335733 243311 335767
rect 242817 335529 242851 335563
rect 243461 335393 243495 335427
rect 243737 337909 243771 337943
rect 242081 335325 242115 335359
rect 245025 337909 245059 337943
rect 244933 337841 244967 337875
rect 244013 336277 244047 336311
rect 244013 335869 244047 335903
rect 244105 336277 244139 336311
rect 244105 334441 244139 334475
rect 245209 337909 245243 337943
rect 245209 337569 245243 337603
rect 245301 337909 245335 337943
rect 245945 337909 245979 337943
rect 245485 337773 245519 337807
rect 245485 336617 245519 336651
rect 245577 337773 245611 337807
rect 245301 336345 245335 336379
rect 245025 336141 245059 336175
rect 244933 333761 244967 333795
rect 243737 333285 243771 333319
rect 240977 333217 241011 333251
rect 245853 337773 245887 337807
rect 249717 337909 249751 337943
rect 247233 337841 247267 337875
rect 248061 337841 248095 337875
rect 247233 334577 247267 334611
rect 247601 337773 247635 337807
rect 245945 333897 245979 333931
rect 245853 333217 245887 333251
rect 248981 336821 249015 336855
rect 248981 335461 249015 335495
rect 249165 336753 249199 336787
rect 249165 335393 249199 335427
rect 249717 333965 249751 333999
rect 249901 337909 249935 337943
rect 248061 333149 248095 333183
rect 247601 333013 247635 333047
rect 250361 337841 250395 337875
rect 250085 337705 250119 337739
rect 250361 334849 250395 334883
rect 250085 334781 250119 334815
rect 274557 337977 274591 338011
rect 251557 337909 251591 337943
rect 251281 337705 251315 337739
rect 252201 337909 252235 337943
rect 251557 337501 251591 337535
rect 251741 337841 251775 337875
rect 251281 335665 251315 335699
rect 250545 333149 250579 333183
rect 251741 333149 251775 333183
rect 254225 337909 254259 337943
rect 252753 337841 252787 337875
rect 253029 337841 253063 337875
rect 253029 336413 253063 336447
rect 253489 337773 253523 337807
rect 252753 336073 252787 336107
rect 252201 332809 252235 332843
rect 257169 337909 257203 337943
rect 255513 337841 255547 337875
rect 255605 337841 255639 337875
rect 257537 337909 257571 337943
rect 257721 337909 257755 337943
rect 257537 337637 257571 337671
rect 257629 337773 257663 337807
rect 257169 337569 257203 337603
rect 255605 337501 255639 337535
rect 255513 337433 255547 337467
rect 259285 337909 259319 337943
rect 257721 336141 257755 336175
rect 258089 337841 258123 337875
rect 257629 335937 257663 335971
rect 254225 335733 254259 335767
rect 260573 337909 260607 337943
rect 260481 337841 260515 337875
rect 260481 336345 260515 336379
rect 259285 335257 259319 335291
rect 260573 333965 260607 333999
rect 261861 337909 261895 337943
rect 258089 333421 258123 333455
rect 253489 332741 253523 332775
rect 263333 337909 263367 337943
rect 263241 337841 263275 337875
rect 262965 337773 262999 337807
rect 262229 336073 262263 336107
rect 262873 335937 262907 335971
rect 262965 335869 262999 335903
rect 262781 335801 262815 335835
rect 262873 335801 262907 335835
rect 263241 335733 263275 335767
rect 262781 335665 262815 335699
rect 262229 334441 262263 334475
rect 262873 335529 262907 335563
rect 261861 332741 261895 332775
rect 249901 332401 249935 332435
rect 266645 337909 266679 337943
rect 263425 337841 263459 337875
rect 263885 337773 263919 337807
rect 263425 336073 263459 336107
rect 263517 336413 263551 336447
rect 263517 335325 263551 335359
rect 266093 336821 266127 336855
rect 267381 337909 267415 337943
rect 266645 336209 266679 336243
rect 267105 337841 267139 337875
rect 266093 335665 266127 335699
rect 263885 333149 263919 333183
rect 268117 337909 268151 337943
rect 267381 336277 267415 336311
rect 267657 337841 267691 337875
rect 267473 335733 267507 335767
rect 267473 335597 267507 335631
rect 267933 337841 267967 337875
rect 267657 333897 267691 333931
rect 267749 337705 267783 337739
rect 267749 333285 267783 333319
rect 268117 337365 268151 337399
rect 270049 337909 270083 337943
rect 269129 336617 269163 336651
rect 269313 336141 269347 336175
rect 269865 335733 269899 335767
rect 268945 335529 268979 335563
rect 269865 335257 269899 335291
rect 269957 335597 269991 335631
rect 269957 335189 269991 335223
rect 268945 335121 268979 335155
rect 270417 337909 270451 337943
rect 270233 336005 270267 336039
rect 270325 335325 270359 335359
rect 270049 335121 270083 335155
rect 271061 337909 271095 337943
rect 270785 336685 270819 336719
rect 270969 336481 271003 336515
rect 270877 336141 270911 336175
rect 270693 335801 270727 335835
rect 270693 335529 270727 335563
rect 270417 333557 270451 333591
rect 267933 333285 267967 333319
rect 267105 333013 267139 333047
rect 263333 332401 263367 332435
rect 262873 332333 262907 332367
rect 271061 333489 271095 333523
rect 271429 337909 271463 337943
rect 272809 337909 272843 337943
rect 271981 337841 272015 337875
rect 272165 337841 272199 337875
rect 271797 337773 271831 337807
rect 271429 333421 271463 333455
rect 271705 335665 271739 335699
rect 271705 333353 271739 333387
rect 272073 336753 272107 336787
rect 272165 336753 272199 336787
rect 272165 336209 272199 336243
rect 272073 335529 272107 335563
rect 271981 335461 272015 335495
rect 271797 333285 271831 333319
rect 271429 333149 271463 333183
rect 272165 332877 272199 332911
rect 270877 332265 270911 332299
rect 245577 332197 245611 332231
rect 240885 331925 240919 331959
rect 272257 330225 272291 330259
rect 272625 337773 272659 337807
rect 274097 337909 274131 337943
rect 272809 337501 272843 337535
rect 273361 337841 273395 337875
rect 273361 337229 273395 337263
rect 272993 337025 273027 337059
rect 272901 336957 272935 336991
rect 272901 336617 272935 336651
rect 273361 337025 273395 337059
rect 272993 336549 273027 336583
rect 273085 336549 273119 336583
rect 273453 336957 273487 336991
rect 273453 336209 273487 336243
rect 273361 336141 273395 336175
rect 272993 335937 273027 335971
rect 273177 335937 273211 335971
rect 273085 335733 273119 335767
rect 273821 334781 273855 334815
rect 273729 334645 273763 334679
rect 273821 334577 273855 334611
rect 274005 334645 274039 334679
rect 274373 337773 274407 337807
rect 274373 337569 274407 337603
rect 276397 337909 276431 337943
rect 275293 337841 275327 337875
rect 274557 336685 274591 336719
rect 274741 336753 274775 336787
rect 274741 335937 274775 335971
rect 276397 337501 276431 337535
rect 277225 337909 277259 337943
rect 275937 336209 275971 336243
rect 275293 335257 275327 335291
rect 275845 336073 275879 336107
rect 275937 335937 275971 335971
rect 276949 336073 276983 336107
rect 278789 337909 278823 337943
rect 277501 337841 277535 337875
rect 277409 337161 277443 337195
rect 277225 335733 277259 335767
rect 277317 335869 277351 335903
rect 276949 335325 276983 335359
rect 277317 335189 277351 335223
rect 278697 336889 278731 336923
rect 277593 336209 277627 336243
rect 278421 336141 278455 336175
rect 278605 336073 278639 336107
rect 277777 335937 277811 335971
rect 278697 335937 278731 335971
rect 277501 335869 277535 335903
rect 277409 335189 277443 335223
rect 279433 337909 279467 337943
rect 279617 337637 279651 337671
rect 279893 337909 279927 337943
rect 280721 337909 280755 337943
rect 279893 337365 279927 337399
rect 280537 337841 280571 337875
rect 280445 335869 280479 335903
rect 279525 335121 279559 335155
rect 278789 334917 278823 334951
rect 275845 334781 275879 334815
rect 280537 335665 280571 335699
rect 280537 334781 280571 334815
rect 280721 334713 280755 334747
rect 281181 337841 281215 337875
rect 274097 334577 274131 334611
rect 280077 332265 280111 332299
rect 280445 332265 280479 332299
rect 282009 337841 282043 337875
rect 281181 330565 281215 330599
rect 281825 337773 281859 337807
rect 282653 338045 282687 338079
rect 282561 336957 282595 336991
rect 282561 336685 282595 336719
rect 282469 336073 282503 336107
rect 282009 334577 282043 334611
rect 282377 335257 282411 335291
rect 282469 335121 282503 335155
rect 282469 334917 282503 334951
rect 282561 334917 282595 334951
rect 282561 334441 282595 334475
rect 282377 334305 282411 334339
rect 282837 337093 282871 337127
rect 282745 335597 282779 335631
rect 282745 335393 282779 335427
rect 285597 336957 285631 336991
rect 282929 335597 282963 335631
rect 283021 335869 283055 335903
rect 282837 335393 282871 335427
rect 283113 335801 283147 335835
rect 284769 335665 284803 335699
rect 284769 335529 284803 335563
rect 284309 335393 284343 335427
rect 285413 335393 285447 335427
rect 282929 335325 282963 335359
rect 287345 335869 287379 335903
rect 286517 335801 286551 335835
rect 286517 335597 286551 335631
rect 287345 335529 287379 335563
rect 285597 335325 285631 335359
rect 282653 334305 282687 334339
rect 284861 331653 284895 331687
rect 284861 331245 284895 331279
rect 281825 330497 281859 330531
rect 272625 330157 272659 330191
rect 240701 326417 240735 326451
rect 240701 321045 240735 321079
rect 441537 239853 441571 239887
rect 456717 239649 456751 239683
rect 441353 239309 441387 239343
rect 441537 239309 441571 239343
rect 441261 239241 441295 239275
rect 456717 236045 456751 236079
rect 298293 5457 298327 5491
rect 298109 5389 298143 5423
rect 282285 5049 282319 5083
rect 282101 4981 282135 5015
rect 282377 4981 282411 5015
rect 281733 4845 281767 4879
rect 293049 4709 293083 4743
rect 293785 4709 293819 4743
rect 233893 4097 233927 4131
rect 128369 3009 128403 3043
rect 128369 2873 128403 2907
rect 296085 3961 296119 3995
rect 239137 3689 239171 3723
rect 296269 3621 296303 3655
rect 239137 3349 239171 3383
rect 233893 2805 233927 2839
<< metal1 >>
rect 105446 700952 105452 701004
rect 105504 700992 105510 701004
rect 262214 700992 262220 701004
rect 105504 700964 262220 700992
rect 105504 700952 105510 700964
rect 262214 700952 262220 700964
rect 262272 700952 262278 701004
rect 256510 700884 256516 700936
rect 256568 700924 256574 700936
rect 429838 700924 429844 700936
rect 256568 700896 429844 700924
rect 256568 700884 256574 700896
rect 429838 700884 429844 700896
rect 429896 700884 429902 700936
rect 89162 700816 89168 700868
rect 89220 700856 89226 700868
rect 262306 700856 262312 700868
rect 89220 700828 262312 700856
rect 89220 700816 89226 700828
rect 262306 700816 262312 700828
rect 262364 700816 262370 700868
rect 72970 700748 72976 700800
rect 73028 700788 73034 700800
rect 262490 700788 262496 700800
rect 73028 700760 262496 700788
rect 73028 700748 73034 700760
rect 262490 700748 262496 700760
rect 262548 700748 262554 700800
rect 256418 700680 256424 700732
rect 256476 700720 256482 700732
rect 462314 700720 462320 700732
rect 256476 700692 462320 700720
rect 256476 700680 256482 700692
rect 462314 700680 462320 700692
rect 462372 700680 462378 700732
rect 256602 700612 256608 700664
rect 256660 700652 256666 700664
rect 478506 700652 478512 700664
rect 256660 700624 478512 700652
rect 256660 700612 256666 700624
rect 478506 700612 478512 700624
rect 478564 700612 478570 700664
rect 40494 700544 40500 700596
rect 40552 700584 40558 700596
rect 263686 700584 263692 700596
rect 40552 700556 263692 700584
rect 40552 700544 40558 700556
rect 263686 700544 263692 700556
rect 263744 700544 263750 700596
rect 24302 700476 24308 700528
rect 24360 700516 24366 700528
rect 263594 700516 263600 700528
rect 24360 700488 263600 700516
rect 24360 700476 24366 700488
rect 263594 700476 263600 700488
rect 263652 700476 263658 700528
rect 283650 700476 283656 700528
rect 283708 700516 283714 700528
rect 300118 700516 300124 700528
rect 283708 700488 300124 700516
rect 283708 700476 283714 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 8110 700408 8116 700460
rect 8168 700448 8174 700460
rect 263778 700448 263784 700460
rect 8168 700420 263784 700448
rect 8168 700408 8174 700420
rect 263778 700408 263784 700420
rect 263836 700408 263842 700460
rect 269758 700408 269764 700460
rect 269816 700448 269822 700460
rect 283834 700448 283840 700460
rect 269816 700420 283840 700448
rect 269816 700408 269822 700420
rect 283834 700408 283840 700420
rect 283892 700408 283898 700460
rect 283926 700408 283932 700460
rect 283984 700448 283990 700460
rect 364978 700448 364984 700460
rect 283984 700420 364984 700448
rect 283984 700408 283990 700420
rect 364978 700408 364984 700420
rect 365036 700408 365042 700460
rect 255130 700340 255136 700392
rect 255188 700380 255194 700392
rect 527174 700380 527180 700392
rect 255188 700352 527180 700380
rect 255188 700340 255194 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 255038 700272 255044 700324
rect 255096 700312 255102 700324
rect 543458 700312 543464 700324
rect 255096 700284 543464 700312
rect 255096 700272 255102 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 257706 700204 257712 700256
rect 257764 700244 257770 700256
rect 413646 700244 413652 700256
rect 257764 700216 413652 700244
rect 257764 700204 257770 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 257798 700136 257804 700188
rect 257856 700176 257862 700188
rect 397454 700176 397460 700188
rect 257856 700148 397460 700176
rect 257856 700136 257862 700148
rect 397454 700136 397460 700148
rect 397512 700136 397518 700188
rect 137830 700068 137836 700120
rect 137888 700108 137894 700120
rect 260926 700108 260932 700120
rect 137888 700080 260932 700108
rect 137888 700068 137894 700080
rect 260926 700068 260932 700080
rect 260984 700068 260990 700120
rect 154114 700000 154120 700052
rect 154172 700040 154178 700052
rect 262398 700040 262404 700052
rect 154172 700012 262404 700040
rect 154172 700000 154178 700012
rect 262398 700000 262404 700012
rect 262456 700000 262462 700052
rect 170306 699932 170312 699984
rect 170364 699972 170370 699984
rect 260834 699972 260840 699984
rect 170364 699944 260840 699972
rect 170364 699932 170370 699944
rect 260834 699932 260840 699944
rect 260892 699932 260898 699984
rect 259178 699864 259184 699916
rect 259236 699904 259242 699916
rect 348786 699904 348792 699916
rect 259236 699876 348792 699904
rect 259236 699864 259242 699876
rect 348786 699864 348792 699876
rect 348844 699864 348850 699916
rect 235166 699796 235172 699848
rect 235224 699836 235230 699848
rect 235902 699836 235908 699848
rect 235224 699808 235908 699836
rect 235224 699796 235230 699808
rect 235902 699796 235908 699808
rect 235960 699796 235966 699848
rect 257890 699796 257896 699848
rect 257948 699836 257954 699848
rect 332502 699836 332508 699848
rect 257948 699808 332508 699836
rect 257948 699796 257954 699808
rect 332502 699796 332508 699808
rect 332560 699796 332566 699848
rect 202782 699728 202788 699780
rect 202840 699768 202846 699780
rect 259638 699768 259644 699780
rect 202840 699740 259644 699768
rect 202840 699728 202846 699740
rect 259638 699728 259644 699740
rect 259696 699728 259702 699780
rect 218974 699660 218980 699712
rect 219032 699700 219038 699712
rect 261018 699700 261024 699712
rect 219032 699672 261024 699700
rect 219032 699660 219038 699672
rect 261018 699660 261024 699672
rect 261076 699660 261082 699712
rect 261478 699660 261484 699712
rect 261536 699700 261542 699712
rect 267642 699700 267648 699712
rect 261536 699672 267648 699700
rect 261536 699660 261542 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 283558 699660 283564 699712
rect 283616 699700 283622 699712
rect 283926 699700 283932 699712
rect 283616 699672 283932 699700
rect 283616 699660 283622 699672
rect 283926 699660 283932 699672
rect 283984 699660 283990 699712
rect 253566 696940 253572 696992
rect 253624 696980 253630 696992
rect 580166 696980 580172 696992
rect 253624 696952 580172 696980
rect 253624 696940 253630 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 264974 683244 264980 683256
rect 3476 683216 264980 683244
rect 3476 683204 3482 683216
rect 264974 683204 264980 683216
rect 265032 683204 265038 683256
rect 253750 683136 253756 683188
rect 253808 683176 253814 683188
rect 580166 683176 580172 683188
rect 253808 683148 580172 683176
rect 253808 683136 253814 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3418 670760 3424 670812
rect 3476 670800 3482 670812
rect 265066 670800 265072 670812
rect 3476 670772 265072 670800
rect 3476 670760 3482 670772
rect 265066 670760 265072 670772
rect 265124 670760 265130 670812
rect 253658 670692 253664 670744
rect 253716 670732 253722 670744
rect 580166 670732 580172 670744
rect 253716 670704 580172 670732
rect 253716 670692 253722 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 265158 656928 265164 656940
rect 3476 656900 265164 656928
rect 3476 656888 3482 656900
rect 265158 656888 265164 656900
rect 265216 656888 265222 656940
rect 252462 643084 252468 643136
rect 252520 643124 252526 643136
rect 580166 643124 580172 643136
rect 252520 643096 580172 643124
rect 252520 643084 252526 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 266354 632108 266360 632120
rect 3476 632080 266360 632108
rect 3476 632068 3482 632080
rect 266354 632068 266360 632080
rect 266412 632068 266418 632120
rect 252370 630640 252376 630692
rect 252428 630680 252434 630692
rect 580166 630680 580172 630692
rect 252428 630652 580172 630680
rect 252428 630640 252434 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 266446 618304 266452 618316
rect 3200 618276 266452 618304
rect 3200 618264 3206 618276
rect 266446 618264 266452 618276
rect 266504 618264 266510 618316
rect 252278 616836 252284 616888
rect 252336 616876 252342 616888
rect 580166 616876 580172 616888
rect 252336 616848 580172 616876
rect 252336 616836 252342 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 266538 605860 266544 605872
rect 3292 605832 266544 605860
rect 3292 605820 3298 605832
rect 266538 605820 266544 605832
rect 266596 605820 266602 605872
rect 251082 590656 251088 590708
rect 251140 590696 251146 590708
rect 579798 590696 579804 590708
rect 251140 590668 579804 590696
rect 251140 590656 251146 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 266630 579680 266636 579692
rect 3384 579652 266636 579680
rect 3384 579640 3390 579652
rect 266630 579640 266636 579652
rect 266688 579640 266694 579692
rect 250990 576852 250996 576904
rect 251048 576892 251054 576904
rect 580166 576892 580172 576904
rect 251048 576864 580172 576892
rect 251048 576852 251054 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 267734 565876 267740 565888
rect 3476 565848 267740 565876
rect 3476 565836 3482 565848
rect 267734 565836 267740 565848
rect 267792 565836 267798 565888
rect 250898 563048 250904 563100
rect 250956 563088 250962 563100
rect 579798 563088 579804 563100
rect 250956 563060 579804 563088
rect 250956 563048 250962 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 267826 553432 267832 553444
rect 3476 553404 267832 553432
rect 3476 553392 3482 553404
rect 267826 553392 267832 553404
rect 267884 553392 267890 553444
rect 249702 536800 249708 536852
rect 249760 536840 249766 536852
rect 580166 536840 580172 536852
rect 249760 536812 580172 536840
rect 249760 536800 249766 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 267918 527184 267924 527196
rect 3476 527156 267924 527184
rect 3476 527144 3482 527156
rect 267918 527144 267924 527156
rect 267976 527144 267982 527196
rect 249610 524424 249616 524476
rect 249668 524464 249674 524476
rect 580166 524464 580172 524476
rect 249668 524436 580172 524464
rect 249668 524424 249674 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 269114 514808 269120 514820
rect 3476 514780 269120 514808
rect 3476 514768 3482 514780
rect 269114 514768 269120 514780
rect 269172 514768 269178 514820
rect 249518 510620 249524 510672
rect 249576 510660 249582 510672
rect 580166 510660 580172 510672
rect 249576 510632 580172 510660
rect 249576 510620 249582 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 269206 501004 269212 501016
rect 3108 500976 269212 501004
rect 3108 500964 3114 500976
rect 269206 500964 269212 500976
rect 269264 500964 269270 501016
rect 248322 484372 248328 484424
rect 248380 484412 248386 484424
rect 580166 484412 580172 484424
rect 248380 484384 580172 484412
rect 248380 484372 248386 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 269298 474756 269304 474768
rect 3476 474728 269304 474756
rect 3476 474716 3482 474728
rect 269298 474716 269304 474728
rect 269356 474716 269362 474768
rect 249426 470568 249432 470620
rect 249484 470608 249490 470620
rect 579982 470608 579988 470620
rect 249484 470580 579988 470608
rect 249484 470568 249490 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 270770 462380 270776 462392
rect 3292 462352 270776 462380
rect 3292 462340 3298 462352
rect 270770 462340 270776 462352
rect 270828 462340 270834 462392
rect 248230 456764 248236 456816
rect 248288 456804 248294 456816
rect 580166 456804 580172 456816
rect 248288 456776 580172 456804
rect 248288 456764 248294 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 270586 448576 270592 448588
rect 3200 448548 270592 448576
rect 3200 448536 3206 448548
rect 270586 448536 270592 448548
rect 270644 448536 270650 448588
rect 259270 434664 259276 434716
rect 259328 434704 259334 434716
rect 261478 434704 261484 434716
rect 259328 434676 261484 434704
rect 259328 434664 259334 434676
rect 261478 434664 261484 434676
rect 261536 434664 261542 434716
rect 246942 430584 246948 430636
rect 247000 430624 247006 430636
rect 580166 430624 580172 430636
rect 247000 430596 580172 430624
rect 247000 430584 247006 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 270678 422328 270684 422340
rect 3476 422300 270684 422328
rect 3476 422288 3482 422300
rect 270678 422288 270684 422300
rect 270736 422288 270742 422340
rect 248138 418140 248144 418192
rect 248196 418180 248202 418192
rect 580166 418180 580172 418192
rect 248196 418152 580172 418180
rect 248196 418140 248202 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 271874 409884 271880 409896
rect 3200 409856 271880 409884
rect 3200 409844 3206 409856
rect 271874 409844 271880 409856
rect 271932 409844 271938 409896
rect 246850 404336 246856 404388
rect 246908 404376 246914 404388
rect 580166 404376 580172 404388
rect 246908 404348 580172 404376
rect 246908 404336 246914 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 270494 397508 270500 397520
rect 3476 397480 270500 397508
rect 3476 397468 3482 397480
rect 270494 397468 270500 397480
rect 270552 397468 270558 397520
rect 260834 391620 260840 391672
rect 260892 391660 260898 391672
rect 261110 391660 261116 391672
rect 260892 391632 261116 391660
rect 260892 391620 260898 391632
rect 261110 391620 261116 391632
rect 261168 391620 261174 391672
rect 259822 391592 259828 391604
rect 238726 391564 259828 391592
rect 235902 391484 235908 391536
rect 235960 391524 235966 391536
rect 238726 391524 238754 391564
rect 259822 391552 259828 391564
rect 259880 391552 259886 391604
rect 235960 391496 238754 391524
rect 235960 391484 235966 391496
rect 259638 391484 259644 391536
rect 259696 391524 259702 391536
rect 269758 391524 269764 391536
rect 259696 391496 269764 391524
rect 259696 391484 259702 391496
rect 269758 391484 269764 391496
rect 269816 391484 269822 391536
rect 259178 391416 259184 391468
rect 259236 391456 259242 391468
rect 283650 391456 283656 391468
rect 259236 391428 283656 391456
rect 259236 391416 259242 391428
rect 283650 391416 283656 391428
rect 283708 391416 283714 391468
rect 257890 391348 257896 391400
rect 257948 391388 257954 391400
rect 283558 391388 283564 391400
rect 257948 391360 283564 391388
rect 257948 391348 257954 391360
rect 283558 391348 283564 391360
rect 283616 391348 283622 391400
rect 255222 391280 255228 391332
rect 255280 391320 255286 391332
rect 494054 391320 494060 391332
rect 255280 391292 494060 391320
rect 255280 391280 255286 391292
rect 494054 391280 494060 391292
rect 494112 391280 494118 391332
rect 253842 391212 253848 391264
rect 253900 391252 253906 391264
rect 558914 391252 558920 391264
rect 253900 391224 558920 391252
rect 253900 391212 253906 391224
rect 558914 391212 558920 391224
rect 558972 391212 558978 391264
rect 257893 390643 257951 390649
rect 257893 390640 257905 390643
rect 248616 390612 257905 390640
rect 242066 390464 242072 390516
rect 242124 390504 242130 390516
rect 248616 390504 248644 390612
rect 257893 390609 257905 390612
rect 257939 390609 257951 390643
rect 257893 390603 257951 390609
rect 262306 390600 262312 390652
rect 262364 390640 262370 390652
rect 263226 390640 263232 390652
rect 262364 390612 263232 390640
rect 262364 390600 262370 390612
rect 263226 390600 263232 390612
rect 263284 390600 263290 390652
rect 249334 390532 249340 390584
rect 249392 390572 249398 390584
rect 249702 390572 249708 390584
rect 249392 390544 249708 390572
rect 249392 390532 249398 390544
rect 249702 390532 249708 390544
rect 249760 390532 249766 390584
rect 250806 390532 250812 390584
rect 250864 390572 250870 390584
rect 251082 390572 251088 390584
rect 250864 390544 251088 390572
rect 250864 390532 250870 390544
rect 251082 390532 251088 390544
rect 251140 390532 251146 390584
rect 260926 390532 260932 390584
rect 260984 390572 260990 390584
rect 261570 390572 261576 390584
rect 260984 390544 261576 390572
rect 260984 390532 260990 390544
rect 261570 390532 261576 390544
rect 261628 390532 261634 390584
rect 262214 390532 262220 390584
rect 262272 390572 262278 390584
rect 262490 390572 262496 390584
rect 262272 390544 262496 390572
rect 262272 390532 262278 390544
rect 262490 390532 262496 390544
rect 262548 390532 262554 390584
rect 263594 390532 263600 390584
rect 263652 390572 263658 390584
rect 264422 390572 264428 390584
rect 263652 390544 264428 390572
rect 263652 390532 263658 390544
rect 264422 390532 264428 390544
rect 264480 390532 264486 390584
rect 265066 390532 265072 390584
rect 265124 390572 265130 390584
rect 265710 390572 265716 390584
rect 265124 390544 265716 390572
rect 265124 390532 265130 390544
rect 265710 390532 265716 390544
rect 265768 390532 265774 390584
rect 266446 390532 266452 390584
rect 266504 390572 266510 390584
rect 266906 390572 266912 390584
rect 266504 390544 266912 390572
rect 266504 390532 266510 390544
rect 266906 390532 266912 390544
rect 266964 390532 266970 390584
rect 267734 390532 267740 390584
rect 267792 390572 267798 390584
rect 268194 390572 268200 390584
rect 267792 390544 268200 390572
rect 267792 390532 267798 390544
rect 268194 390532 268200 390544
rect 268252 390532 268258 390584
rect 269114 390532 269120 390584
rect 269172 390572 269178 390584
rect 269482 390572 269488 390584
rect 269172 390544 269488 390572
rect 269172 390532 269178 390544
rect 269482 390532 269488 390544
rect 269540 390532 269546 390584
rect 270678 390532 270684 390584
rect 270736 390572 270742 390584
rect 271138 390572 271144 390584
rect 270736 390544 271144 390572
rect 270736 390532 270742 390544
rect 271138 390532 271144 390544
rect 271196 390532 271202 390584
rect 289078 390504 289084 390516
rect 242124 390476 248644 390504
rect 248708 390476 289084 390504
rect 242124 390464 242130 390476
rect 246298 390396 246304 390448
rect 246356 390436 246362 390448
rect 248708 390436 248736 390476
rect 289078 390464 289084 390476
rect 289136 390464 289142 390516
rect 288986 390436 288992 390448
rect 246356 390408 248736 390436
rect 248800 390408 288992 390436
rect 246356 390396 246362 390408
rect 245010 390328 245016 390380
rect 245068 390368 245074 390380
rect 248800 390368 248828 390408
rect 288986 390396 288992 390408
rect 289044 390396 289050 390448
rect 537478 390368 537484 390380
rect 245068 390340 248828 390368
rect 248892 390340 537484 390368
rect 245068 390328 245074 390340
rect 240042 390260 240048 390312
rect 240100 390300 240106 390312
rect 247405 390303 247463 390309
rect 247405 390300 247417 390303
rect 240100 390272 247417 390300
rect 240100 390260 240106 390272
rect 247405 390269 247417 390272
rect 247451 390269 247463 390303
rect 247405 390263 247463 390269
rect 247494 390260 247500 390312
rect 247552 390300 247558 390312
rect 248138 390300 248144 390312
rect 247552 390272 248144 390300
rect 247552 390260 247558 390272
rect 248138 390260 248144 390272
rect 248196 390260 248202 390312
rect 248892 390300 248920 390340
rect 537478 390328 537484 390340
rect 537536 390328 537542 390380
rect 248248 390272 248920 390300
rect 243814 390192 243820 390244
rect 243872 390232 243878 390244
rect 248248 390232 248276 390272
rect 248966 390260 248972 390312
rect 249024 390300 249030 390312
rect 249426 390300 249432 390312
rect 249024 390272 249432 390300
rect 249024 390260 249030 390272
rect 249426 390260 249432 390272
rect 249484 390260 249490 390312
rect 250438 390260 250444 390312
rect 250496 390300 250502 390312
rect 250898 390300 250904 390312
rect 250496 390272 250904 390300
rect 250496 390260 250502 390272
rect 250898 390260 250904 390272
rect 250956 390260 250962 390312
rect 252094 390260 252100 390312
rect 252152 390300 252158 390312
rect 252462 390300 252468 390312
rect 252152 390272 252468 390300
rect 252152 390260 252158 390272
rect 252462 390260 252468 390272
rect 252520 390260 252526 390312
rect 252922 390260 252928 390312
rect 252980 390300 252986 390312
rect 253658 390300 253664 390312
rect 252980 390272 253664 390300
rect 252980 390260 252986 390272
rect 253658 390260 253664 390272
rect 253716 390260 253722 390312
rect 254578 390260 254584 390312
rect 254636 390300 254642 390312
rect 255130 390300 255136 390312
rect 254636 390272 255136 390300
rect 254636 390260 254642 390272
rect 255130 390260 255136 390272
rect 255188 390260 255194 390312
rect 256234 390260 256240 390312
rect 256292 390300 256298 390312
rect 256602 390300 256608 390312
rect 256292 390272 256608 390300
rect 256292 390260 256298 390272
rect 256602 390260 256608 390272
rect 256660 390260 256666 390312
rect 257062 390260 257068 390312
rect 257120 390300 257126 390312
rect 257798 390300 257804 390312
rect 257120 390272 257804 390300
rect 257120 390260 257126 390272
rect 257798 390260 257804 390272
rect 257856 390260 257862 390312
rect 257893 390303 257951 390309
rect 257893 390269 257905 390303
rect 257939 390300 257951 390303
rect 286962 390300 286968 390312
rect 257939 390272 286968 390300
rect 257939 390269 257951 390272
rect 257893 390263 257951 390269
rect 286962 390260 286968 390272
rect 287020 390260 287026 390312
rect 243872 390204 248276 390232
rect 248325 390235 248383 390241
rect 243872 390192 243878 390204
rect 248325 390201 248337 390235
rect 248371 390232 248383 390235
rect 286778 390232 286784 390244
rect 248371 390204 286784 390232
rect 248371 390201 248383 390204
rect 248325 390195 248383 390201
rect 286778 390192 286784 390204
rect 286836 390192 286842 390244
rect 242526 390124 242532 390176
rect 242584 390164 242590 390176
rect 289722 390164 289728 390176
rect 242584 390136 289728 390164
rect 242584 390124 242590 390136
rect 289722 390124 289728 390136
rect 289780 390124 289786 390176
rect 238662 390056 238668 390108
rect 238720 390096 238726 390108
rect 286594 390096 286600 390108
rect 238720 390068 286600 390096
rect 238720 390056 238726 390068
rect 286594 390056 286600 390068
rect 286652 390056 286658 390108
rect 241146 389988 241152 390040
rect 241204 390028 241210 390040
rect 289630 390028 289636 390040
rect 241204 390000 289636 390028
rect 241204 389988 241210 390000
rect 289630 389988 289636 390000
rect 289688 389988 289694 390040
rect 4706 389920 4712 389972
rect 4764 389960 4770 389972
rect 4764 389932 270448 389960
rect 4764 389920 4770 389932
rect 5350 389852 5356 389904
rect 5408 389892 5414 389904
rect 270420 389892 270448 389932
rect 270494 389920 270500 389972
rect 270552 389960 270558 389972
rect 271506 389960 271512 389972
rect 270552 389932 271512 389960
rect 270552 389920 270558 389932
rect 271506 389920 271512 389932
rect 271564 389920 271570 389972
rect 271598 389920 271604 389972
rect 271656 389960 271662 389972
rect 276934 389960 276940 389972
rect 271656 389932 276940 389960
rect 271656 389920 271662 389932
rect 276934 389920 276940 389932
rect 276992 389920 276998 389972
rect 273254 389892 273260 389904
rect 5408 389864 270356 389892
rect 270420 389864 273260 389892
rect 5408 389852 5414 389864
rect 6546 389784 6552 389836
rect 6604 389824 6610 389836
rect 270218 389824 270224 389836
rect 6604 389796 270224 389824
rect 6604 389784 6610 389796
rect 270218 389784 270224 389796
rect 270276 389784 270282 389836
rect 270328 389824 270356 389864
rect 273254 389852 273260 389864
rect 273312 389852 273318 389904
rect 275646 389824 275652 389836
rect 270328 389796 275652 389824
rect 275646 389784 275652 389796
rect 275704 389784 275710 389836
rect 5166 389716 5172 389768
rect 5224 389756 5230 389768
rect 276474 389756 276480 389768
rect 5224 389728 276480 389756
rect 5224 389716 5230 389728
rect 276474 389716 276480 389728
rect 276532 389716 276538 389768
rect 6454 389648 6460 389700
rect 6512 389688 6518 389700
rect 278222 389688 278228 389700
rect 6512 389660 278228 389688
rect 6512 389648 6518 389660
rect 278222 389648 278228 389660
rect 278280 389648 278286 389700
rect 5074 389580 5080 389632
rect 5132 389620 5138 389632
rect 277762 389620 277768 389632
rect 5132 389592 277768 389620
rect 5132 389580 5138 389592
rect 277762 389580 277768 389592
rect 277820 389580 277826 389632
rect 284202 389580 284208 389632
rect 284260 389620 284266 389632
rect 292206 389620 292212 389632
rect 284260 389592 292212 389620
rect 284260 389580 284266 389592
rect 292206 389580 292212 389592
rect 292264 389580 292270 389632
rect 6362 389512 6368 389564
rect 6420 389552 6426 389564
rect 279418 389552 279424 389564
rect 6420 389524 279424 389552
rect 6420 389512 6426 389524
rect 279418 389512 279424 389524
rect 279476 389512 279482 389564
rect 284110 389512 284116 389564
rect 284168 389552 284174 389564
rect 292114 389552 292120 389564
rect 284168 389524 292120 389552
rect 284168 389512 284174 389524
rect 292114 389512 292120 389524
rect 292172 389512 292178 389564
rect 4982 389444 4988 389496
rect 5040 389484 5046 389496
rect 279050 389484 279056 389496
rect 5040 389456 279056 389484
rect 5040 389444 5046 389456
rect 279050 389444 279056 389456
rect 279108 389444 279114 389496
rect 283742 389444 283748 389496
rect 283800 389484 283806 389496
rect 298830 389484 298836 389496
rect 283800 389456 298836 389484
rect 283800 389444 283806 389456
rect 298830 389444 298836 389456
rect 298888 389444 298894 389496
rect 6270 389376 6276 389428
rect 6328 389416 6334 389428
rect 280706 389416 280712 389428
rect 6328 389388 280712 389416
rect 6328 389376 6334 389388
rect 280706 389376 280712 389388
rect 280764 389376 280770 389428
rect 285030 389376 285036 389428
rect 285088 389416 285094 389428
rect 292022 389416 292028 389428
rect 285088 389388 292028 389416
rect 285088 389376 285094 389388
rect 292022 389376 292028 389388
rect 292080 389376 292086 389428
rect 4890 389308 4896 389360
rect 4948 389348 4954 389360
rect 280246 389348 280252 389360
rect 4948 389320 280252 389348
rect 4948 389308 4954 389320
rect 280246 389308 280252 389320
rect 280304 389308 280310 389360
rect 283282 389308 283288 389360
rect 283340 389348 283346 389360
rect 294598 389348 294604 389360
rect 283340 389320 294604 389348
rect 283340 389308 283346 389320
rect 294598 389308 294604 389320
rect 294656 389308 294662 389360
rect 243354 389240 243360 389292
rect 243412 389280 243418 389292
rect 537570 389280 537576 389292
rect 243412 389252 537576 389280
rect 243412 389240 243418 389252
rect 537570 389240 537576 389252
rect 537628 389240 537634 389292
rect 6638 389172 6644 389224
rect 6696 389212 6702 389224
rect 274634 389212 274640 389224
rect 6696 389184 274640 389212
rect 6696 389172 6702 389184
rect 274634 389172 274640 389184
rect 274692 389172 274698 389224
rect 282822 389172 282828 389224
rect 282880 389212 282886 389224
rect 293310 389212 293316 389224
rect 282880 389184 293316 389212
rect 282880 389172 282886 389184
rect 293310 389172 293316 389184
rect 293368 389172 293374 389224
rect 5442 389104 5448 389156
rect 5500 389144 5506 389156
rect 272794 389144 272800 389156
rect 5500 389116 272800 389144
rect 5500 389104 5506 389116
rect 272794 389104 272800 389116
rect 272852 389104 272858 389156
rect 3326 389036 3332 389088
rect 3384 389076 3390 389088
rect 272334 389076 272340 389088
rect 3384 389048 272340 389076
rect 3384 389036 3390 389048
rect 272334 389036 272340 389048
rect 272392 389036 272398 389088
rect 4062 388968 4068 389020
rect 4120 389008 4126 389020
rect 273622 389008 273628 389020
rect 4120 388980 273628 389008
rect 4120 388968 4126 388980
rect 273622 388968 273628 388980
rect 273680 388968 273686 389020
rect 245470 388900 245476 388952
rect 245528 388940 245534 388952
rect 286410 388940 286416 388952
rect 245528 388912 286416 388940
rect 245528 388900 245534 388912
rect 286410 388900 286416 388912
rect 286468 388900 286474 388952
rect 239582 388832 239588 388884
rect 239640 388872 239646 388884
rect 286870 388872 286876 388884
rect 239640 388844 286876 388872
rect 239640 388832 239646 388844
rect 286870 388832 286876 388844
rect 286928 388832 286934 388884
rect 239214 388764 239220 388816
rect 239272 388804 239278 388816
rect 286686 388804 286692 388816
rect 239272 388776 286692 388804
rect 239272 388764 239278 388776
rect 286686 388764 286692 388776
rect 286744 388764 286750 388816
rect 3970 388696 3976 388748
rect 4028 388736 4034 388748
rect 273990 388736 273996 388748
rect 4028 388708 273996 388736
rect 4028 388696 4034 388708
rect 273990 388696 273996 388708
rect 274048 388696 274054 388748
rect 5258 388628 5264 388680
rect 5316 388668 5322 388680
rect 275278 388668 275284 388680
rect 5316 388640 275284 388668
rect 5316 388628 5322 388640
rect 275278 388628 275284 388640
rect 275336 388628 275342 388680
rect 3878 388560 3884 388612
rect 3936 388600 3942 388612
rect 274818 388600 274824 388612
rect 3936 388572 274824 388600
rect 3936 388560 3942 388572
rect 274818 388560 274824 388572
rect 274876 388560 274882 388612
rect 3786 388492 3792 388544
rect 3844 388532 3850 388544
rect 276106 388532 276112 388544
rect 3844 388504 276112 388532
rect 3844 388492 3850 388504
rect 276106 388492 276112 388504
rect 276164 388492 276170 388544
rect 3694 388424 3700 388476
rect 3752 388464 3758 388476
rect 277486 388464 277492 388476
rect 3752 388436 277492 388464
rect 3752 388424 3758 388436
rect 277486 388424 277492 388436
rect 277544 388424 277550 388476
rect 3602 388356 3608 388408
rect 3660 388396 3666 388408
rect 278774 388396 278780 388408
rect 3660 388368 278780 388396
rect 3660 388356 3666 388368
rect 278774 388356 278780 388368
rect 278832 388356 278838 388408
rect 3510 388288 3516 388340
rect 3568 388328 3574 388340
rect 279878 388328 279884 388340
rect 3568 388300 279884 388328
rect 3568 388288 3574 388300
rect 279878 388288 279884 388300
rect 279936 388288 279942 388340
rect 245562 388220 245568 388272
rect 245620 388260 245626 388272
rect 580166 388260 580172 388272
rect 245620 388232 580172 388260
rect 245620 388220 245626 388232
rect 580166 388220 580172 388232
rect 580224 388220 580230 388272
rect 244320 388152 244326 388204
rect 244378 388192 244384 388204
rect 249061 388195 249119 388201
rect 249061 388192 249073 388195
rect 244378 388164 249073 388192
rect 244378 388152 244384 388164
rect 249061 388161 249073 388164
rect 249107 388161 249119 388195
rect 249061 388155 249119 388161
rect 249150 388152 249156 388204
rect 249208 388192 249214 388204
rect 249518 388192 249524 388204
rect 249208 388164 249524 388192
rect 249208 388152 249214 388164
rect 249518 388152 249524 388164
rect 249576 388152 249582 388204
rect 249613 388195 249671 388201
rect 249613 388161 249625 388195
rect 249659 388192 249671 388195
rect 580902 388192 580908 388204
rect 249659 388164 580908 388192
rect 249659 388161 249671 388164
rect 249613 388155 249671 388161
rect 580902 388152 580908 388164
rect 580960 388152 580966 388204
rect 243952 388084 243958 388136
rect 244010 388124 244016 388136
rect 580810 388124 580816 388136
rect 244010 388096 580816 388124
rect 244010 388084 244016 388096
rect 580810 388084 580816 388096
rect 580868 388084 580874 388136
rect 242802 388016 242808 388068
rect 242860 388056 242866 388068
rect 580718 388056 580724 388068
rect 242860 388028 580724 388056
rect 242860 388016 242866 388028
rect 580718 388016 580724 388028
rect 580776 388016 580782 388068
rect 240410 387948 240416 388000
rect 240468 387988 240474 388000
rect 240468 387960 241192 387988
rect 240468 387948 240474 387960
rect 240870 387920 240876 387932
rect 240831 387892 240876 387920
rect 240870 387880 240876 387892
rect 240928 387880 240934 387932
rect 241164 387920 241192 387960
rect 241238 387948 241244 388000
rect 241296 387988 241302 388000
rect 580626 387988 580632 388000
rect 241296 387960 580632 387988
rect 241296 387948 241302 387960
rect 580626 387948 580632 387960
rect 580684 387948 580690 388000
rect 580534 387920 580540 387932
rect 241164 387892 580540 387920
rect 580534 387880 580540 387892
rect 580592 387880 580598 387932
rect 236730 387852 236736 387864
rect 236691 387824 236736 387852
rect 236730 387812 236736 387824
rect 236788 387812 236794 387864
rect 238386 387812 238392 387864
rect 238444 387852 238450 387864
rect 580442 387852 580448 387864
rect 238444 387824 580448 387852
rect 238444 387812 238450 387824
rect 580442 387812 580448 387824
rect 580500 387812 580506 387864
rect 287606 387132 287612 387184
rect 287664 387172 287670 387184
rect 294690 387172 294696 387184
rect 287664 387144 294696 387172
rect 287664 387132 287670 387144
rect 294690 387132 294696 387144
rect 294748 387132 294754 387184
rect 298738 386696 298744 386708
rect 277366 386668 298744 386696
rect 240873 386563 240931 386569
rect 240873 386529 240885 386563
rect 240919 386560 240931 386563
rect 277366 386560 277394 386668
rect 298738 386656 298744 386668
rect 298796 386656 298802 386708
rect 295978 386628 295984 386640
rect 240919 386532 277394 386560
rect 287440 386600 295984 386628
rect 240919 386529 240931 386532
rect 240873 386523 240931 386529
rect 234890 386452 234896 386504
rect 234948 386492 234954 386504
rect 287440 386492 287468 386600
rect 295978 386588 295984 386600
rect 296036 386588 296042 386640
rect 234948 386464 287468 386492
rect 234948 386452 234954 386464
rect 287606 386452 287612 386504
rect 287664 386492 287670 386504
rect 293402 386492 293408 386504
rect 287664 386464 293408 386492
rect 287664 386452 287670 386464
rect 293402 386452 293408 386464
rect 293460 386452 293466 386504
rect 236733 386427 236791 386433
rect 236733 386393 236745 386427
rect 236779 386424 236791 386427
rect 580258 386424 580264 386436
rect 236779 386396 580264 386424
rect 236779 386393 236791 386396
rect 236733 386387 236791 386393
rect 580258 386384 580264 386396
rect 580316 386384 580322 386436
rect 287514 385636 287520 385688
rect 287572 385676 287578 385688
rect 293494 385676 293500 385688
rect 287572 385648 293500 385676
rect 287572 385636 287578 385648
rect 293494 385636 293500 385648
rect 293552 385636 293558 385688
rect 287606 385364 287612 385416
rect 287664 385404 287670 385416
rect 293586 385404 293592 385416
rect 287664 385376 293592 385404
rect 287664 385364 287670 385376
rect 293586 385364 293592 385376
rect 293644 385364 293650 385416
rect 288342 385024 288348 385076
rect 288400 385064 288406 385076
rect 438118 385064 438124 385076
rect 288400 385036 438124 385064
rect 288400 385024 288406 385036
rect 438118 385024 438124 385036
rect 438176 385024 438182 385076
rect 288342 383664 288348 383716
rect 288400 383704 288406 383716
rect 299014 383704 299020 383716
rect 288400 383676 299020 383704
rect 288400 383664 288406 383676
rect 299014 383664 299020 383676
rect 299072 383664 299078 383716
rect 287606 382372 287612 382424
rect 287664 382412 287670 382424
rect 294874 382412 294880 382424
rect 287664 382384 294880 382412
rect 287664 382372 287670 382384
rect 294874 382372 294880 382384
rect 294932 382372 294938 382424
rect 288342 382304 288348 382356
rect 288400 382344 288406 382356
rect 294782 382344 294788 382356
rect 288400 382316 294788 382344
rect 288400 382304 288406 382316
rect 294782 382304 294788 382316
rect 294840 382304 294846 382356
rect 288158 380944 288164 380996
rect 288216 380984 288222 380996
rect 298922 380984 298928 380996
rect 288216 380956 298928 380984
rect 288216 380944 288222 380956
rect 298922 380944 298928 380956
rect 298980 380944 298986 380996
rect 288342 380876 288348 380928
rect 288400 380916 288406 380928
rect 537110 380916 537116 380928
rect 288400 380888 537116 380916
rect 288400 380876 288406 380888
rect 537110 380876 537116 380888
rect 537168 380876 537174 380928
rect 288342 379720 288348 379772
rect 288400 379760 288406 379772
rect 290826 379760 290832 379772
rect 288400 379732 290832 379760
rect 288400 379720 288406 379732
rect 290826 379720 290832 379732
rect 290884 379720 290890 379772
rect 288250 379516 288256 379568
rect 288308 379556 288314 379568
rect 370498 379556 370504 379568
rect 288308 379528 370504 379556
rect 288308 379516 288314 379528
rect 370498 379516 370504 379528
rect 370556 379516 370562 379568
rect 288342 378224 288348 378276
rect 288400 378264 288406 378276
rect 353938 378264 353944 378276
rect 288400 378236 353944 378264
rect 288400 378224 288406 378236
rect 353938 378224 353944 378236
rect 353996 378224 354002 378276
rect 288250 378156 288256 378208
rect 288308 378196 288314 378208
rect 356698 378196 356704 378208
rect 288308 378168 356704 378196
rect 288308 378156 288314 378168
rect 356698 378156 356704 378168
rect 356756 378156 356762 378208
rect 288342 376796 288348 376848
rect 288400 376836 288406 376848
rect 349798 376836 349804 376848
rect 288400 376808 349804 376836
rect 288400 376796 288406 376808
rect 349798 376796 349804 376808
rect 349856 376796 349862 376848
rect 288250 376728 288256 376780
rect 288308 376768 288314 376780
rect 352650 376768 352656 376780
rect 288308 376740 352656 376768
rect 288308 376728 288314 376740
rect 352650 376728 352656 376740
rect 352708 376728 352714 376780
rect 288158 375436 288164 375488
rect 288216 375476 288222 375488
rect 342898 375476 342904 375488
rect 288216 375448 342904 375476
rect 288216 375436 288222 375448
rect 342898 375436 342904 375448
rect 342956 375436 342962 375488
rect 288342 375368 288348 375420
rect 288400 375408 288406 375420
rect 345658 375408 345664 375420
rect 288400 375380 345664 375408
rect 288400 375368 288406 375380
rect 345658 375368 345664 375380
rect 345716 375368 345722 375420
rect 288158 374076 288164 374128
rect 288216 374116 288222 374128
rect 338758 374116 338764 374128
rect 288216 374088 338764 374116
rect 288216 374076 288222 374088
rect 338758 374076 338764 374088
rect 338816 374076 338822 374128
rect 288342 374008 288348 374060
rect 288400 374048 288406 374060
rect 340138 374048 340144 374060
rect 288400 374020 340144 374048
rect 288400 374008 288406 374020
rect 340138 374008 340144 374020
rect 340196 374008 340202 374060
rect 288342 372716 288348 372768
rect 288400 372756 288406 372768
rect 453298 372756 453304 372768
rect 288400 372728 453304 372756
rect 288400 372716 288406 372728
rect 453298 372716 453304 372728
rect 453356 372716 453362 372768
rect 288158 372648 288164 372700
rect 288216 372688 288222 372700
rect 454678 372688 454684 372700
rect 288216 372660 454684 372688
rect 288216 372648 288222 372660
rect 454678 372648 454684 372660
rect 454736 372648 454742 372700
rect 288250 372580 288256 372632
rect 288308 372620 288314 372632
rect 496814 372620 496820 372632
rect 288308 372592 496820 372620
rect 288308 372580 288314 372592
rect 496814 372580 496820 372592
rect 496872 372580 496878 372632
rect 288250 371220 288256 371272
rect 288308 371260 288314 371272
rect 450538 371260 450544 371272
rect 288308 371232 450544 371260
rect 288308 371220 288314 371232
rect 450538 371220 450544 371232
rect 450596 371220 450602 371272
rect 287606 369928 287612 369980
rect 287664 369968 287670 369980
rect 488534 369968 488540 369980
rect 287664 369940 488540 369968
rect 287664 369928 287670 369940
rect 488534 369928 488540 369940
rect 488592 369928 488598 369980
rect 288342 369860 288348 369912
rect 288400 369900 288406 369912
rect 489914 369900 489920 369912
rect 288400 369872 489920 369900
rect 288400 369860 288406 369872
rect 489914 369860 489920 369872
rect 489972 369860 489978 369912
rect 287606 368568 287612 368620
rect 287664 368608 287670 368620
rect 485038 368608 485044 368620
rect 287664 368580 485044 368608
rect 287664 368568 287670 368580
rect 485038 368568 485044 368580
rect 485096 368568 485102 368620
rect 288250 368500 288256 368552
rect 288308 368540 288314 368552
rect 486418 368540 486424 368552
rect 288308 368512 486424 368540
rect 288308 368500 288314 368512
rect 486418 368500 486424 368512
rect 486476 368500 486482 368552
rect 287974 367140 287980 367192
rect 288032 367180 288038 367192
rect 440970 367180 440976 367192
rect 288032 367152 440976 367180
rect 288032 367140 288038 367152
rect 440970 367140 440976 367152
rect 441028 367140 441034 367192
rect 288342 367072 288348 367124
rect 288400 367112 288406 367124
rect 440878 367112 440884 367124
rect 288400 367084 440884 367112
rect 288400 367072 288406 367084
rect 440878 367072 440884 367084
rect 440936 367072 440942 367124
rect 289078 365644 289084 365696
rect 289136 365684 289142 365696
rect 580166 365684 580172 365696
rect 289136 365656 580172 365684
rect 289136 365644 289142 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 288342 364352 288348 364404
rect 288400 364392 288406 364404
rect 478874 364392 478880 364404
rect 288400 364364 478880 364392
rect 288400 364352 288406 364364
rect 478874 364352 478880 364364
rect 478932 364352 478938 364404
rect 288158 362992 288164 363044
rect 288216 363032 288222 363044
rect 363598 363032 363604 363044
rect 288216 363004 363604 363032
rect 288216 362992 288222 363004
rect 363598 362992 363604 363004
rect 363656 362992 363662 363044
rect 287146 362924 287152 362976
rect 287204 362964 287210 362976
rect 367738 362964 367744 362976
rect 287204 362936 367744 362964
rect 287204 362924 287210 362936
rect 367738 362924 367744 362936
rect 367796 362924 367802 362976
rect 288250 361700 288256 361752
rect 288308 361740 288314 361752
rect 360838 361740 360844 361752
rect 288308 361712 360844 361740
rect 288308 361700 288314 361712
rect 360838 361700 360844 361712
rect 360896 361700 360902 361752
rect 288342 361632 288348 361684
rect 288400 361672 288406 361684
rect 472066 361672 472072 361684
rect 288400 361644 472072 361672
rect 288400 361632 288406 361644
rect 472066 361632 472072 361644
rect 472124 361632 472130 361684
rect 288158 361564 288164 361616
rect 288216 361604 288222 361616
rect 474734 361604 474740 361616
rect 288216 361576 474740 361604
rect 288216 361564 288222 361576
rect 474734 361564 474740 361576
rect 474792 361564 474798 361616
rect 288158 360272 288164 360324
rect 288216 360312 288222 360324
rect 359458 360312 359464 360324
rect 288216 360284 359464 360312
rect 288216 360272 288222 360284
rect 359458 360272 359464 360284
rect 359516 360272 359522 360324
rect 288342 360204 288348 360256
rect 288400 360244 288406 360256
rect 470594 360244 470600 360256
rect 288400 360216 470600 360244
rect 288400 360204 288406 360216
rect 470594 360204 470600 360216
rect 470652 360204 470658 360256
rect 288342 358776 288348 358828
rect 288400 358816 288406 358828
rect 449158 358816 449164 358828
rect 288400 358788 449164 358816
rect 288400 358776 288406 358788
rect 449158 358776 449164 358788
rect 449216 358776 449222 358828
rect 2774 358436 2780 358488
rect 2832 358476 2838 358488
rect 4706 358476 4712 358488
rect 2832 358448 4712 358476
rect 2832 358436 2838 358448
rect 4706 358436 4712 358448
rect 4764 358436 4770 358488
rect 288158 358300 288164 358352
rect 288216 358340 288222 358352
rect 467834 358340 467840 358352
rect 288216 358312 467840 358340
rect 288216 358300 288222 358312
rect 467834 358300 467840 358312
rect 467892 358300 467898 358352
rect 287330 358232 287336 358284
rect 287388 358272 287394 358284
rect 480254 358272 480260 358284
rect 287388 358244 480260 358272
rect 287388 358232 287394 358244
rect 480254 358232 480260 358244
rect 480312 358232 480318 358284
rect 287422 358164 287428 358216
rect 287480 358204 287486 358216
rect 481634 358204 481640 358216
rect 287480 358176 481640 358204
rect 287480 358164 287486 358176
rect 481634 358164 481640 358176
rect 481692 358164 481698 358216
rect 287514 358096 287520 358148
rect 287572 358136 287578 358148
rect 483014 358136 483020 358148
rect 287572 358108 483020 358136
rect 287572 358096 287578 358108
rect 483014 358096 483020 358108
rect 483072 358096 483078 358148
rect 287698 358028 287704 358080
rect 287756 358068 287762 358080
rect 491294 358068 491300 358080
rect 287756 358040 491300 358068
rect 287756 358028 287762 358040
rect 491294 358028 491300 358040
rect 491352 358028 491358 358080
rect 288250 357484 288256 357536
rect 288308 357524 288314 357536
rect 297450 357524 297456 357536
rect 288308 357496 297456 357524
rect 288308 357484 288314 357496
rect 297450 357484 297456 357496
rect 297508 357484 297514 357536
rect 288342 357416 288348 357468
rect 288400 357456 288406 357468
rect 297358 357456 297364 357468
rect 288400 357428 297364 357456
rect 288400 357416 288406 357428
rect 297358 357416 297364 357428
rect 297416 357416 297422 357468
rect 287606 356260 287612 356312
rect 287664 356300 287670 356312
rect 296254 356300 296260 356312
rect 287664 356272 296260 356300
rect 287664 356260 287670 356272
rect 296254 356260 296260 356272
rect 296312 356260 296318 356312
rect 287422 356056 287428 356108
rect 287480 356096 287486 356108
rect 296162 356096 296168 356108
rect 287480 356068 296168 356096
rect 287480 356056 287486 356068
rect 296162 356056 296168 356068
rect 296220 356056 296226 356108
rect 287974 354764 287980 354816
rect 288032 354804 288038 354816
rect 300210 354804 300216 354816
rect 288032 354776 300216 354804
rect 288032 354764 288038 354776
rect 300210 354764 300216 354776
rect 300268 354764 300274 354816
rect 288342 354696 288348 354748
rect 288400 354736 288406 354748
rect 438210 354736 438216 354748
rect 288400 354708 438216 354736
rect 288400 354696 288406 354708
rect 438210 354696 438216 354708
rect 438268 354696 438274 354748
rect 287606 353744 287612 353796
rect 287664 353784 287670 353796
rect 296346 353784 296352 353796
rect 287664 353756 296352 353784
rect 287664 353744 287670 353756
rect 296346 353744 296352 353756
rect 296404 353744 296410 353796
rect 286410 353200 286416 353252
rect 286468 353240 286474 353252
rect 580166 353240 580172 353252
rect 286468 353212 580172 353240
rect 286468 353200 286474 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 288342 351908 288348 351960
rect 288400 351948 288406 351960
rect 300394 351948 300400 351960
rect 288400 351920 300400 351948
rect 288400 351908 288406 351920
rect 300394 351908 300400 351920
rect 300452 351908 300458 351960
rect 288342 350616 288348 350668
rect 288400 350656 288406 350668
rect 300302 350656 300308 350668
rect 288400 350628 300308 350656
rect 288400 350616 288406 350628
rect 300302 350616 300308 350628
rect 300360 350616 300366 350668
rect 288066 350548 288072 350600
rect 288124 350588 288130 350600
rect 439682 350588 439688 350600
rect 288124 350560 439688 350588
rect 288124 350548 288130 350560
rect 439682 350548 439688 350560
rect 439740 350548 439746 350600
rect 287698 350276 287704 350328
rect 287756 350316 287762 350328
rect 287974 350316 287980 350328
rect 287756 350288 287980 350316
rect 287756 350276 287762 350288
rect 287974 350276 287980 350288
rect 288032 350276 288038 350328
rect 288250 349256 288256 349308
rect 288308 349296 288314 349308
rect 296438 349296 296444 349308
rect 288308 349268 296444 349296
rect 288308 349256 288314 349268
rect 296438 349256 296444 349268
rect 296496 349256 296502 349308
rect 288342 349120 288348 349172
rect 288400 349160 288406 349172
rect 300486 349160 300492 349172
rect 288400 349132 300492 349160
rect 288400 349120 288406 349132
rect 300486 349120 300492 349132
rect 300544 349120 300550 349172
rect 288250 347896 288256 347948
rect 288308 347936 288314 347948
rect 296530 347936 296536 347948
rect 288308 347908 296536 347936
rect 288308 347896 288314 347908
rect 296530 347896 296536 347908
rect 296588 347896 296594 347948
rect 288342 347760 288348 347812
rect 288400 347800 288406 347812
rect 299106 347800 299112 347812
rect 288400 347772 299112 347800
rect 288400 347760 288406 347772
rect 299106 347760 299112 347772
rect 299164 347760 299170 347812
rect 288342 346672 288348 346724
rect 288400 346712 288406 346724
rect 294966 346712 294972 346724
rect 288400 346684 294972 346712
rect 288400 346672 288406 346684
rect 294966 346672 294972 346684
rect 295024 346672 295030 346724
rect 287606 346400 287612 346452
rect 287664 346440 287670 346452
rect 295058 346440 295064 346452
rect 287664 346412 295064 346440
rect 287664 346400 287670 346412
rect 295058 346400 295064 346412
rect 295116 346400 295122 346452
rect 2774 345856 2780 345908
rect 2832 345896 2838 345908
rect 5442 345896 5448 345908
rect 2832 345868 5448 345896
rect 2832 345856 2838 345868
rect 5442 345856 5448 345868
rect 5500 345856 5506 345908
rect 287330 345108 287336 345160
rect 287388 345148 287394 345160
rect 299290 345148 299296 345160
rect 287388 345120 299296 345148
rect 287388 345108 287394 345120
rect 299290 345108 299296 345120
rect 299348 345108 299354 345160
rect 288342 345040 288348 345092
rect 288400 345080 288406 345092
rect 352558 345080 352564 345092
rect 288400 345052 352564 345080
rect 288400 345040 288406 345052
rect 352558 345040 352564 345052
rect 352616 345040 352622 345092
rect 288158 343680 288164 343732
rect 288216 343720 288222 343732
rect 295150 343720 295156 343732
rect 288216 343692 295156 343720
rect 288216 343680 288222 343692
rect 295150 343680 295156 343692
rect 295208 343680 295214 343732
rect 288342 342252 288348 342304
rect 288400 342292 288406 342304
rect 299198 342292 299204 342304
rect 288400 342264 299204 342292
rect 288400 342252 288406 342264
rect 299198 342252 299204 342264
rect 299256 342252 299262 342304
rect 288342 340960 288348 341012
rect 288400 341000 288406 341012
rect 297634 341000 297640 341012
rect 288400 340972 297640 341000
rect 288400 340960 288406 340972
rect 297634 340960 297640 340972
rect 297692 340960 297698 341012
rect 287698 340892 287704 340944
rect 287756 340932 287762 340944
rect 297542 340932 297548 340944
rect 287756 340904 297548 340932
rect 287756 340892 287762 340904
rect 297542 340892 297548 340904
rect 297600 340892 297606 340944
rect 288342 339532 288348 339584
rect 288400 339572 288406 339584
rect 296622 339572 296628 339584
rect 288400 339544 296628 339572
rect 288400 339532 288406 339544
rect 296622 339532 296628 339544
rect 296680 339532 296686 339584
rect 288250 339464 288256 339516
rect 288308 339504 288314 339516
rect 297726 339504 297732 339516
rect 288308 339476 297732 339504
rect 288308 339464 288314 339476
rect 297726 339464 297732 339476
rect 297784 339464 297790 339516
rect 288250 338172 288256 338224
rect 288308 338212 288314 338224
rect 300578 338212 300584 338224
rect 288308 338184 300584 338212
rect 288308 338172 288314 338184
rect 300578 338172 300584 338184
rect 300636 338172 300642 338224
rect 269712 338104 269718 338156
rect 269770 338144 269776 338156
rect 282457 338147 282515 338153
rect 282457 338144 282469 338147
rect 269770 338116 282469 338144
rect 269770 338104 269776 338116
rect 282457 338113 282469 338116
rect 282503 338113 282515 338147
rect 282457 338107 282515 338113
rect 288342 338104 288348 338156
rect 288400 338144 288406 338156
rect 439774 338144 439780 338156
rect 288400 338116 439780 338144
rect 288400 338104 288406 338116
rect 439774 338104 439780 338116
rect 439832 338104 439838 338156
rect 279605 338079 279663 338085
rect 279605 338045 279617 338079
rect 279651 338076 279663 338079
rect 282641 338079 282699 338085
rect 282641 338076 282653 338079
rect 279651 338048 282653 338076
rect 279651 338045 279663 338048
rect 279605 338039 279663 338045
rect 282641 338045 282653 338048
rect 282687 338045 282699 338079
rect 282641 338039 282699 338045
rect 235077 338011 235135 338017
rect 235077 337977 235089 338011
rect 235123 338008 235135 338011
rect 250533 338011 250591 338017
rect 235123 337980 238662 338008
rect 235123 337977 235135 337980
rect 235077 337971 235135 337977
rect 238634 337952 238662 337980
rect 250533 337977 250545 338011
rect 250579 338008 250591 338011
rect 274545 338011 274603 338017
rect 274545 338008 274557 338011
rect 250579 337980 250806 338008
rect 250579 337977 250591 337980
rect 250533 337971 250591 337977
rect 250778 337952 250806 337980
rect 270650 337980 274557 338008
rect 270650 337952 270678 337980
rect 274545 337977 274557 337980
rect 274591 337977 274603 338011
rect 274545 337971 274603 337977
rect 234798 337900 234804 337952
rect 234856 337940 234862 337952
rect 235212 337940 235218 337952
rect 234856 337912 235218 337940
rect 234856 337900 234862 337912
rect 235212 337900 235218 337912
rect 235270 337900 235276 337952
rect 235672 337900 235678 337952
rect 235730 337900 235736 337952
rect 235948 337940 235954 337952
rect 235920 337900 235954 337940
rect 236006 337900 236012 337952
rect 236500 337900 236506 337952
rect 236558 337900 236564 337952
rect 237512 337900 237518 337952
rect 237570 337900 237576 337952
rect 237604 337900 237610 337952
rect 237662 337940 237668 337952
rect 237662 337912 238432 337940
rect 237662 337900 237668 337912
rect 234982 337832 234988 337884
rect 235040 337872 235046 337884
rect 235690 337872 235718 337900
rect 235040 337844 235718 337872
rect 235040 337832 235046 337844
rect 235810 337628 235816 337680
rect 235868 337668 235874 337680
rect 235920 337668 235948 337900
rect 235868 337640 235948 337668
rect 235868 337628 235874 337640
rect 236518 337544 236546 337900
rect 236641 337875 236699 337881
rect 236641 337841 236653 337875
rect 236687 337872 236699 337875
rect 236776 337872 236782 337884
rect 236687 337844 236782 337872
rect 236687 337841 236699 337844
rect 236641 337835 236699 337841
rect 236776 337832 236782 337844
rect 236834 337832 236840 337884
rect 236960 337832 236966 337884
rect 237018 337832 237024 337884
rect 236978 337680 237006 337832
rect 237530 337736 237558 337900
rect 237880 337881 237886 337884
rect 237837 337875 237886 337881
rect 237837 337841 237849 337875
rect 237883 337841 237886 337875
rect 237837 337835 237886 337841
rect 237880 337832 237886 337835
rect 237938 337832 237944 337884
rect 237972 337804 237978 337816
rect 237944 337764 237978 337804
rect 238030 337764 238036 337816
rect 237530 337708 237696 337736
rect 237668 337680 237696 337708
rect 236914 337628 236920 337680
rect 236972 337640 237006 337680
rect 236972 337628 236978 337640
rect 237650 337628 237656 337680
rect 237708 337628 237714 337680
rect 237944 337612 237972 337764
rect 238404 337680 238432 337912
rect 238616 337900 238622 337952
rect 238674 337900 238680 337952
rect 238800 337949 238806 337952
rect 238757 337943 238806 337949
rect 238757 337909 238769 337943
rect 238803 337909 238806 337943
rect 238757 337903 238806 337909
rect 238800 337900 238806 337903
rect 238858 337900 238864 337952
rect 238892 337900 238898 337952
rect 238950 337900 238956 337952
rect 239444 337900 239450 337952
rect 239502 337900 239508 337952
rect 240456 337949 240462 337952
rect 240413 337943 240462 337949
rect 240413 337909 240425 337943
rect 240459 337909 240462 337943
rect 240413 337903 240462 337909
rect 240456 337900 240462 337903
rect 240514 337900 240520 337952
rect 241744 337900 241750 337952
rect 241802 337900 241808 337952
rect 242112 337900 242118 337952
rect 242170 337900 242176 337952
rect 242345 337943 242403 337949
rect 242345 337909 242357 337943
rect 242391 337940 242403 337943
rect 242664 337940 242670 337952
rect 242391 337912 242670 337940
rect 242391 337909 242403 337912
rect 242345 337903 242403 337909
rect 242664 337900 242670 337912
rect 242722 337900 242728 337952
rect 242848 337949 242854 337952
rect 242805 337943 242854 337949
rect 242805 337909 242817 337943
rect 242851 337909 242854 337943
rect 242805 337903 242854 337909
rect 242848 337900 242854 337903
rect 242906 337900 242912 337952
rect 243308 337949 243314 337952
rect 243265 337943 243314 337949
rect 243265 337909 243277 337943
rect 243311 337909 243314 337943
rect 243265 337903 243314 337909
rect 243308 337900 243314 337903
rect 243366 337900 243372 337952
rect 243492 337949 243498 337952
rect 243449 337943 243498 337949
rect 243449 337909 243461 337943
rect 243495 337909 243498 337943
rect 243449 337903 243498 337909
rect 243492 337900 243498 337903
rect 243550 337900 243556 337952
rect 243768 337949 243774 337952
rect 243725 337943 243774 337949
rect 243725 337909 243737 337943
rect 243771 337909 243774 337943
rect 243725 337903 243774 337909
rect 243768 337900 243774 337903
rect 243826 337900 243832 337952
rect 244504 337900 244510 337952
rect 244562 337900 244568 337952
rect 245056 337949 245062 337952
rect 245013 337943 245062 337949
rect 245013 337909 245025 337943
rect 245059 337909 245062 337943
rect 245013 337903 245062 337909
rect 245056 337900 245062 337903
rect 245114 337900 245120 337952
rect 245148 337900 245154 337952
rect 245206 337949 245212 337952
rect 245332 337949 245338 337952
rect 245206 337943 245255 337949
rect 245206 337909 245209 337943
rect 245243 337909 245255 337943
rect 245206 337903 245255 337909
rect 245289 337943 245338 337949
rect 245289 337909 245301 337943
rect 245335 337909 245338 337943
rect 245289 337903 245338 337909
rect 245206 337900 245212 337903
rect 245332 337900 245338 337903
rect 245390 337900 245396 337952
rect 245933 337943 245991 337949
rect 245933 337909 245945 337943
rect 245979 337940 245991 337943
rect 247356 337940 247362 337952
rect 245979 337912 247362 337940
rect 245979 337909 245991 337912
rect 245933 337903 245991 337909
rect 247356 337900 247362 337912
rect 247414 337900 247420 337952
rect 248184 337900 248190 337952
rect 248242 337900 248248 337952
rect 249748 337949 249754 337952
rect 249705 337943 249754 337949
rect 249705 337909 249717 337943
rect 249751 337909 249754 337943
rect 249705 337903 249754 337909
rect 249748 337900 249754 337903
rect 249806 337900 249812 337952
rect 249840 337900 249846 337952
rect 249898 337949 249904 337952
rect 249898 337943 249947 337949
rect 249898 337909 249901 337943
rect 249935 337909 249947 337943
rect 249898 337903 249947 337909
rect 249898 337900 249904 337903
rect 250760 337900 250766 337952
rect 250818 337900 250824 337952
rect 250852 337900 250858 337952
rect 250910 337900 250916 337952
rect 251496 337900 251502 337952
rect 251554 337949 251560 337952
rect 251554 337943 251603 337949
rect 251554 337909 251557 337943
rect 251591 337909 251603 337943
rect 251554 337903 251603 337909
rect 252189 337943 252247 337949
rect 252189 337909 252201 337943
rect 252235 337940 252247 337943
rect 252600 337940 252606 337952
rect 252235 337912 252606 337940
rect 252235 337909 252247 337912
rect 252189 337903 252247 337909
rect 251554 337900 251560 337903
rect 252600 337900 252606 337912
rect 252658 337900 252664 337952
rect 254256 337949 254262 337952
rect 254213 337943 254262 337949
rect 254213 337909 254225 337943
rect 254259 337909 254262 337943
rect 254213 337903 254262 337909
rect 254256 337900 254262 337903
rect 254314 337900 254320 337952
rect 254900 337900 254906 337952
rect 254958 337900 254964 337952
rect 255084 337900 255090 337952
rect 255142 337900 255148 337952
rect 256188 337900 256194 337952
rect 256246 337900 256252 337952
rect 257157 337943 257215 337949
rect 257157 337909 257169 337943
rect 257203 337940 257215 337943
rect 257384 337940 257390 337952
rect 257203 337912 257390 337940
rect 257203 337909 257215 337912
rect 257157 337903 257215 337909
rect 257384 337900 257390 337912
rect 257442 337900 257448 337952
rect 257568 337949 257574 337952
rect 257525 337943 257574 337949
rect 257525 337909 257537 337943
rect 257571 337909 257574 337943
rect 257525 337903 257574 337909
rect 257568 337900 257574 337903
rect 257626 337900 257632 337952
rect 257752 337949 257758 337952
rect 257709 337943 257758 337949
rect 257709 337909 257721 337943
rect 257755 337909 257758 337943
rect 257709 337903 257758 337909
rect 257752 337900 257758 337903
rect 257810 337900 257816 337952
rect 257844 337900 257850 337952
rect 257902 337900 257908 337952
rect 258856 337900 258862 337952
rect 258914 337900 258920 337952
rect 259132 337900 259138 337952
rect 259190 337940 259196 337952
rect 259273 337943 259331 337949
rect 259273 337940 259285 337943
rect 259190 337912 259285 337940
rect 259190 337900 259196 337912
rect 259273 337909 259285 337912
rect 259319 337909 259331 337943
rect 259273 337903 259331 337909
rect 260144 337900 260150 337952
rect 260202 337900 260208 337952
rect 260236 337900 260242 337952
rect 260294 337940 260300 337952
rect 260561 337943 260619 337949
rect 260561 337940 260573 337943
rect 260294 337912 260573 337940
rect 260294 337900 260300 337912
rect 260561 337909 260573 337912
rect 260607 337909 260619 337943
rect 260561 337903 260619 337909
rect 261800 337900 261806 337952
rect 261858 337949 261864 337952
rect 261858 337943 261907 337949
rect 261858 337909 261861 337943
rect 261895 337909 261907 337943
rect 261858 337903 261907 337909
rect 261858 337900 261864 337903
rect 261984 337900 261990 337952
rect 262042 337940 262048 337952
rect 263321 337943 263379 337949
rect 263321 337940 263333 337943
rect 262042 337912 263333 337940
rect 262042 337900 262048 337912
rect 263321 337909 263333 337912
rect 263367 337909 263379 337943
rect 263321 337903 263379 337909
rect 263640 337900 263646 337952
rect 263698 337900 263704 337952
rect 264928 337900 264934 337952
rect 264986 337940 264992 337952
rect 266633 337943 266691 337949
rect 266633 337940 266645 337943
rect 264986 337912 266645 337940
rect 264986 337900 264992 337912
rect 266633 337909 266645 337912
rect 266679 337909 266691 337943
rect 266633 337903 266691 337909
rect 267228 337900 267234 337952
rect 267286 337900 267292 337952
rect 267320 337900 267326 337952
rect 267378 337949 267384 337952
rect 267378 337943 267427 337949
rect 267378 337909 267381 337943
rect 267415 337909 267427 337943
rect 267378 337903 267427 337909
rect 268105 337943 268163 337949
rect 268105 337909 268117 337943
rect 268151 337940 268163 337943
rect 268240 337940 268246 337952
rect 268151 337912 268246 337940
rect 268151 337909 268163 337912
rect 268105 337903 268163 337909
rect 267378 337900 267384 337903
rect 268240 337900 268246 337912
rect 268298 337900 268304 337952
rect 269988 337900 269994 337952
rect 270046 337949 270052 337952
rect 270046 337943 270095 337949
rect 270046 337909 270049 337943
rect 270083 337909 270095 337943
rect 270046 337903 270095 337909
rect 270046 337900 270052 337903
rect 270172 337900 270178 337952
rect 270230 337940 270236 337952
rect 270405 337943 270463 337949
rect 270405 337940 270417 337943
rect 270230 337912 270417 337940
rect 270230 337900 270236 337912
rect 270405 337909 270417 337912
rect 270451 337909 270463 337943
rect 270405 337903 270463 337909
rect 270632 337900 270638 337952
rect 270690 337900 270696 337952
rect 270724 337900 270730 337952
rect 270782 337940 270788 337952
rect 271049 337943 271107 337949
rect 271049 337940 271061 337943
rect 270782 337912 271061 337940
rect 270782 337900 270788 337912
rect 271049 337909 271061 337912
rect 271095 337909 271107 337943
rect 271049 337903 271107 337909
rect 271276 337900 271282 337952
rect 271334 337900 271340 337952
rect 271368 337900 271374 337952
rect 271426 337949 271432 337952
rect 271426 337943 271475 337949
rect 271426 337909 271429 337943
rect 271463 337909 271475 337943
rect 271426 337903 271475 337909
rect 271426 337900 271432 337903
rect 272656 337900 272662 337952
rect 272714 337940 272720 337952
rect 272797 337943 272855 337949
rect 272797 337940 272809 337943
rect 272714 337912 272809 337940
rect 272714 337900 272720 337912
rect 272797 337909 272809 337912
rect 272843 337909 272855 337943
rect 274085 337943 274143 337949
rect 274085 337940 274097 337943
rect 272797 337903 272855 337909
rect 272904 337912 274097 337940
rect 238910 337816 238938 337900
rect 239168 337832 239174 337884
rect 239226 337832 239232 337884
rect 238846 337764 238852 337816
rect 238904 337776 238938 337816
rect 238904 337764 238910 337776
rect 238386 337628 238392 337680
rect 238444 337628 238450 337680
rect 239030 337628 239036 337680
rect 239088 337668 239094 337680
rect 239186 337668 239214 337832
rect 239462 337816 239490 337900
rect 240689 337875 240747 337881
rect 240689 337841 240701 337875
rect 240735 337872 240747 337875
rect 241100 337872 241106 337884
rect 240735 337844 241106 337872
rect 240735 337841 240747 337844
rect 240689 337835 240747 337841
rect 241100 337832 241106 337844
rect 241158 337832 241164 337884
rect 241468 337832 241474 337884
rect 241526 337832 241532 337884
rect 239462 337776 239496 337816
rect 239490 337764 239496 337776
rect 239548 337764 239554 337816
rect 240548 337764 240554 337816
rect 240606 337804 240612 337816
rect 240965 337807 241023 337813
rect 240965 337804 240977 337807
rect 240606 337776 240977 337804
rect 240606 337764 240612 337776
rect 240965 337773 240977 337776
rect 241011 337773 241023 337807
rect 240965 337767 241023 337773
rect 240870 337736 240876 337748
rect 240831 337708 240876 337736
rect 240870 337696 240876 337708
rect 240928 337696 240934 337748
rect 239088 337640 239214 337668
rect 239088 337628 239094 337640
rect 240502 337628 240508 337680
rect 240560 337668 240566 337680
rect 241486 337668 241514 337832
rect 241762 337680 241790 337900
rect 240560 337640 241514 337668
rect 240560 337628 240566 337640
rect 241698 337628 241704 337680
rect 241756 337640 241790 337680
rect 241756 337628 241762 337640
rect 237926 337560 237932 337612
rect 237984 337560 237990 337612
rect 236454 337492 236460 337544
rect 236512 337504 236546 337544
rect 240686 337532 240692 337544
rect 240647 337504 240692 337532
rect 236512 337492 236518 337504
rect 240686 337492 240692 337504
rect 240744 337492 240750 337544
rect 241514 337492 241520 337544
rect 241572 337532 241578 337544
rect 242130 337532 242158 337900
rect 242480 337832 242486 337884
rect 242538 337872 242544 337884
rect 242538 337832 242572 337872
rect 243170 337832 243176 337884
rect 243228 337832 243234 337884
rect 243952 337832 243958 337884
rect 244010 337832 244016 337884
rect 244228 337832 244234 337884
rect 244286 337832 244292 337884
rect 242296 337764 242302 337816
rect 242354 337764 242360 337816
rect 242314 337736 242342 337764
rect 242268 337708 242342 337736
rect 242268 337680 242296 337708
rect 242544 337680 242572 337832
rect 242621 337807 242679 337813
rect 242621 337773 242633 337807
rect 242667 337804 242679 337807
rect 242940 337804 242946 337816
rect 242667 337776 242946 337804
rect 242667 337773 242679 337776
rect 242621 337767 242679 337773
rect 242940 337764 242946 337776
rect 242998 337764 243004 337816
rect 243188 337736 243216 337832
rect 243400 337813 243406 337816
rect 243357 337807 243406 337813
rect 243357 337773 243369 337807
rect 243403 337773 243406 337807
rect 243357 337767 243406 337773
rect 243400 337764 243406 337767
rect 243458 337764 243464 337816
rect 243188 337708 243492 337736
rect 243464 337680 243492 337708
rect 243970 337680 243998 337832
rect 242250 337628 242256 337680
rect 242308 337628 242314 337680
rect 242526 337628 242532 337680
rect 242584 337628 242590 337680
rect 243446 337628 243452 337680
rect 243504 337628 243510 337680
rect 243906 337628 243912 337680
rect 243964 337640 243998 337680
rect 243964 337628 243970 337640
rect 244090 337628 244096 337680
rect 244148 337668 244154 337680
rect 244246 337668 244274 337832
rect 244522 337736 244550 337900
rect 244688 337832 244694 337884
rect 244746 337832 244752 337884
rect 244872 337832 244878 337884
rect 244930 337881 244936 337884
rect 244930 337875 244979 337881
rect 244930 337841 244933 337875
rect 244967 337841 244979 337875
rect 244930 337835 244979 337841
rect 244930 337832 244936 337835
rect 246344 337832 246350 337884
rect 246402 337832 246408 337884
rect 246528 337832 246534 337884
rect 246586 337832 246592 337884
rect 247264 337881 247270 337884
rect 247221 337875 247270 337881
rect 247221 337841 247233 337875
rect 247267 337841 247270 337875
rect 247221 337835 247270 337841
rect 247264 337832 247270 337835
rect 247322 337832 247328 337884
rect 247448 337832 247454 337884
rect 247506 337832 247512 337884
rect 247770 337832 247776 337884
rect 247828 337832 247834 337884
rect 248092 337881 248098 337884
rect 248049 337875 248098 337881
rect 248049 337841 248061 337875
rect 248095 337841 248098 337875
rect 248049 337835 248098 337841
rect 248092 337832 248098 337835
rect 248150 337832 248156 337884
rect 244522 337708 244596 337736
rect 244568 337680 244596 337708
rect 244706 337680 244734 337832
rect 244780 337764 244786 337816
rect 244838 337804 244844 337816
rect 245470 337804 245476 337816
rect 244838 337764 244872 337804
rect 245431 337776 245476 337804
rect 245470 337764 245476 337776
rect 245528 337764 245534 337816
rect 245608 337813 245614 337816
rect 245565 337807 245614 337813
rect 245565 337773 245577 337807
rect 245611 337773 245614 337807
rect 245565 337767 245614 337773
rect 245608 337764 245614 337767
rect 245666 337764 245672 337816
rect 245792 337764 245798 337816
rect 245850 337813 245856 337816
rect 245850 337807 245899 337813
rect 245850 337773 245853 337807
rect 245887 337773 245899 337807
rect 245850 337767 245899 337773
rect 245850 337764 245856 337767
rect 244844 337680 244872 337764
rect 246362 337680 246390 337832
rect 246546 337680 246574 337832
rect 247080 337764 247086 337816
rect 247138 337764 247144 337816
rect 247098 337736 247126 337764
rect 247052 337708 247126 337736
rect 247052 337680 247080 337708
rect 244148 337640 244274 337668
rect 244148 337628 244154 337640
rect 244550 337628 244556 337680
rect 244608 337628 244614 337680
rect 244706 337640 244740 337680
rect 244734 337628 244740 337640
rect 244792 337628 244798 337680
rect 244826 337628 244832 337680
rect 244884 337628 244890 337680
rect 246362 337640 246396 337680
rect 246390 337628 246396 337640
rect 246448 337628 246454 337680
rect 246482 337628 246488 337680
rect 246540 337640 246574 337680
rect 246540 337628 246546 337640
rect 247034 337628 247040 337680
rect 247092 337628 247098 337680
rect 247310 337628 247316 337680
rect 247368 337668 247374 337680
rect 247466 337668 247494 337832
rect 247632 337813 247638 337816
rect 247589 337807 247638 337813
rect 247589 337773 247601 337807
rect 247635 337773 247638 337807
rect 247589 337767 247638 337773
rect 247632 337764 247638 337767
rect 247690 337764 247696 337816
rect 247788 337736 247816 337832
rect 248202 337804 248230 337900
rect 248368 337872 248374 337884
rect 248156 337776 248230 337804
rect 248340 337832 248374 337872
rect 248426 337832 248432 337884
rect 248552 337832 248558 337884
rect 248610 337832 248616 337884
rect 250392 337881 250398 337884
rect 250349 337875 250398 337881
rect 250349 337841 250361 337875
rect 250395 337841 250398 337875
rect 250349 337835 250398 337841
rect 250392 337832 250398 337835
rect 250450 337832 250456 337884
rect 247788 337708 248000 337736
rect 247972 337680 248000 337708
rect 247368 337640 247494 337668
rect 247368 337628 247374 337640
rect 247954 337628 247960 337680
rect 248012 337628 248018 337680
rect 248156 337612 248184 337776
rect 248340 337748 248368 337832
rect 248322 337696 248328 337748
rect 248380 337696 248386 337748
rect 248570 337736 248598 337832
rect 250870 337816 250898 337900
rect 251036 337832 251042 337884
rect 251094 337832 251100 337884
rect 251680 337832 251686 337884
rect 251738 337881 251744 337884
rect 251738 337875 251787 337881
rect 251738 337841 251741 337875
rect 251775 337841 251787 337875
rect 252048 337872 252054 337884
rect 251738 337835 251787 337841
rect 251836 337844 252054 337872
rect 251738 337832 251744 337835
rect 250208 337764 250214 337816
rect 250266 337804 250272 337816
rect 250266 337764 250300 337804
rect 250806 337764 250812 337816
rect 250864 337776 250898 337816
rect 250864 337764 250870 337776
rect 250070 337736 250076 337748
rect 248432 337708 248598 337736
rect 250031 337708 250076 337736
rect 248432 337680 248460 337708
rect 250070 337696 250076 337708
rect 250128 337696 250134 337748
rect 250272 337680 250300 337764
rect 248414 337628 248420 337680
rect 248472 337628 248478 337680
rect 250254 337628 250260 337680
rect 250312 337628 250318 337680
rect 242802 337600 242808 337612
rect 242763 337572 242808 337600
rect 242802 337560 242808 337572
rect 242860 337560 242866 337612
rect 245194 337600 245200 337612
rect 245155 337572 245200 337600
rect 245194 337560 245200 337572
rect 245252 337560 245258 337612
rect 248138 337560 248144 337612
rect 248196 337560 248202 337612
rect 250070 337560 250076 337612
rect 250128 337600 250134 337612
rect 251054 337600 251082 337832
rect 251266 337736 251272 337748
rect 251227 337708 251272 337736
rect 251266 337696 251272 337708
rect 251324 337696 251330 337748
rect 251836 337612 251864 337844
rect 252048 337832 252054 337844
rect 252106 337832 252112 337884
rect 252784 337881 252790 337884
rect 252741 337875 252790 337881
rect 252741 337841 252753 337875
rect 252787 337841 252790 337875
rect 252741 337835 252790 337841
rect 252784 337832 252790 337835
rect 252842 337832 252848 337884
rect 253060 337881 253066 337884
rect 253017 337875 253066 337881
rect 253017 337841 253029 337875
rect 253063 337841 253066 337875
rect 253017 337835 253066 337841
rect 253060 337832 253066 337835
rect 253118 337832 253124 337884
rect 253336 337832 253342 337884
rect 253394 337832 253400 337884
rect 254440 337872 254446 337884
rect 254412 337832 254446 337872
rect 254498 337832 254504 337884
rect 253198 337628 253204 337680
rect 253256 337668 253262 337680
rect 253354 337668 253382 337832
rect 253477 337807 253535 337813
rect 253477 337773 253489 337807
rect 253523 337804 253535 337807
rect 254072 337804 254078 337816
rect 253523 337776 254078 337804
rect 253523 337773 253535 337776
rect 253477 337767 253535 337773
rect 254072 337764 254078 337776
rect 254130 337764 254136 337816
rect 254412 337680 254440 337832
rect 254918 337736 254946 337900
rect 254918 337708 254992 337736
rect 254964 337680 254992 337708
rect 255102 337680 255130 337900
rect 255360 337832 255366 337884
rect 255418 337832 255424 337884
rect 255452 337832 255458 337884
rect 255510 337881 255516 337884
rect 255510 337875 255559 337881
rect 255510 337841 255513 337875
rect 255547 337841 255559 337875
rect 255510 337835 255559 337841
rect 255593 337875 255651 337881
rect 255593 337841 255605 337875
rect 255639 337872 255651 337875
rect 255820 337872 255826 337884
rect 255639 337844 255826 337872
rect 255639 337841 255651 337844
rect 255593 337835 255651 337841
rect 255510 337832 255516 337835
rect 255820 337832 255826 337844
rect 255878 337832 255884 337884
rect 256096 337832 256102 337884
rect 256154 337832 256160 337884
rect 253256 337640 253382 337668
rect 253256 337628 253262 337640
rect 254394 337628 254400 337680
rect 254452 337628 254458 337680
rect 254946 337628 254952 337680
rect 255004 337628 255010 337680
rect 255038 337628 255044 337680
rect 255096 337640 255130 337680
rect 255096 337628 255102 337640
rect 250128 337572 251082 337600
rect 250128 337560 250134 337572
rect 251818 337560 251824 337612
rect 251876 337560 251882 337612
rect 255378 337600 255406 337832
rect 255774 337600 255780 337612
rect 255378 337572 255780 337600
rect 255774 337560 255780 337572
rect 255832 337560 255838 337612
rect 241572 337504 242158 337532
rect 251545 337535 251603 337541
rect 241572 337492 241578 337504
rect 251545 337501 251557 337535
rect 251591 337532 251603 337535
rect 251634 337532 251640 337544
rect 251591 337504 251640 337532
rect 251591 337501 251603 337504
rect 251545 337495 251603 337501
rect 251634 337492 251640 337504
rect 251692 337492 251698 337544
rect 255590 337532 255596 337544
rect 255551 337504 255596 337532
rect 255590 337492 255596 337504
rect 255648 337492 255654 337544
rect 255866 337492 255872 337544
rect 255924 337532 255930 337544
rect 256114 337532 256142 337832
rect 255924 337504 256142 337532
rect 256206 337544 256234 337900
rect 257862 337872 257890 337900
rect 257816 337844 257890 337872
rect 257476 337764 257482 337816
rect 257534 337804 257540 337816
rect 257617 337807 257675 337813
rect 257617 337804 257629 337807
rect 257534 337776 257629 337804
rect 257534 337764 257540 337776
rect 257617 337773 257629 337776
rect 257663 337773 257675 337807
rect 257617 337767 257675 337773
rect 257816 337748 257844 337844
rect 258028 337832 258034 337884
rect 258086 337881 258092 337884
rect 258086 337875 258135 337881
rect 258086 337841 258089 337875
rect 258123 337841 258135 337875
rect 258086 337835 258135 337841
rect 258086 337832 258092 337835
rect 258580 337832 258586 337884
rect 258638 337832 258644 337884
rect 257798 337696 257804 337748
rect 257856 337696 257862 337748
rect 257525 337671 257583 337677
rect 257525 337637 257537 337671
rect 257571 337668 257583 337671
rect 257614 337668 257620 337680
rect 257571 337640 257620 337668
rect 257571 337637 257583 337640
rect 257525 337631 257583 337637
rect 257614 337628 257620 337640
rect 257672 337628 257678 337680
rect 257154 337600 257160 337612
rect 257115 337572 257160 337600
rect 257154 337560 257160 337572
rect 257212 337560 257218 337612
rect 258598 337600 258626 337832
rect 258874 337668 258902 337900
rect 259868 337832 259874 337884
rect 259926 337832 259932 337884
rect 260052 337832 260058 337884
rect 260110 337832 260116 337884
rect 260162 337872 260190 337900
rect 260469 337875 260527 337881
rect 260469 337872 260481 337875
rect 260162 337844 260481 337872
rect 260469 337841 260481 337844
rect 260515 337841 260527 337875
rect 260469 337835 260527 337841
rect 260880 337832 260886 337884
rect 260938 337832 260944 337884
rect 261432 337832 261438 337884
rect 261490 337832 261496 337884
rect 262168 337832 262174 337884
rect 262226 337832 262232 337884
rect 262628 337832 262634 337884
rect 262686 337872 262692 337884
rect 263456 337881 263462 337884
rect 263229 337875 263287 337881
rect 263229 337872 263241 337875
rect 262686 337844 263241 337872
rect 262686 337832 262692 337844
rect 263229 337841 263241 337844
rect 263275 337841 263287 337875
rect 263229 337835 263287 337841
rect 263413 337875 263462 337881
rect 263413 337841 263425 337875
rect 263459 337841 263462 337875
rect 263413 337835 263462 337841
rect 263456 337832 263462 337835
rect 263514 337832 263520 337884
rect 258994 337668 259000 337680
rect 258874 337640 259000 337668
rect 258994 337628 259000 337640
rect 259052 337628 259058 337680
rect 259886 337612 259914 337832
rect 259178 337600 259184 337612
rect 258598 337572 259184 337600
rect 259178 337560 259184 337572
rect 259236 337560 259242 337612
rect 259886 337572 259920 337612
rect 259914 337560 259920 337572
rect 259972 337560 259978 337612
rect 256206 337504 256240 337544
rect 255924 337492 255930 337504
rect 256234 337492 256240 337504
rect 256292 337492 256298 337544
rect 260070 337532 260098 337832
rect 260898 337612 260926 337832
rect 261450 337668 261478 337832
rect 261754 337764 261760 337816
rect 261812 337804 261818 337816
rect 262076 337804 262082 337816
rect 261812 337776 262082 337804
rect 261812 337764 261818 337776
rect 262076 337764 262082 337776
rect 262134 337764 262140 337816
rect 262186 337680 262214 337832
rect 262536 337764 262542 337816
rect 262594 337804 262600 337816
rect 262953 337807 263011 337813
rect 262953 337804 262965 337807
rect 262594 337776 262965 337804
rect 262594 337764 262600 337776
rect 262953 337773 262965 337776
rect 262999 337773 263011 337807
rect 262953 337767 263011 337773
rect 261570 337668 261576 337680
rect 261450 337640 261576 337668
rect 261570 337628 261576 337640
rect 261628 337628 261634 337680
rect 262122 337628 262128 337680
rect 262180 337640 262214 337680
rect 263658 337668 263686 337900
rect 264192 337872 264198 337884
rect 264072 337844 264198 337872
rect 263824 337764 263830 337816
rect 263882 337813 263888 337816
rect 263882 337807 263931 337813
rect 263882 337773 263885 337807
rect 263919 337773 263931 337807
rect 263882 337767 263931 337773
rect 263882 337764 263888 337767
rect 263778 337668 263784 337680
rect 263658 337640 263784 337668
rect 262180 337628 262186 337640
rect 263778 337628 263784 337640
rect 263836 337628 263842 337680
rect 264072 337612 264100 337844
rect 264192 337832 264198 337844
rect 264250 337832 264256 337884
rect 264560 337832 264566 337884
rect 264618 337832 264624 337884
rect 265664 337832 265670 337884
rect 265722 337832 265728 337884
rect 265848 337832 265854 337884
rect 265906 337832 265912 337884
rect 266860 337832 266866 337884
rect 266918 337832 266924 337884
rect 266952 337832 266958 337884
rect 267010 337832 267016 337884
rect 267136 337881 267142 337884
rect 267093 337875 267142 337881
rect 267093 337841 267105 337875
rect 267139 337841 267142 337875
rect 267093 337835 267142 337841
rect 267136 337832 267142 337835
rect 267194 337832 267200 337884
rect 260834 337560 260840 337612
rect 260892 337572 260926 337612
rect 260892 337560 260898 337572
rect 264054 337560 264060 337612
rect 264112 337560 264118 337612
rect 264422 337560 264428 337612
rect 264480 337600 264486 337612
rect 264578 337600 264606 337832
rect 265682 337680 265710 337832
rect 265682 337640 265716 337680
rect 265710 337628 265716 337640
rect 265768 337628 265774 337680
rect 265866 337668 265894 337832
rect 266878 337680 266906 337832
rect 265986 337668 265992 337680
rect 265866 337640 265992 337668
rect 265986 337628 265992 337640
rect 266044 337628 266050 337680
rect 266814 337628 266820 337680
rect 266872 337640 266906 337680
rect 266970 337680 266998 337832
rect 267246 337804 267274 337900
rect 267458 337832 267464 337884
rect 267516 337872 267522 337884
rect 267645 337875 267703 337881
rect 267645 337872 267657 337875
rect 267516 337844 267657 337872
rect 267516 337832 267522 337844
rect 267645 337841 267657 337844
rect 267691 337841 267703 337875
rect 267645 337835 267703 337841
rect 267872 337832 267878 337884
rect 267930 337881 267936 337884
rect 267930 337875 267979 337881
rect 267930 337841 267933 337875
rect 267967 337841 267979 337875
rect 267930 337835 267979 337841
rect 267930 337832 267936 337835
rect 268884 337832 268890 337884
rect 268942 337832 268948 337884
rect 269252 337832 269258 337884
rect 269310 337832 269316 337884
rect 269436 337832 269442 337884
rect 269494 337832 269500 337884
rect 269758 337832 269764 337884
rect 269816 337872 269822 337884
rect 270264 337872 270270 337884
rect 269816 337844 270270 337872
rect 269816 337832 269822 337844
rect 270264 337832 270270 337844
rect 270322 337832 270328 337884
rect 270540 337832 270546 337884
rect 270598 337832 270604 337884
rect 271294 337872 271322 337900
rect 271969 337875 272027 337881
rect 271969 337872 271981 337875
rect 271294 337844 271981 337872
rect 271969 337841 271981 337844
rect 272015 337841 272027 337875
rect 271969 337835 272027 337841
rect 272104 337832 272110 337884
rect 272162 337881 272168 337884
rect 272162 337875 272211 337881
rect 272162 337841 272165 337875
rect 272199 337841 272211 337875
rect 272162 337835 272211 337841
rect 272162 337832 272168 337835
rect 272288 337832 272294 337884
rect 272346 337832 272352 337884
rect 272472 337832 272478 337884
rect 272530 337872 272536 337884
rect 272904 337872 272932 337912
rect 274085 337909 274097 337912
rect 274131 337909 274143 337943
rect 274085 337903 274143 337909
rect 276336 337900 276342 337952
rect 276394 337949 276400 337952
rect 276394 337943 276443 337949
rect 276394 337909 276397 337943
rect 276431 337909 276443 337943
rect 276394 337903 276443 337909
rect 276394 337900 276400 337903
rect 276520 337900 276526 337952
rect 276578 337940 276584 337952
rect 277213 337943 277271 337949
rect 277213 337940 277225 337943
rect 276578 337912 277225 337940
rect 276578 337900 276584 337912
rect 277213 337909 277225 337912
rect 277259 337909 277271 337943
rect 277213 337903 277271 337909
rect 278268 337900 278274 337952
rect 278326 337940 278332 337952
rect 279464 337949 279470 337952
rect 278777 337943 278835 337949
rect 278777 337940 278789 337943
rect 278326 337912 278789 337940
rect 278326 337900 278332 337912
rect 278777 337909 278789 337912
rect 278823 337909 278835 337943
rect 278777 337903 278835 337909
rect 279421 337943 279470 337949
rect 279421 337909 279433 337943
rect 279467 337909 279470 337943
rect 279421 337903 279470 337909
rect 279464 337900 279470 337903
rect 279522 337900 279528 337952
rect 279648 337900 279654 337952
rect 279706 337940 279712 337952
rect 279881 337943 279939 337949
rect 279881 337940 279893 337943
rect 279706 337912 279893 337940
rect 279706 337900 279712 337912
rect 279881 337909 279893 337912
rect 279927 337909 279939 337943
rect 279881 337903 279939 337909
rect 280660 337900 280666 337952
rect 280718 337949 280724 337952
rect 280718 337943 280767 337949
rect 280718 337909 280721 337943
rect 280755 337909 280767 337943
rect 280718 337903 280767 337909
rect 280718 337900 280724 337903
rect 281856 337900 281862 337952
rect 281914 337900 281920 337952
rect 283144 337900 283150 337952
rect 283202 337900 283208 337952
rect 283328 337900 283334 337952
rect 283386 337900 283392 337952
rect 283420 337900 283426 337952
rect 283478 337900 283484 337952
rect 284064 337900 284070 337952
rect 284122 337940 284128 337952
rect 286410 337940 286416 337952
rect 284122 337912 286416 337940
rect 284122 337900 284128 337912
rect 286410 337900 286416 337912
rect 286468 337900 286474 337952
rect 272530 337844 272932 337872
rect 272530 337832 272536 337844
rect 273024 337832 273030 337884
rect 273082 337832 273088 337884
rect 273349 337875 273407 337881
rect 273349 337841 273361 337875
rect 273395 337872 273407 337875
rect 273760 337872 273766 337884
rect 273395 337844 273766 337872
rect 273395 337841 273407 337844
rect 273349 337835 273407 337841
rect 273760 337832 273766 337844
rect 273818 337832 273824 337884
rect 274220 337832 274226 337884
rect 274278 337832 274284 337884
rect 274864 337832 274870 337884
rect 274922 337832 274928 337884
rect 275140 337832 275146 337884
rect 275198 337832 275204 337884
rect 275232 337832 275238 337884
rect 275290 337881 275296 337884
rect 275290 337875 275339 337881
rect 275290 337841 275293 337875
rect 275327 337841 275339 337875
rect 275290 337835 275339 337841
rect 275290 337832 275296 337835
rect 277348 337832 277354 337884
rect 277406 337832 277412 337884
rect 277489 337875 277547 337881
rect 277489 337841 277501 337875
rect 277535 337872 277547 337875
rect 277900 337872 277906 337884
rect 277535 337844 277906 337872
rect 277535 337841 277547 337844
rect 277489 337835 277547 337841
rect 277900 337832 277906 337844
rect 277958 337832 277964 337884
rect 278452 337872 278458 337884
rect 278148 337844 278458 337872
rect 267246 337776 267504 337804
rect 267476 337748 267504 337776
rect 267458 337696 267464 337748
rect 267516 337696 267522 337748
rect 267737 337739 267795 337745
rect 267737 337705 267749 337739
rect 267783 337736 267795 337739
rect 268286 337736 268292 337748
rect 267783 337708 268292 337736
rect 267783 337705 267795 337708
rect 267737 337699 267795 337705
rect 268286 337696 268292 337708
rect 268344 337696 268350 337748
rect 266970 337640 267004 337680
rect 266872 337628 266878 337640
rect 266998 337628 267004 337640
rect 267056 337628 267062 337680
rect 264480 337572 264606 337600
rect 264480 337560 264486 337572
rect 268286 337560 268292 337612
rect 268344 337600 268350 337612
rect 268902 337600 268930 337832
rect 269270 337668 269298 337832
rect 269454 337736 269482 337832
rect 269454 337708 269620 337736
rect 269390 337668 269396 337680
rect 269270 337640 269396 337668
rect 269390 337628 269396 337640
rect 269448 337628 269454 337680
rect 269592 337612 269620 337708
rect 268344 337572 268930 337600
rect 268344 337560 268350 337572
rect 269574 337560 269580 337612
rect 269632 337560 269638 337612
rect 260190 337532 260196 337544
rect 260070 337504 260196 337532
rect 260190 337492 260196 337504
rect 260248 337492 260254 337544
rect 270558 337532 270586 337832
rect 271644 337764 271650 337816
rect 271702 337804 271708 337816
rect 271785 337807 271843 337813
rect 271785 337804 271797 337807
rect 271702 337776 271797 337804
rect 271702 337764 271708 337776
rect 271785 337773 271797 337776
rect 271831 337773 271843 337807
rect 271785 337767 271843 337773
rect 272306 337600 272334 337832
rect 272564 337764 272570 337816
rect 272622 337813 272628 337816
rect 272622 337807 272671 337813
rect 272622 337773 272625 337807
rect 272659 337773 272671 337807
rect 272622 337767 272671 337773
rect 272622 337764 272628 337767
rect 272840 337764 272846 337816
rect 272898 337764 272904 337816
rect 272858 337680 272886 337764
rect 272858 337640 272892 337680
rect 272886 337628 272892 337640
rect 272944 337628 272950 337680
rect 272426 337600 272432 337612
rect 272306 337572 272432 337600
rect 272426 337560 272432 337572
rect 272484 337560 272490 337612
rect 273042 337600 273070 337832
rect 274036 337764 274042 337816
rect 274094 337764 274100 337816
rect 272536 337572 273070 337600
rect 272536 337544 272564 337572
rect 274054 337544 274082 337764
rect 274238 337668 274266 337832
rect 274361 337807 274419 337813
rect 274361 337773 274373 337807
rect 274407 337804 274419 337807
rect 274450 337804 274456 337816
rect 274407 337776 274456 337804
rect 274407 337773 274419 337776
rect 274361 337767 274419 337773
rect 274450 337764 274456 337776
rect 274508 337764 274514 337816
rect 274450 337668 274456 337680
rect 274238 337640 274456 337668
rect 274450 337628 274456 337640
rect 274508 337628 274514 337680
rect 274358 337600 274364 337612
rect 274319 337572 274364 337600
rect 274358 337560 274364 337572
rect 274416 337560 274422 337612
rect 274726 337560 274732 337612
rect 274784 337600 274790 337612
rect 274882 337600 274910 337832
rect 274784 337572 274910 337600
rect 274784 337560 274790 337572
rect 270770 337532 270776 337544
rect 270558 337504 270776 337532
rect 270770 337492 270776 337504
rect 270828 337492 270834 337544
rect 272518 337492 272524 337544
rect 272576 337492 272582 337544
rect 272794 337532 272800 337544
rect 272755 337504 272800 337532
rect 272794 337492 272800 337504
rect 272852 337492 272858 337544
rect 274054 337504 274088 337544
rect 274082 337492 274088 337504
rect 274140 337492 274146 337544
rect 275158 337532 275186 337832
rect 277210 337560 277216 337612
rect 277268 337600 277274 337612
rect 277366 337600 277394 337832
rect 278148 337612 278176 337844
rect 278452 337832 278458 337844
rect 278510 337832 278516 337884
rect 279740 337832 279746 337884
rect 279798 337832 279804 337884
rect 280016 337832 280022 337884
rect 280074 337832 280080 337884
rect 280568 337881 280574 337884
rect 280525 337875 280574 337881
rect 280525 337841 280537 337875
rect 280571 337841 280574 337875
rect 280525 337835 280574 337841
rect 280568 337832 280574 337835
rect 280626 337832 280632 337884
rect 280844 337872 280850 337884
rect 280816 337832 280850 337872
rect 280902 337832 280908 337884
rect 280936 337832 280942 337884
rect 280994 337832 281000 337884
rect 281120 337832 281126 337884
rect 281178 337881 281184 337884
rect 281178 337875 281227 337881
rect 281178 337841 281181 337875
rect 281215 337841 281227 337875
rect 281178 337835 281227 337841
rect 281178 337832 281184 337835
rect 281534 337832 281540 337884
rect 281592 337832 281598 337884
rect 281874 337872 281902 337900
rect 281997 337875 282055 337881
rect 281997 337872 282009 337875
rect 281874 337844 282009 337872
rect 281997 337841 282009 337844
rect 282043 337841 282055 337875
rect 281997 337835 282055 337841
rect 282132 337832 282138 337884
rect 282190 337832 282196 337884
rect 282776 337832 282782 337884
rect 282834 337832 282840 337884
rect 279602 337668 279608 337680
rect 279563 337640 279608 337668
rect 279602 337628 279608 337640
rect 279660 337628 279666 337680
rect 279758 337668 279786 337832
rect 279878 337668 279884 337680
rect 279758 337640 279884 337668
rect 279878 337628 279884 337640
rect 279936 337628 279942 337680
rect 277268 337572 277394 337600
rect 277268 337560 277274 337572
rect 278130 337560 278136 337612
rect 278188 337560 278194 337612
rect 280034 337600 280062 337832
rect 280816 337668 280844 337832
rect 280954 337748 280982 337832
rect 280890 337696 280896 337748
rect 280948 337708 280982 337748
rect 280948 337696 280954 337708
rect 281074 337668 281080 337680
rect 280816 337640 281080 337668
rect 281074 337628 281080 337640
rect 281132 337628 281138 337680
rect 279252 337572 280062 337600
rect 279252 337544 279280 337572
rect 275462 337532 275468 337544
rect 275158 337504 275468 337532
rect 275462 337492 275468 337504
rect 275520 337492 275526 337544
rect 276385 337535 276443 337541
rect 276385 337501 276397 337535
rect 276431 337532 276443 337535
rect 276750 337532 276756 337544
rect 276431 337504 276756 337532
rect 276431 337501 276443 337504
rect 276385 337495 276443 337501
rect 276750 337492 276756 337504
rect 276808 337492 276814 337544
rect 279234 337492 279240 337544
rect 279292 337492 279298 337544
rect 281552 337532 281580 337832
rect 281764 337764 281770 337816
rect 281822 337813 281828 337816
rect 281822 337807 281871 337813
rect 281822 337773 281825 337807
rect 281859 337773 281871 337807
rect 281822 337767 281871 337773
rect 281822 337764 281828 337767
rect 281626 337560 281632 337612
rect 281684 337600 281690 337612
rect 282150 337600 282178 337832
rect 282794 337680 282822 337832
rect 283162 337680 283190 337900
rect 283346 337736 283374 337900
rect 283300 337708 283374 337736
rect 283300 337680 283328 337708
rect 283438 337680 283466 337900
rect 284156 337832 284162 337884
rect 284214 337832 284220 337884
rect 284432 337832 284438 337884
rect 284490 337872 284496 337884
rect 284938 337872 284944 337884
rect 284490 337844 284944 337872
rect 284490 337832 284496 337844
rect 284938 337832 284944 337844
rect 284996 337832 285002 337884
rect 282794 337640 282828 337680
rect 282822 337628 282828 337640
rect 282880 337628 282886 337680
rect 283162 337640 283196 337680
rect 283190 337628 283196 337640
rect 283248 337628 283254 337680
rect 283282 337628 283288 337680
rect 283340 337628 283346 337680
rect 283438 337640 283472 337680
rect 283466 337628 283472 337640
rect 283524 337628 283530 337680
rect 281684 337572 282178 337600
rect 281684 337560 281690 337572
rect 281718 337532 281724 337544
rect 281552 337504 281724 337532
rect 281718 337492 281724 337504
rect 281776 337492 281782 337544
rect 255498 337464 255504 337476
rect 255459 337436 255504 337464
rect 255498 337424 255504 337436
rect 255556 337424 255562 337476
rect 273254 337464 273260 337476
rect 271892 337436 273260 337464
rect 271892 337408 271920 337436
rect 273254 337424 273260 337436
rect 273312 337424 273318 337476
rect 283742 337424 283748 337476
rect 283800 337464 283806 337476
rect 284174 337464 284202 337832
rect 283800 337436 284202 337464
rect 283800 337424 283806 337436
rect 268105 337399 268163 337405
rect 268105 337365 268117 337399
rect 268151 337396 268163 337399
rect 268194 337396 268200 337408
rect 268151 337368 268200 337396
rect 268151 337365 268163 337368
rect 268105 337359 268163 337365
rect 268194 337356 268200 337368
rect 268252 337356 268258 337408
rect 271874 337356 271880 337408
rect 271932 337356 271938 337408
rect 278774 337356 278780 337408
rect 278832 337396 278838 337408
rect 279881 337399 279939 337405
rect 279881 337396 279893 337399
rect 278832 337368 279893 337396
rect 278832 337356 278838 337368
rect 279881 337365 279893 337368
rect 279927 337365 279939 337399
rect 279881 337359 279939 337365
rect 273346 337260 273352 337272
rect 273307 337232 273352 337260
rect 273346 337220 273352 337232
rect 273404 337220 273410 337272
rect 270954 337152 270960 337204
rect 271012 337192 271018 337204
rect 277397 337195 277455 337201
rect 277397 337192 277409 337195
rect 271012 337164 277409 337192
rect 271012 337152 271018 337164
rect 277397 337161 277409 337164
rect 277443 337161 277455 337195
rect 277397 337155 277455 337161
rect 273714 337084 273720 337136
rect 273772 337124 273778 337136
rect 282825 337127 282883 337133
rect 282825 337124 282837 337127
rect 273772 337096 282837 337124
rect 273772 337084 273778 337096
rect 282825 337093 282837 337096
rect 282871 337093 282883 337127
rect 282825 337087 282883 337093
rect 236638 337016 236644 337068
rect 236696 337056 236702 337068
rect 237190 337056 237196 337068
rect 236696 337028 237196 337056
rect 236696 337016 236702 337028
rect 237190 337016 237196 337028
rect 237248 337056 237254 337068
rect 241333 337059 241391 337065
rect 241333 337056 241345 337059
rect 237248 337028 241345 337056
rect 237248 337016 237254 337028
rect 241333 337025 241345 337028
rect 241379 337025 241391 337059
rect 241333 337019 241391 337025
rect 272981 337059 273039 337065
rect 272981 337025 272993 337059
rect 273027 337056 273039 337059
rect 273349 337059 273407 337065
rect 273349 337056 273361 337059
rect 273027 337028 273361 337056
rect 273027 337025 273039 337028
rect 272981 337019 273039 337025
rect 273349 337025 273361 337028
rect 273395 337025 273407 337059
rect 273349 337019 273407 337025
rect 278866 337016 278872 337068
rect 278924 337056 278930 337068
rect 278924 337028 292574 337056
rect 278924 337016 278930 337028
rect 237834 336988 237840 337000
rect 237795 336960 237840 336988
rect 237834 336948 237840 336960
rect 237892 336948 237898 337000
rect 272889 336991 272947 336997
rect 272889 336957 272901 336991
rect 272935 336988 272947 336991
rect 273441 336991 273499 336997
rect 273441 336988 273453 336991
rect 272935 336960 273453 336988
rect 272935 336957 272947 336960
rect 272889 336951 272947 336957
rect 273441 336957 273453 336960
rect 273487 336957 273499 336991
rect 273441 336951 273499 336957
rect 282549 336991 282607 336997
rect 282549 336957 282561 336991
rect 282595 336988 282607 336991
rect 285585 336991 285643 336997
rect 285585 336988 285597 336991
rect 282595 336960 285597 336988
rect 282595 336957 282607 336960
rect 282549 336951 282607 336957
rect 285585 336957 285597 336960
rect 285631 336957 285643 336991
rect 292546 336988 292574 337028
rect 439498 336988 439504 337000
rect 292546 336960 439504 336988
rect 285585 336951 285643 336957
rect 439498 336948 439504 336960
rect 439556 336948 439562 337000
rect 271506 336880 271512 336932
rect 271564 336920 271570 336932
rect 278685 336923 278743 336929
rect 278685 336920 278697 336923
rect 271564 336892 278697 336920
rect 271564 336880 271570 336892
rect 278685 336889 278697 336892
rect 278731 336889 278743 336923
rect 278685 336883 278743 336889
rect 282454 336880 282460 336932
rect 282512 336920 282518 336932
rect 282512 336892 282914 336920
rect 282512 336880 282518 336892
rect 248969 336855 249027 336861
rect 248969 336852 248981 336855
rect 242820 336824 248981 336852
rect 235258 336744 235264 336796
rect 235316 336784 235322 336796
rect 235994 336784 236000 336796
rect 235316 336756 236000 336784
rect 235316 336744 235322 336756
rect 235994 336744 236000 336756
rect 236052 336744 236058 336796
rect 236178 336744 236184 336796
rect 236236 336784 236242 336796
rect 237098 336784 237104 336796
rect 236236 336756 237104 336784
rect 236236 336744 236242 336756
rect 237098 336744 237104 336756
rect 237156 336744 237162 336796
rect 237742 336744 237748 336796
rect 237800 336784 237806 336796
rect 242820 336784 242848 336824
rect 248969 336821 248981 336824
rect 249015 336821 249027 336855
rect 248969 336815 249027 336821
rect 261662 336812 261668 336864
rect 261720 336852 261726 336864
rect 266081 336855 266139 336861
rect 266081 336852 266093 336855
rect 261720 336824 266093 336852
rect 261720 336812 261726 336824
rect 266081 336821 266093 336824
rect 266127 336821 266139 336855
rect 266081 336815 266139 336821
rect 282886 336796 282914 336892
rect 283098 336880 283104 336932
rect 283156 336920 283162 336932
rect 568574 336920 568580 336932
rect 283156 336892 568580 336920
rect 283156 336880 283162 336892
rect 568574 336880 568580 336892
rect 568632 336880 568638 336932
rect 283190 336812 283196 336864
rect 283248 336852 283254 336864
rect 569954 336852 569960 336864
rect 283248 336824 569960 336852
rect 283248 336812 283254 336824
rect 569954 336812 569960 336824
rect 570012 336812 570018 336864
rect 237800 336756 242848 336784
rect 242897 336787 242955 336793
rect 237800 336744 237806 336756
rect 242897 336753 242909 336787
rect 242943 336784 242955 336787
rect 249153 336787 249211 336793
rect 249153 336784 249165 336787
rect 242943 336756 249165 336784
rect 242943 336753 242955 336756
rect 242897 336747 242955 336753
rect 249153 336753 249165 336756
rect 249199 336753 249211 336787
rect 272061 336787 272119 336793
rect 272061 336784 272073 336787
rect 249153 336747 249211 336753
rect 266096 336756 272073 336784
rect 86862 336676 86868 336728
rect 86920 336716 86926 336728
rect 239033 336719 239091 336725
rect 239033 336716 239045 336719
rect 86920 336688 239045 336716
rect 86920 336676 86926 336688
rect 239033 336685 239045 336688
rect 239079 336685 239091 336719
rect 239033 336679 239091 336685
rect 239309 336719 239367 336725
rect 239309 336685 239321 336719
rect 239355 336716 239367 336719
rect 242158 336716 242164 336728
rect 239355 336688 242164 336716
rect 239355 336685 239367 336688
rect 239309 336679 239367 336685
rect 242158 336676 242164 336688
rect 242216 336676 242222 336728
rect 264606 336676 264612 336728
rect 264664 336716 264670 336728
rect 266096 336716 266124 336756
rect 272061 336753 272073 336756
rect 272107 336753 272119 336787
rect 272061 336747 272119 336753
rect 272153 336787 272211 336793
rect 272153 336753 272165 336787
rect 272199 336784 272211 336787
rect 274729 336787 274787 336793
rect 272199 336756 272932 336784
rect 272199 336753 272211 336756
rect 272153 336747 272211 336753
rect 264664 336688 266124 336716
rect 264664 336676 264670 336688
rect 266170 336676 266176 336728
rect 266228 336716 266234 336728
rect 270773 336719 270831 336725
rect 270773 336716 270785 336719
rect 266228 336688 270785 336716
rect 266228 336676 266234 336688
rect 270773 336685 270785 336688
rect 270819 336685 270831 336719
rect 272904 336716 272932 336756
rect 274729 336753 274741 336787
rect 274775 336784 274787 336787
rect 274775 336756 282684 336784
rect 282886 336756 282920 336796
rect 274775 336753 274787 336756
rect 274729 336747 274787 336753
rect 274545 336719 274603 336725
rect 272904 336688 273024 336716
rect 270773 336679 270831 336685
rect 100662 336608 100668 336660
rect 100720 336648 100726 336660
rect 235261 336651 235319 336657
rect 235261 336648 235273 336651
rect 100720 336620 235273 336648
rect 100720 336608 100726 336620
rect 235261 336617 235273 336620
rect 235307 336617 235319 336651
rect 235261 336611 235319 336617
rect 235350 336608 235356 336660
rect 235408 336648 235414 336660
rect 236549 336651 236607 336657
rect 236549 336648 236561 336651
rect 235408 336620 236561 336648
rect 235408 336608 235414 336620
rect 236549 336617 236561 336620
rect 236595 336617 236607 336651
rect 236549 336611 236607 336617
rect 239217 336651 239275 336657
rect 239217 336617 239229 336651
rect 239263 336648 239275 336651
rect 245473 336651 245531 336657
rect 245473 336648 245485 336651
rect 239263 336620 245485 336648
rect 239263 336617 239275 336620
rect 239217 336611 239275 336617
rect 245473 336617 245485 336620
rect 245519 336617 245531 336651
rect 269117 336651 269175 336657
rect 269117 336648 269129 336651
rect 245473 336611 245531 336617
rect 268488 336620 269129 336648
rect 82722 336540 82728 336592
rect 82780 336580 82786 336592
rect 241882 336580 241888 336592
rect 82780 336552 241888 336580
rect 82780 336540 82786 336552
rect 241882 336540 241888 336552
rect 241940 336540 241946 336592
rect 265250 336540 265256 336592
rect 265308 336580 265314 336592
rect 268488 336580 268516 336620
rect 269117 336617 269129 336620
rect 269163 336617 269175 336651
rect 269117 336611 269175 336617
rect 269206 336608 269212 336660
rect 269264 336648 269270 336660
rect 272889 336651 272947 336657
rect 272889 336648 272901 336651
rect 269264 336620 272901 336648
rect 269264 336608 269270 336620
rect 272889 336617 272901 336620
rect 272935 336617 272947 336651
rect 272996 336648 273024 336688
rect 274545 336685 274557 336719
rect 274591 336716 274603 336719
rect 282549 336719 282607 336725
rect 282549 336716 282561 336719
rect 274591 336688 282561 336716
rect 274591 336685 274603 336688
rect 274545 336679 274603 336685
rect 282549 336685 282561 336688
rect 282595 336685 282607 336719
rect 282656 336716 282684 336756
rect 282914 336744 282920 336756
rect 282972 336744 282978 336796
rect 283282 336744 283288 336796
rect 283340 336784 283346 336796
rect 572714 336784 572720 336796
rect 283340 336756 572720 336784
rect 283340 336744 283346 336756
rect 572714 336744 572720 336756
rect 572772 336744 572778 336796
rect 347774 336716 347780 336728
rect 282656 336688 347780 336716
rect 282549 336679 282607 336685
rect 347774 336676 347780 336688
rect 347832 336676 347838 336728
rect 354674 336648 354680 336660
rect 272996 336620 354680 336648
rect 272889 336611 272947 336617
rect 354674 336608 354680 336620
rect 354732 336608 354738 336660
rect 265308 336552 268516 336580
rect 265308 336540 265314 336552
rect 268562 336540 268568 336592
rect 268620 336580 268626 336592
rect 272981 336583 273039 336589
rect 272981 336580 272993 336583
rect 268620 336552 272993 336580
rect 268620 336540 268626 336552
rect 272981 336549 272993 336552
rect 273027 336549 273039 336583
rect 272981 336543 273039 336549
rect 273073 336583 273131 336589
rect 273073 336549 273085 336583
rect 273119 336580 273131 336583
rect 361574 336580 361580 336592
rect 273119 336552 361580 336580
rect 273119 336549 273131 336552
rect 273073 336543 273131 336549
rect 361574 336540 361580 336552
rect 361632 336540 361638 336592
rect 44082 336472 44088 336524
rect 44140 336512 44146 336524
rect 235077 336515 235135 336521
rect 235077 336512 235089 336515
rect 44140 336484 235089 336512
rect 44140 336472 44146 336484
rect 235077 336481 235089 336484
rect 235123 336481 235135 336515
rect 235077 336475 235135 336481
rect 235261 336515 235319 336521
rect 235261 336481 235273 336515
rect 235307 336512 235319 336515
rect 243357 336515 243415 336521
rect 243357 336512 243369 336515
rect 235307 336484 243369 336512
rect 235307 336481 235319 336484
rect 235261 336475 235319 336481
rect 243357 336481 243369 336484
rect 243403 336481 243415 336515
rect 243357 336475 243415 336481
rect 244274 336472 244280 336524
rect 244332 336512 244338 336524
rect 249150 336512 249156 336524
rect 244332 336484 249156 336512
rect 244332 336472 244338 336484
rect 249150 336472 249156 336484
rect 249208 336472 249214 336524
rect 251174 336472 251180 336524
rect 251232 336512 251238 336524
rect 254486 336512 254492 336524
rect 251232 336484 254492 336512
rect 251232 336472 251238 336484
rect 254486 336472 254492 336484
rect 254544 336472 254550 336524
rect 260742 336472 260748 336524
rect 260800 336512 260806 336524
rect 270862 336512 270868 336524
rect 260800 336484 270868 336512
rect 260800 336472 260806 336484
rect 270862 336472 270868 336484
rect 270920 336472 270926 336524
rect 270957 336515 271015 336521
rect 270957 336481 270969 336515
rect 271003 336512 271015 336515
rect 368474 336512 368480 336524
rect 271003 336484 368480 336512
rect 271003 336481 271015 336484
rect 270957 336475 271015 336481
rect 368474 336472 368480 336484
rect 368532 336472 368538 336524
rect 75822 336404 75828 336456
rect 75880 336444 75886 336456
rect 241238 336444 241244 336456
rect 75880 336416 233924 336444
rect 75880 336404 75886 336416
rect 42702 336336 42708 336388
rect 42760 336376 42766 336388
rect 233789 336379 233847 336385
rect 233789 336376 233801 336379
rect 42760 336348 233801 336376
rect 42760 336336 42766 336348
rect 233789 336345 233801 336348
rect 233835 336345 233847 336379
rect 233896 336376 233924 336416
rect 238680 336416 241244 336444
rect 238680 336376 238708 336416
rect 241238 336404 241244 336416
rect 241296 336404 241302 336456
rect 241333 336447 241391 336453
rect 241333 336413 241345 336447
rect 241379 336444 241391 336447
rect 242897 336447 242955 336453
rect 242897 336444 242909 336447
rect 241379 336416 242909 336444
rect 241379 336413 241391 336416
rect 241333 336407 241391 336413
rect 242897 336413 242909 336416
rect 242943 336413 242955 336447
rect 242897 336407 242955 336413
rect 242986 336404 242992 336456
rect 243044 336444 243050 336456
rect 253017 336447 253075 336453
rect 253017 336444 253029 336447
rect 243044 336416 253029 336444
rect 243044 336404 243050 336416
rect 253017 336413 253029 336416
rect 253063 336413 253075 336447
rect 253017 336407 253075 336413
rect 260834 336404 260840 336456
rect 260892 336444 260898 336456
rect 263505 336447 263563 336453
rect 263505 336444 263517 336447
rect 260892 336416 263517 336444
rect 260892 336404 260898 336416
rect 263505 336413 263517 336416
rect 263551 336413 263563 336447
rect 263505 336407 263563 336413
rect 266446 336404 266452 336456
rect 266504 336444 266510 336456
rect 372614 336444 372620 336456
rect 266504 336416 372620 336444
rect 266504 336404 266510 336416
rect 372614 336404 372620 336416
rect 372672 336404 372678 336456
rect 233896 336348 238708 336376
rect 239309 336379 239367 336385
rect 233789 336339 233847 336345
rect 239309 336345 239321 336379
rect 239355 336376 239367 336379
rect 241149 336379 241207 336385
rect 241149 336376 241161 336379
rect 239355 336348 241161 336376
rect 239355 336345 239367 336348
rect 239309 336339 239367 336345
rect 241149 336345 241161 336348
rect 241195 336345 241207 336379
rect 241149 336339 241207 336345
rect 241425 336379 241483 336385
rect 241425 336345 241437 336379
rect 241471 336376 241483 336379
rect 245289 336379 245347 336385
rect 245289 336376 245301 336379
rect 241471 336348 245301 336376
rect 241471 336345 241483 336348
rect 241425 336339 241483 336345
rect 245289 336345 245301 336348
rect 245335 336345 245347 336379
rect 245289 336339 245347 336345
rect 245562 336336 245568 336388
rect 245620 336376 245626 336388
rect 253934 336376 253940 336388
rect 245620 336348 253940 336376
rect 245620 336336 245626 336348
rect 253934 336336 253940 336348
rect 253992 336336 253998 336388
rect 260469 336379 260527 336385
rect 260469 336345 260481 336379
rect 260515 336376 260527 336379
rect 260515 336348 266492 336376
rect 260515 336345 260527 336348
rect 260469 336339 260527 336345
rect 266464 336320 266492 336348
rect 266906 336336 266912 336388
rect 266964 336376 266970 336388
rect 375374 336376 375380 336388
rect 266964 336348 375380 336376
rect 266964 336336 266970 336348
rect 375374 336336 375380 336348
rect 375432 336336 375438 336388
rect 28902 336268 28908 336320
rect 28960 336308 28966 336320
rect 237282 336308 237288 336320
rect 28960 336280 237288 336308
rect 28960 336268 28966 336280
rect 237282 336268 237288 336280
rect 237340 336268 237346 336320
rect 241698 336268 241704 336320
rect 241756 336308 241762 336320
rect 241882 336308 241888 336320
rect 241756 336280 241888 336308
rect 241756 336268 241762 336280
rect 241882 336268 241888 336280
rect 241940 336268 241946 336320
rect 241977 336311 242035 336317
rect 241977 336277 241989 336311
rect 242023 336308 242035 336311
rect 244001 336311 244059 336317
rect 244001 336308 244013 336311
rect 242023 336280 244013 336308
rect 242023 336277 242035 336280
rect 241977 336271 242035 336277
rect 244001 336277 244013 336280
rect 244047 336277 244059 336311
rect 244001 336271 244059 336277
rect 244093 336311 244151 336317
rect 244093 336277 244105 336311
rect 244139 336308 244151 336311
rect 248874 336308 248880 336320
rect 244139 336280 248880 336308
rect 244139 336277 244151 336280
rect 244093 336271 244151 336277
rect 248874 336268 248880 336280
rect 248932 336268 248938 336320
rect 266446 336268 266452 336320
rect 266504 336268 266510 336320
rect 266538 336268 266544 336320
rect 266596 336308 266602 336320
rect 266722 336308 266728 336320
rect 266596 336280 266728 336308
rect 266596 336268 266602 336280
rect 266722 336268 266728 336280
rect 266780 336268 266786 336320
rect 267369 336311 267427 336317
rect 267369 336277 267381 336311
rect 267415 336308 267427 336311
rect 382274 336308 382280 336320
rect 267415 336280 382280 336308
rect 267415 336277 267427 336280
rect 267369 336271 267427 336277
rect 382274 336268 382280 336280
rect 382332 336268 382338 336320
rect 20622 336200 20628 336252
rect 20680 336240 20686 336252
rect 236546 336240 236552 336252
rect 20680 336212 236552 336240
rect 20680 336200 20686 336212
rect 236546 336200 236552 336212
rect 236604 336200 236610 336252
rect 237006 336200 237012 336252
rect 237064 336240 237070 336252
rect 242621 336243 242679 336249
rect 242621 336240 242633 336243
rect 237064 336212 242633 336240
rect 237064 336200 237070 336212
rect 242621 336209 242633 336212
rect 242667 336209 242679 336243
rect 242621 336203 242679 336209
rect 243354 336200 243360 336252
rect 243412 336240 243418 336252
rect 258810 336240 258816 336252
rect 243412 336212 258816 336240
rect 243412 336200 243418 336212
rect 258810 336200 258816 336212
rect 258868 336200 258874 336252
rect 266633 336243 266691 336249
rect 266633 336209 266645 336243
rect 266679 336240 266691 336243
rect 272153 336243 272211 336249
rect 272153 336240 272165 336243
rect 266679 336212 272165 336240
rect 266679 336209 266691 336212
rect 266633 336203 266691 336209
rect 272153 336209 272165 336212
rect 272199 336209 272211 336243
rect 272153 336203 272211 336209
rect 273441 336243 273499 336249
rect 273441 336209 273453 336243
rect 273487 336240 273499 336243
rect 275925 336243 275983 336249
rect 275925 336240 275937 336243
rect 273487 336212 275937 336240
rect 273487 336209 273499 336212
rect 273441 336203 273499 336209
rect 275925 336209 275937 336212
rect 275971 336209 275983 336243
rect 275925 336203 275983 336209
rect 276014 336200 276020 336252
rect 276072 336240 276078 336252
rect 276934 336240 276940 336252
rect 276072 336212 276940 336240
rect 276072 336200 276078 336212
rect 276934 336200 276940 336212
rect 276992 336200 276998 336252
rect 277581 336243 277639 336249
rect 277581 336240 277593 336243
rect 277044 336212 277593 336240
rect 233789 336175 233847 336181
rect 233789 336141 233801 336175
rect 233835 336172 233847 336175
rect 238478 336172 238484 336184
rect 233835 336144 238484 336172
rect 233835 336141 233847 336144
rect 233789 336135 233847 336141
rect 238478 336132 238484 336144
rect 238536 336132 238542 336184
rect 245013 336175 245071 336181
rect 245013 336172 245025 336175
rect 238588 336144 245025 336172
rect 7558 336064 7564 336116
rect 7616 336104 7622 336116
rect 235534 336104 235540 336116
rect 7616 336076 235540 336104
rect 7616 336064 7622 336076
rect 235534 336064 235540 336076
rect 235592 336064 235598 336116
rect 235629 336107 235687 336113
rect 235629 336073 235641 336107
rect 235675 336104 235687 336107
rect 238588 336104 238616 336144
rect 245013 336141 245025 336144
rect 245059 336141 245071 336175
rect 245013 336135 245071 336141
rect 250530 336132 250536 336184
rect 250588 336172 250594 336184
rect 254946 336172 254952 336184
rect 250588 336144 254952 336172
rect 250588 336132 250594 336144
rect 254946 336132 254952 336144
rect 255004 336132 255010 336184
rect 257709 336175 257767 336181
rect 257709 336141 257721 336175
rect 257755 336172 257767 336175
rect 263870 336172 263876 336184
rect 257755 336144 263876 336172
rect 257755 336141 257767 336144
rect 257709 336135 257767 336141
rect 263870 336132 263876 336144
rect 263928 336132 263934 336184
rect 269301 336175 269359 336181
rect 269301 336141 269313 336175
rect 269347 336172 269359 336175
rect 270865 336175 270923 336181
rect 270865 336172 270877 336175
rect 269347 336144 270877 336172
rect 269347 336141 269359 336144
rect 269301 336135 269359 336141
rect 270865 336141 270877 336144
rect 270911 336141 270923 336175
rect 270865 336135 270923 336141
rect 273349 336175 273407 336181
rect 273349 336141 273361 336175
rect 273395 336172 273407 336175
rect 277044 336172 277072 336212
rect 277581 336209 277593 336212
rect 277627 336209 277639 336243
rect 277581 336203 277639 336209
rect 277670 336200 277676 336252
rect 277728 336240 277734 336252
rect 278682 336240 278688 336252
rect 277728 336212 278688 336240
rect 277728 336200 277734 336212
rect 278682 336200 278688 336212
rect 278740 336200 278746 336252
rect 397454 336240 397460 336252
rect 278792 336212 397460 336240
rect 273395 336144 277072 336172
rect 278409 336175 278467 336181
rect 273395 336141 273407 336144
rect 273349 336135 273407 336141
rect 278409 336141 278421 336175
rect 278455 336172 278467 336175
rect 278792 336172 278820 336212
rect 397454 336200 397460 336212
rect 397512 336200 397518 336252
rect 404354 336172 404360 336184
rect 278455 336144 278820 336172
rect 278884 336144 404360 336172
rect 278455 336141 278467 336144
rect 278409 336135 278467 336141
rect 235675 336076 238616 336104
rect 238665 336107 238723 336113
rect 235675 336073 235687 336076
rect 235629 336067 235687 336073
rect 238665 336073 238677 336107
rect 238711 336104 238723 336107
rect 241609 336107 241667 336113
rect 241609 336104 241621 336107
rect 238711 336076 241621 336104
rect 238711 336073 238723 336076
rect 238665 336067 238723 336073
rect 241609 336073 241621 336076
rect 241655 336073 241667 336107
rect 241609 336067 241667 336073
rect 241698 336064 241704 336116
rect 241756 336104 241762 336116
rect 252741 336107 252799 336113
rect 252741 336104 252753 336107
rect 241756 336076 252753 336104
rect 241756 336064 241762 336076
rect 252741 336073 252753 336076
rect 252787 336073 252799 336107
rect 252741 336067 252799 336073
rect 257246 336064 257252 336116
rect 257304 336104 257310 336116
rect 262217 336107 262275 336113
rect 262217 336104 262229 336107
rect 257304 336076 262229 336104
rect 257304 336064 257310 336076
rect 262217 336073 262229 336076
rect 262263 336073 262275 336107
rect 262217 336067 262275 336073
rect 263413 336107 263471 336113
rect 263413 336073 263425 336107
rect 263459 336104 263471 336107
rect 272242 336104 272248 336116
rect 263459 336076 272248 336104
rect 263459 336073 263471 336076
rect 263413 336067 263471 336073
rect 272242 336064 272248 336076
rect 272300 336064 272306 336116
rect 274910 336064 274916 336116
rect 274968 336104 274974 336116
rect 275738 336104 275744 336116
rect 274968 336076 275744 336104
rect 274968 336064 274974 336076
rect 275738 336064 275744 336076
rect 275796 336064 275802 336116
rect 275830 336064 275836 336116
rect 275888 336104 275894 336116
rect 275888 336076 275933 336104
rect 275888 336064 275894 336076
rect 276106 336064 276112 336116
rect 276164 336104 276170 336116
rect 276937 336107 276995 336113
rect 276937 336104 276949 336107
rect 276164 336076 276949 336104
rect 276164 336064 276170 336076
rect 276937 336073 276949 336076
rect 276983 336073 276995 336107
rect 276937 336067 276995 336073
rect 277578 336064 277584 336116
rect 277636 336104 277642 336116
rect 278498 336104 278504 336116
rect 277636 336076 278504 336104
rect 277636 336064 277642 336076
rect 278498 336064 278504 336076
rect 278556 336064 278562 336116
rect 278593 336107 278651 336113
rect 278593 336073 278605 336107
rect 278639 336104 278651 336107
rect 278884 336104 278912 336144
rect 404354 336132 404360 336144
rect 404412 336132 404418 336184
rect 278639 336076 278912 336104
rect 278639 336073 278651 336076
rect 278593 336067 278651 336073
rect 280338 336064 280344 336116
rect 280396 336104 280402 336116
rect 281258 336104 281264 336116
rect 280396 336076 281264 336104
rect 280396 336064 280402 336076
rect 281258 336064 281264 336076
rect 281316 336064 281322 336116
rect 282457 336107 282515 336113
rect 282457 336073 282469 336107
rect 282503 336104 282515 336107
rect 411254 336104 411260 336116
rect 282503 336076 411260 336104
rect 282503 336073 282515 336076
rect 282457 336067 282515 336073
rect 411254 336064 411260 336076
rect 411312 336064 411318 336116
rect 5442 335996 5448 336048
rect 5500 336036 5506 336048
rect 235442 336036 235448 336048
rect 5500 336008 235448 336036
rect 5500 335996 5506 336008
rect 235442 335996 235448 336008
rect 235500 335996 235506 336048
rect 236641 336039 236699 336045
rect 236641 336005 236653 336039
rect 236687 336036 236699 336039
rect 238481 336039 238539 336045
rect 238481 336036 238493 336039
rect 236687 336008 238493 336036
rect 236687 336005 236699 336008
rect 236641 335999 236699 336005
rect 238481 336005 238493 336008
rect 238527 336005 238539 336039
rect 238481 335999 238539 336005
rect 238570 335996 238576 336048
rect 238628 336036 238634 336048
rect 242345 336039 242403 336045
rect 242345 336036 242357 336039
rect 238628 336008 242357 336036
rect 238628 335996 238634 336008
rect 242345 336005 242357 336008
rect 242391 336005 242403 336039
rect 242345 335999 242403 336005
rect 242437 336039 242495 336045
rect 242437 336005 242449 336039
rect 242483 336036 242495 336039
rect 252554 336036 252560 336048
rect 242483 336008 252560 336036
rect 242483 336005 242495 336008
rect 242437 335999 242495 336005
rect 252554 335996 252560 336008
rect 252612 335996 252618 336048
rect 261386 335996 261392 336048
rect 261444 336036 261450 336048
rect 263594 336036 263600 336048
rect 261444 336008 263600 336036
rect 261444 335996 261450 336008
rect 263594 335996 263600 336008
rect 263652 335996 263658 336048
rect 265986 335996 265992 336048
rect 266044 336036 266050 336048
rect 270221 336039 270279 336045
rect 270221 336036 270233 336039
rect 266044 336008 270233 336036
rect 266044 335996 266050 336008
rect 270221 336005 270233 336008
rect 270267 336005 270279 336039
rect 270221 335999 270279 336005
rect 270310 335996 270316 336048
rect 270368 336036 270374 336048
rect 418154 336036 418160 336048
rect 270368 336008 418160 336036
rect 270368 335996 270374 336008
rect 418154 335996 418160 336008
rect 418212 335996 418218 336048
rect 93762 335928 93768 335980
rect 93820 335968 93826 335980
rect 241974 335968 241980 335980
rect 93820 335940 241980 335968
rect 93820 335928 93826 335940
rect 241974 335928 241980 335940
rect 242032 335928 242038 335980
rect 242805 335971 242863 335977
rect 242805 335937 242817 335971
rect 242851 335968 242863 335971
rect 243814 335968 243820 335980
rect 242851 335940 243820 335968
rect 242851 335937 242863 335940
rect 242805 335931 242863 335937
rect 243814 335928 243820 335940
rect 243872 335928 243878 335980
rect 244366 335928 244372 335980
rect 244424 335968 244430 335980
rect 253474 335968 253480 335980
rect 244424 335940 253480 335968
rect 244424 335928 244430 335940
rect 253474 335928 253480 335940
rect 253532 335928 253538 335980
rect 257617 335971 257675 335977
rect 257617 335937 257629 335971
rect 257663 335968 257675 335971
rect 262861 335971 262919 335977
rect 262861 335968 262873 335971
rect 257663 335940 262873 335968
rect 257663 335937 257675 335940
rect 257617 335931 257675 335937
rect 262861 335937 262873 335940
rect 262907 335937 262919 335971
rect 262861 335931 262919 335937
rect 264146 335928 264152 335980
rect 264204 335968 264210 335980
rect 264698 335968 264704 335980
rect 264204 335940 264704 335968
rect 264204 335928 264210 335940
rect 264698 335928 264704 335940
rect 264756 335928 264762 335980
rect 265618 335928 265624 335980
rect 265676 335968 265682 335980
rect 272981 335971 273039 335977
rect 272981 335968 272993 335971
rect 265676 335940 272993 335968
rect 265676 335928 265682 335940
rect 272981 335937 272993 335940
rect 273027 335937 273039 335971
rect 272981 335931 273039 335937
rect 273165 335971 273223 335977
rect 273165 335937 273177 335971
rect 273211 335968 273223 335971
rect 274729 335971 274787 335977
rect 274729 335968 274741 335971
rect 273211 335940 274741 335968
rect 273211 335937 273223 335940
rect 273165 335931 273223 335937
rect 274729 335937 274741 335940
rect 274775 335937 274787 335971
rect 274729 335931 274787 335937
rect 274818 335928 274824 335980
rect 274876 335968 274882 335980
rect 275830 335968 275836 335980
rect 274876 335940 275836 335968
rect 274876 335928 274882 335940
rect 275830 335928 275836 335940
rect 275888 335928 275894 335980
rect 275925 335971 275983 335977
rect 275925 335937 275937 335971
rect 275971 335968 275983 335971
rect 277765 335971 277823 335977
rect 277765 335968 277777 335971
rect 275971 335940 277777 335968
rect 275971 335937 275983 335940
rect 275925 335931 275983 335937
rect 277765 335937 277777 335940
rect 277811 335937 277823 335971
rect 277765 335931 277823 335937
rect 278685 335971 278743 335977
rect 278685 335937 278697 335971
rect 278731 335968 278743 335971
rect 300118 335968 300124 335980
rect 278731 335940 300124 335968
rect 278731 335937 278743 335940
rect 278685 335931 278743 335937
rect 300118 335928 300124 335940
rect 300176 335928 300182 335980
rect 107562 335860 107568 335912
rect 107620 335900 107626 335912
rect 243906 335900 243912 335912
rect 107620 335872 243912 335900
rect 107620 335860 107626 335872
rect 243906 335860 243912 335872
rect 243964 335860 243970 335912
rect 244001 335903 244059 335909
rect 244001 335869 244013 335903
rect 244047 335900 244059 335903
rect 257246 335900 257252 335912
rect 244047 335872 257252 335900
rect 244047 335869 244059 335872
rect 244001 335863 244059 335869
rect 257246 335860 257252 335872
rect 257304 335860 257310 335912
rect 260466 335860 260472 335912
rect 260524 335900 260530 335912
rect 262398 335900 262404 335912
rect 260524 335872 262404 335900
rect 260524 335860 260530 335872
rect 262398 335860 262404 335872
rect 262456 335860 262462 335912
rect 262953 335903 263011 335909
rect 262953 335869 262965 335903
rect 262999 335900 263011 335903
rect 270494 335900 270500 335912
rect 262999 335872 270500 335900
rect 262999 335869 263011 335872
rect 262953 335863 263011 335869
rect 270494 335860 270500 335872
rect 270552 335860 270558 335912
rect 275094 335860 275100 335912
rect 275152 335900 275158 335912
rect 275738 335900 275744 335912
rect 275152 335872 275744 335900
rect 275152 335860 275158 335872
rect 275738 335860 275744 335872
rect 275796 335860 275802 335912
rect 276106 335860 276112 335912
rect 276164 335900 276170 335912
rect 276842 335900 276848 335912
rect 276164 335872 276848 335900
rect 276164 335860 276170 335872
rect 276842 335860 276848 335872
rect 276900 335860 276906 335912
rect 277210 335860 277216 335912
rect 277268 335900 277274 335912
rect 277305 335903 277363 335909
rect 277305 335900 277317 335903
rect 277268 335872 277317 335900
rect 277268 335860 277274 335872
rect 277305 335869 277317 335872
rect 277351 335869 277363 335903
rect 277305 335863 277363 335869
rect 277489 335903 277547 335909
rect 277489 335869 277501 335903
rect 277535 335900 277547 335903
rect 277578 335900 277584 335912
rect 277535 335872 277584 335900
rect 277535 335869 277547 335872
rect 277489 335863 277547 335869
rect 277578 335860 277584 335872
rect 277636 335860 277642 335912
rect 280246 335860 280252 335912
rect 280304 335900 280310 335912
rect 280433 335903 280491 335909
rect 280433 335900 280445 335903
rect 280304 335872 280445 335900
rect 280304 335860 280310 335872
rect 280433 335869 280445 335872
rect 280479 335869 280491 335903
rect 280433 335863 280491 335869
rect 283009 335903 283067 335909
rect 283009 335869 283021 335903
rect 283055 335900 283067 335903
rect 287333 335903 287391 335909
rect 287333 335900 287345 335903
rect 283055 335872 287345 335900
rect 283055 335869 283067 335872
rect 283009 335863 283067 335869
rect 287333 335869 287345 335872
rect 287379 335869 287391 335903
rect 287333 335863 287391 335869
rect 287606 335860 287612 335912
rect 287664 335900 287670 335912
rect 288250 335900 288256 335912
rect 287664 335872 288256 335900
rect 287664 335860 287670 335872
rect 288250 335860 288256 335872
rect 288308 335860 288314 335912
rect 296070 335900 296076 335912
rect 292546 335872 296076 335900
rect 114462 335792 114468 335844
rect 114520 335832 114526 335844
rect 114520 335804 239444 335832
rect 114520 335792 114526 335804
rect 125502 335724 125508 335776
rect 125560 335764 125566 335776
rect 239217 335767 239275 335773
rect 239217 335764 239229 335767
rect 125560 335736 239229 335764
rect 125560 335724 125566 335736
rect 239217 335733 239229 335736
rect 239263 335733 239275 335767
rect 239217 335727 239275 335733
rect 124122 335656 124128 335708
rect 124180 335696 124186 335708
rect 239309 335699 239367 335705
rect 239309 335696 239321 335699
rect 124180 335668 239321 335696
rect 124180 335656 124186 335668
rect 239309 335665 239321 335668
rect 239355 335665 239367 335699
rect 239416 335696 239444 335804
rect 240778 335792 240784 335844
rect 240836 335832 240842 335844
rect 241514 335832 241520 335844
rect 240836 335804 241520 335832
rect 240836 335792 240842 335804
rect 241514 335792 241520 335804
rect 241572 335792 241578 335844
rect 242342 335792 242348 335844
rect 242400 335832 242406 335844
rect 244182 335832 244188 335844
rect 242400 335804 244188 335832
rect 242400 335792 242406 335804
rect 244182 335792 244188 335804
rect 244240 335792 244246 335844
rect 259730 335792 259736 335844
rect 259788 335832 259794 335844
rect 262769 335835 262827 335841
rect 262769 335832 262781 335835
rect 259788 335804 262781 335832
rect 259788 335792 259794 335804
rect 262769 335801 262781 335804
rect 262815 335801 262827 335835
rect 262769 335795 262827 335801
rect 262861 335835 262919 335841
rect 262861 335801 262873 335835
rect 262907 335832 262919 335835
rect 266538 335832 266544 335844
rect 262907 335804 266544 335832
rect 262907 335801 262919 335804
rect 262861 335795 262919 335801
rect 266538 335792 266544 335804
rect 266596 335792 266602 335844
rect 268010 335792 268016 335844
rect 268068 335832 268074 335844
rect 270681 335835 270739 335841
rect 270681 335832 270693 335835
rect 268068 335804 270693 335832
rect 268068 335792 268074 335804
rect 270681 335801 270693 335804
rect 270727 335801 270739 335835
rect 283101 335835 283159 335841
rect 270681 335795 270739 335801
rect 273226 335804 282914 335832
rect 239493 335767 239551 335773
rect 239493 335733 239505 335767
rect 239539 335764 239551 335767
rect 243265 335767 243323 335773
rect 243265 335764 243277 335767
rect 239539 335736 243277 335764
rect 239539 335733 239551 335736
rect 239493 335727 239551 335733
rect 243265 335733 243277 335736
rect 243311 335733 243323 335767
rect 243265 335727 243323 335733
rect 249150 335724 249156 335776
rect 249208 335764 249214 335776
rect 254213 335767 254271 335773
rect 254213 335764 254225 335767
rect 249208 335736 254225 335764
rect 249208 335724 249214 335736
rect 254213 335733 254225 335736
rect 254259 335733 254271 335767
rect 254213 335727 254271 335733
rect 258074 335724 258080 335776
rect 258132 335764 258138 335776
rect 263226 335764 263232 335776
rect 258132 335736 261708 335764
rect 263187 335736 263232 335764
rect 258132 335724 258138 335736
rect 244642 335696 244648 335708
rect 239416 335668 244648 335696
rect 239309 335659 239367 335665
rect 244642 335656 244648 335668
rect 244700 335656 244706 335708
rect 245102 335656 245108 335708
rect 245160 335696 245166 335708
rect 251269 335699 251327 335705
rect 251269 335696 251281 335699
rect 245160 335668 251281 335696
rect 245160 335656 245166 335668
rect 251269 335665 251281 335668
rect 251315 335665 251327 335699
rect 251269 335659 251327 335665
rect 258166 335656 258172 335708
rect 258224 335696 258230 335708
rect 258350 335696 258356 335708
rect 258224 335668 258356 335696
rect 258224 335656 258230 335668
rect 258350 335656 258356 335668
rect 258408 335656 258414 335708
rect 259454 335656 259460 335708
rect 259512 335696 259518 335708
rect 259730 335696 259736 335708
rect 259512 335668 259736 335696
rect 259512 335656 259518 335668
rect 259730 335656 259736 335668
rect 259788 335656 259794 335708
rect 260006 335656 260012 335708
rect 260064 335696 260070 335708
rect 260374 335696 260380 335708
rect 260064 335668 260380 335696
rect 260064 335656 260070 335668
rect 260374 335656 260380 335668
rect 260432 335656 260438 335708
rect 261680 335696 261708 335736
rect 263226 335724 263232 335736
rect 263284 335724 263290 335776
rect 266630 335724 266636 335776
rect 266688 335764 266694 335776
rect 267090 335764 267096 335776
rect 266688 335736 267096 335764
rect 266688 335724 266694 335736
rect 267090 335724 267096 335736
rect 267148 335724 267154 335776
rect 267461 335767 267519 335773
rect 267461 335733 267473 335767
rect 267507 335764 267519 335767
rect 269114 335764 269120 335776
rect 267507 335736 269120 335764
rect 267507 335733 267519 335736
rect 267461 335727 267519 335733
rect 269114 335724 269120 335736
rect 269172 335724 269178 335776
rect 269853 335767 269911 335773
rect 269853 335733 269865 335767
rect 269899 335764 269911 335767
rect 273073 335767 273131 335773
rect 273073 335764 273085 335767
rect 269899 335736 273085 335764
rect 269899 335733 269911 335736
rect 269853 335727 269911 335733
rect 273073 335733 273085 335736
rect 273119 335733 273131 335767
rect 273073 335727 273131 335733
rect 262674 335696 262680 335708
rect 261680 335668 262680 335696
rect 262674 335656 262680 335668
rect 262732 335656 262738 335708
rect 262769 335699 262827 335705
rect 262769 335665 262781 335699
rect 262815 335696 262827 335699
rect 266081 335699 266139 335705
rect 262815 335668 263594 335696
rect 262815 335665 262827 335668
rect 262769 335659 262827 335665
rect 234246 335588 234252 335640
rect 234304 335628 234310 335640
rect 244550 335628 244556 335640
rect 234304 335600 244556 335628
rect 234304 335588 234310 335600
rect 244550 335588 244556 335600
rect 244608 335588 244614 335640
rect 245378 335588 245384 335640
rect 245436 335628 245442 335640
rect 247770 335628 247776 335640
rect 245436 335600 247776 335628
rect 245436 335588 245442 335600
rect 247770 335588 247776 335600
rect 247828 335588 247834 335640
rect 254946 335588 254952 335640
rect 255004 335628 255010 335640
rect 255130 335628 255136 335640
rect 255004 335600 255136 335628
rect 255004 335588 255010 335600
rect 255130 335588 255136 335600
rect 255188 335588 255194 335640
rect 257062 335588 257068 335640
rect 257120 335628 257126 335640
rect 260098 335628 260104 335640
rect 257120 335600 260104 335628
rect 257120 335588 257126 335600
rect 260098 335588 260104 335600
rect 260156 335588 260162 335640
rect 263566 335628 263594 335668
rect 266081 335665 266093 335699
rect 266127 335696 266139 335699
rect 266127 335668 270540 335696
rect 266127 335665 266139 335668
rect 266081 335659 266139 335665
rect 264146 335628 264152 335640
rect 263566 335600 264152 335628
rect 264146 335588 264152 335600
rect 264204 335588 264210 335640
rect 264698 335588 264704 335640
rect 264756 335628 264762 335640
rect 267461 335631 267519 335637
rect 267461 335628 267473 335631
rect 264756 335600 267473 335628
rect 264756 335588 264762 335600
rect 267461 335597 267473 335600
rect 267507 335597 267519 335631
rect 267461 335591 267519 335597
rect 267642 335588 267648 335640
rect 267700 335628 267706 335640
rect 269945 335631 270003 335637
rect 269945 335628 269957 335631
rect 267700 335600 269957 335628
rect 267700 335588 267706 335600
rect 269945 335597 269957 335600
rect 269991 335597 270003 335631
rect 269945 335591 270003 335597
rect 234062 335520 234068 335572
rect 234120 335560 234126 335572
rect 234985 335563 235043 335569
rect 234985 335560 234997 335563
rect 234120 335532 234997 335560
rect 234120 335520 234126 335532
rect 234985 335529 234997 335532
rect 235031 335529 235043 335563
rect 242805 335563 242863 335569
rect 242805 335560 242817 335563
rect 234985 335523 235043 335529
rect 235092 335532 242817 335560
rect 234154 335452 234160 335504
rect 234212 335492 234218 335504
rect 235092 335492 235120 335532
rect 242805 335529 242817 335532
rect 242851 335529 242863 335563
rect 242805 335523 242863 335529
rect 253906 335532 259316 335560
rect 234212 335464 235120 335492
rect 235169 335495 235227 335501
rect 234212 335452 234218 335464
rect 235169 335461 235181 335495
rect 235215 335492 235227 335495
rect 239493 335495 239551 335501
rect 239493 335492 239505 335495
rect 235215 335464 239505 335492
rect 235215 335461 235227 335464
rect 235169 335455 235227 335461
rect 239493 335461 239505 335464
rect 239539 335461 239551 335495
rect 239493 335455 239551 335461
rect 248969 335495 249027 335501
rect 248969 335461 248981 335495
rect 249015 335492 249027 335495
rect 253906 335492 253934 335532
rect 249015 335464 253934 335492
rect 249015 335461 249027 335464
rect 248969 335455 249027 335461
rect 256786 335452 256792 335504
rect 256844 335492 256850 335504
rect 258074 335492 258080 335504
rect 256844 335464 258080 335492
rect 256844 335452 256850 335464
rect 258074 335452 258080 335464
rect 258132 335452 258138 335504
rect 258258 335452 258264 335504
rect 258316 335492 258322 335504
rect 259288 335492 259316 335532
rect 259454 335520 259460 335572
rect 259512 335560 259518 335572
rect 260282 335560 260288 335572
rect 259512 335532 260288 335560
rect 259512 335520 259518 335532
rect 260282 335520 260288 335532
rect 260340 335520 260346 335572
rect 262858 335560 262864 335572
rect 262819 335532 262864 335560
rect 262858 335520 262864 335532
rect 262916 335520 262922 335572
rect 263134 335520 263140 335572
rect 263192 335560 263198 335572
rect 263192 335532 263410 335560
rect 263192 335520 263198 335532
rect 259546 335492 259552 335504
rect 258316 335464 259224 335492
rect 259288 335464 259552 335492
rect 258316 335452 258322 335464
rect 10962 335384 10968 335436
rect 11020 335424 11026 335436
rect 235718 335424 235724 335436
rect 11020 335396 235724 335424
rect 11020 335384 11026 335396
rect 235718 335384 235724 335396
rect 235776 335384 235782 335436
rect 235994 335384 236000 335436
rect 236052 335424 236058 335436
rect 236362 335424 236368 335436
rect 236052 335396 236368 335424
rect 236052 335384 236058 335396
rect 236362 335384 236368 335396
rect 236420 335424 236426 335436
rect 238757 335427 238815 335433
rect 236420 335396 237328 335424
rect 236420 335384 236426 335396
rect 234338 335316 234344 335368
rect 234396 335356 234402 335368
rect 235169 335359 235227 335365
rect 235169 335356 235181 335359
rect 234396 335328 235181 335356
rect 234396 335316 234402 335328
rect 235169 335325 235181 335328
rect 235215 335325 235227 335359
rect 235169 335319 235227 335325
rect 236178 335316 236184 335368
rect 236236 335356 236242 335368
rect 237190 335356 237196 335368
rect 236236 335328 237196 335356
rect 236236 335316 236242 335328
rect 237190 335316 237196 335328
rect 237248 335316 237254 335368
rect 237300 335356 237328 335396
rect 238757 335393 238769 335427
rect 238803 335424 238815 335427
rect 242986 335424 242992 335436
rect 238803 335396 242992 335424
rect 238803 335393 238815 335396
rect 238757 335387 238815 335393
rect 242986 335384 242992 335396
rect 243044 335384 243050 335436
rect 243170 335384 243176 335436
rect 243228 335424 243234 335436
rect 243449 335427 243507 335433
rect 243449 335424 243461 335427
rect 243228 335396 243461 335424
rect 243228 335384 243234 335396
rect 243449 335393 243461 335396
rect 243495 335393 243507 335427
rect 243449 335387 243507 335393
rect 249153 335427 249211 335433
rect 249153 335393 249165 335427
rect 249199 335424 249211 335427
rect 255130 335424 255136 335436
rect 249199 335396 255136 335424
rect 249199 335393 249211 335396
rect 249153 335387 249211 335393
rect 255130 335384 255136 335396
rect 255188 335384 255194 335436
rect 258442 335384 258448 335436
rect 258500 335424 258506 335436
rect 259086 335424 259092 335436
rect 258500 335396 259092 335424
rect 258500 335384 258506 335396
rect 259086 335384 259092 335396
rect 259144 335384 259150 335436
rect 242069 335359 242127 335365
rect 242069 335356 242081 335359
rect 237300 335328 242081 335356
rect 242069 335325 242081 335328
rect 242115 335325 242127 335359
rect 242069 335319 242127 335325
rect 256602 335316 256608 335368
rect 256660 335356 256666 335368
rect 257062 335356 257068 335368
rect 256660 335328 257068 335356
rect 256660 335316 256666 335328
rect 257062 335316 257068 335328
rect 257120 335316 257126 335368
rect 258350 335316 258356 335368
rect 258408 335356 258414 335368
rect 258718 335356 258724 335368
rect 258408 335328 258724 335356
rect 258408 335316 258414 335328
rect 258718 335316 258724 335328
rect 258776 335316 258782 335368
rect 259196 335356 259224 335464
rect 259546 335452 259552 335464
rect 259604 335452 259610 335504
rect 259822 335452 259828 335504
rect 259880 335492 259886 335504
rect 260466 335492 260472 335504
rect 259880 335464 260472 335492
rect 259880 335452 259886 335464
rect 260466 335452 260472 335464
rect 260524 335452 260530 335504
rect 259270 335384 259276 335436
rect 259328 335424 259334 335436
rect 260006 335424 260012 335436
rect 259328 335396 260012 335424
rect 259328 335384 259334 335396
rect 260006 335384 260012 335396
rect 260064 335384 260070 335436
rect 260834 335384 260840 335436
rect 260892 335424 260898 335436
rect 262122 335424 262128 335436
rect 260892 335396 262128 335424
rect 260892 335384 260898 335396
rect 262122 335384 262128 335396
rect 262180 335384 262186 335436
rect 262490 335384 262496 335436
rect 262548 335424 262554 335436
rect 262858 335424 262864 335436
rect 262548 335396 262864 335424
rect 262548 335384 262554 335396
rect 262858 335384 262864 335396
rect 262916 335384 262922 335436
rect 263382 335424 263410 335532
rect 264514 335520 264520 335572
rect 264572 335560 264578 335572
rect 264572 335532 267136 335560
rect 264572 335520 264578 335532
rect 266906 335492 266912 335504
rect 263750 335464 266912 335492
rect 263750 335424 263778 335464
rect 266906 335452 266912 335464
rect 266964 335452 266970 335504
rect 263382 335396 263778 335424
rect 264238 335384 264244 335436
rect 264296 335424 264302 335436
rect 264698 335424 264704 335436
rect 264296 335396 264704 335424
rect 264296 335384 264302 335396
rect 264698 335384 264704 335396
rect 264756 335384 264762 335436
rect 266354 335384 266360 335436
rect 266412 335424 266418 335436
rect 267108 335424 267136 335532
rect 267182 335520 267188 335572
rect 267240 335560 267246 335572
rect 268470 335560 268476 335572
rect 267240 335532 268476 335560
rect 267240 335520 267246 335532
rect 268470 335520 268476 335532
rect 268528 335520 268534 335572
rect 268562 335520 268568 335572
rect 268620 335560 268626 335572
rect 268933 335563 268991 335569
rect 268933 335560 268945 335563
rect 268620 335532 268945 335560
rect 268620 335520 268626 335532
rect 268933 335529 268945 335532
rect 268979 335529 268991 335563
rect 268933 335523 268991 335529
rect 269114 335520 269120 335572
rect 269172 335560 269178 335572
rect 269482 335560 269488 335572
rect 269172 335532 269488 335560
rect 269172 335520 269178 335532
rect 269482 335520 269488 335532
rect 269540 335520 269546 335572
rect 269850 335560 269856 335572
rect 269638 335532 269856 335560
rect 269206 335452 269212 335504
rect 269264 335492 269270 335504
rect 269638 335492 269666 335532
rect 269850 335520 269856 335532
rect 269908 335520 269914 335572
rect 269264 335464 269666 335492
rect 269264 335452 269270 335464
rect 266412 335396 267044 335424
rect 267108 335396 268516 335424
rect 266412 335384 266418 335396
rect 259104 335328 259224 335356
rect 259104 335300 259132 335328
rect 259914 335316 259920 335368
rect 259972 335356 259978 335368
rect 260374 335356 260380 335368
rect 259972 335328 260380 335356
rect 259972 335316 259978 335328
rect 260374 335316 260380 335328
rect 260432 335316 260438 335368
rect 260650 335356 260656 335368
rect 260484 335328 260656 335356
rect 219342 335248 219348 335300
rect 219400 335288 219406 335300
rect 253198 335288 253204 335300
rect 219400 335260 253204 335288
rect 219400 335248 219406 335260
rect 253198 335248 253204 335260
rect 253256 335248 253262 335300
rect 259086 335248 259092 335300
rect 259144 335248 259150 335300
rect 259270 335288 259276 335300
rect 259231 335260 259276 335288
rect 259270 335248 259276 335260
rect 259328 335248 259334 335300
rect 259822 335248 259828 335300
rect 259880 335288 259886 335300
rect 260484 335288 260512 335328
rect 260650 335316 260656 335328
rect 260708 335316 260714 335368
rect 261294 335316 261300 335368
rect 261352 335356 261358 335368
rect 261570 335356 261576 335368
rect 261352 335328 261576 335356
rect 261352 335316 261358 335328
rect 261570 335316 261576 335328
rect 261628 335316 261634 335368
rect 262582 335316 262588 335368
rect 262640 335356 262646 335368
rect 262950 335356 262956 335368
rect 262640 335328 262956 335356
rect 262640 335316 262646 335328
rect 262950 335316 262956 335328
rect 263008 335316 263014 335368
rect 263134 335316 263140 335368
rect 263192 335356 263198 335368
rect 263410 335356 263416 335368
rect 263192 335328 263416 335356
rect 263192 335316 263198 335328
rect 263410 335316 263416 335328
rect 263468 335316 263474 335368
rect 263505 335359 263563 335365
rect 263505 335325 263517 335359
rect 263551 335356 263563 335359
rect 263686 335356 263692 335368
rect 263551 335328 263692 335356
rect 263551 335325 263563 335328
rect 263505 335319 263563 335325
rect 263686 335316 263692 335328
rect 263744 335316 263750 335368
rect 264606 335316 264612 335368
rect 264664 335356 264670 335368
rect 264882 335356 264888 335368
rect 264664 335328 264888 335356
rect 264664 335316 264670 335328
rect 264882 335316 264888 335328
rect 264940 335316 264946 335368
rect 264974 335316 264980 335368
rect 265032 335356 265038 335368
rect 265894 335356 265900 335368
rect 265032 335328 265900 335356
rect 265032 335316 265038 335328
rect 265894 335316 265900 335328
rect 265952 335316 265958 335368
rect 266630 335316 266636 335368
rect 266688 335356 266694 335368
rect 266814 335356 266820 335368
rect 266688 335328 266820 335356
rect 266688 335316 266694 335328
rect 266814 335316 266820 335328
rect 266872 335316 266878 335368
rect 259880 335260 260512 335288
rect 267016 335288 267044 335396
rect 267090 335316 267096 335368
rect 267148 335356 267154 335368
rect 267550 335356 267556 335368
rect 267148 335328 267556 335356
rect 267148 335316 267154 335328
rect 267550 335316 267556 335328
rect 267608 335316 267614 335368
rect 267918 335316 267924 335368
rect 267976 335356 267982 335368
rect 268378 335356 268384 335368
rect 267976 335328 268384 335356
rect 267976 335316 267982 335328
rect 268378 335316 268384 335328
rect 268436 335316 268442 335368
rect 268488 335356 268516 335396
rect 268562 335384 268568 335436
rect 268620 335424 268626 335436
rect 269022 335424 269028 335436
rect 268620 335396 269028 335424
rect 268620 335384 268626 335396
rect 269022 335384 269028 335396
rect 269080 335384 269086 335436
rect 269298 335384 269304 335436
rect 269356 335424 269362 335436
rect 269850 335424 269856 335436
rect 269356 335396 269856 335424
rect 269356 335384 269362 335396
rect 269850 335384 269856 335396
rect 269908 335384 269914 335436
rect 270034 335384 270040 335436
rect 270092 335424 270098 335436
rect 270402 335424 270408 335436
rect 270092 335396 270408 335424
rect 270092 335384 270098 335396
rect 270402 335384 270408 335396
rect 270460 335384 270466 335436
rect 270512 335424 270540 335668
rect 271046 335656 271052 335708
rect 271104 335696 271110 335708
rect 271693 335699 271751 335705
rect 271693 335696 271705 335699
rect 271104 335668 271705 335696
rect 271104 335656 271110 335668
rect 271693 335665 271705 335668
rect 271739 335665 271751 335699
rect 271693 335659 271751 335665
rect 270681 335563 270739 335569
rect 270681 335529 270693 335563
rect 270727 335560 270739 335563
rect 272061 335563 272119 335569
rect 270727 335532 271920 335560
rect 270727 335529 270739 335532
rect 270681 335523 270739 335529
rect 271322 335424 271328 335436
rect 270512 335396 271328 335424
rect 271322 335384 271328 335396
rect 271380 335384 271386 335436
rect 271892 335424 271920 335532
rect 272061 335529 272073 335563
rect 272107 335560 272119 335563
rect 273226 335560 273254 335804
rect 277210 335764 277216 335776
rect 277171 335736 277216 335764
rect 277210 335724 277216 335736
rect 277268 335724 277274 335776
rect 278866 335724 278872 335776
rect 278924 335764 278930 335776
rect 280062 335764 280068 335776
rect 278924 335736 280068 335764
rect 278924 335724 278930 335736
rect 280062 335724 280068 335736
rect 280120 335724 280126 335776
rect 280614 335724 280620 335776
rect 280672 335764 280678 335776
rect 281442 335764 281448 335776
rect 280672 335736 281448 335764
rect 280672 335724 280678 335736
rect 281442 335724 281448 335736
rect 281500 335724 281506 335776
rect 281994 335724 282000 335776
rect 282052 335764 282058 335776
rect 282638 335764 282644 335776
rect 282052 335736 282644 335764
rect 282052 335724 282058 335736
rect 282638 335724 282644 335736
rect 282696 335724 282702 335776
rect 280525 335699 280583 335705
rect 278148 335668 278590 335696
rect 273714 335588 273720 335640
rect 273772 335628 273778 335640
rect 278148 335628 278176 335668
rect 273772 335600 278176 335628
rect 273772 335588 273778 335600
rect 272107 335532 273254 335560
rect 272107 335529 272119 335532
rect 272061 335523 272119 335529
rect 273622 335520 273628 335572
rect 273680 335560 273686 335572
rect 274174 335560 274180 335572
rect 273680 335532 274180 335560
rect 273680 335520 273686 335532
rect 274174 335520 274180 335532
rect 274232 335520 274238 335572
rect 275002 335520 275008 335572
rect 275060 335560 275066 335572
rect 275554 335560 275560 335572
rect 275060 335532 275560 335560
rect 275060 335520 275066 335532
rect 275554 335520 275560 335532
rect 275612 335520 275618 335572
rect 277394 335520 277400 335572
rect 277452 335560 277458 335572
rect 278314 335560 278320 335572
rect 277452 335532 278320 335560
rect 277452 335520 277458 335532
rect 278314 335520 278320 335532
rect 278372 335520 278378 335572
rect 278562 335560 278590 335668
rect 280525 335665 280537 335699
rect 280571 335696 280583 335699
rect 281166 335696 281172 335708
rect 280571 335668 281172 335696
rect 280571 335665 280583 335668
rect 280525 335659 280583 335665
rect 281166 335656 281172 335668
rect 281224 335656 281230 335708
rect 282886 335696 282914 335804
rect 283101 335801 283113 335835
rect 283147 335832 283159 335835
rect 286505 335835 286563 335841
rect 286505 335832 286517 335835
rect 283147 335804 286517 335832
rect 283147 335801 283159 335804
rect 283101 335795 283159 335801
rect 286505 335801 286517 335804
rect 286551 335801 286563 335835
rect 286505 335795 286563 335801
rect 287514 335792 287520 335844
rect 287572 335832 287578 335844
rect 288158 335832 288164 335844
rect 287572 335804 288164 335832
rect 287572 335792 287578 335804
rect 288158 335792 288164 335804
rect 288216 335792 288222 335844
rect 289078 335764 289084 335776
rect 283024 335736 289084 335764
rect 283024 335696 283052 335736
rect 289078 335724 289084 335736
rect 289136 335724 289142 335776
rect 282886 335668 283052 335696
rect 284757 335699 284815 335705
rect 284757 335665 284769 335699
rect 284803 335696 284815 335699
rect 289170 335696 289176 335708
rect 284803 335668 289176 335696
rect 284803 335665 284815 335668
rect 284757 335659 284815 335665
rect 289170 335656 289176 335668
rect 289228 335656 289234 335708
rect 279142 335588 279148 335640
rect 279200 335628 279206 335640
rect 282638 335628 282644 335640
rect 279200 335600 282644 335628
rect 279200 335588 279206 335600
rect 282638 335588 282644 335600
rect 282696 335588 282702 335640
rect 282733 335631 282791 335637
rect 282733 335597 282745 335631
rect 282779 335628 282791 335631
rect 282917 335631 282975 335637
rect 282917 335628 282929 335631
rect 282779 335600 282929 335628
rect 282779 335597 282791 335600
rect 282733 335591 282791 335597
rect 282917 335597 282929 335600
rect 282963 335597 282975 335631
rect 282917 335591 282975 335597
rect 283006 335588 283012 335640
rect 283064 335628 283070 335640
rect 286410 335628 286416 335640
rect 283064 335600 286416 335628
rect 283064 335588 283070 335600
rect 286410 335588 286416 335600
rect 286468 335588 286474 335640
rect 286505 335631 286563 335637
rect 286505 335597 286517 335631
rect 286551 335628 286563 335631
rect 289262 335628 289268 335640
rect 286551 335600 289268 335628
rect 286551 335597 286563 335600
rect 286505 335591 286563 335597
rect 289262 335588 289268 335600
rect 289320 335588 289326 335640
rect 284757 335563 284815 335569
rect 284757 335560 284769 335563
rect 278562 335532 284769 335560
rect 284757 335529 284769 335532
rect 284803 335529 284815 335563
rect 284757 335523 284815 335529
rect 284846 335520 284852 335572
rect 284904 335560 284910 335572
rect 285398 335560 285404 335572
rect 284904 335532 285404 335560
rect 284904 335520 284910 335532
rect 285398 335520 285404 335532
rect 285456 335520 285462 335572
rect 287333 335563 287391 335569
rect 287333 335529 287345 335563
rect 287379 335560 287391 335563
rect 291838 335560 291844 335572
rect 287379 335532 291844 335560
rect 287379 335529 287391 335532
rect 287333 335523 287391 335529
rect 291838 335520 291844 335532
rect 291896 335520 291902 335572
rect 271969 335495 272027 335501
rect 271969 335461 271981 335495
rect 272015 335492 272027 335495
rect 292546 335492 292574 335872
rect 296070 335860 296076 335872
rect 296128 335860 296134 335912
rect 272015 335464 292574 335492
rect 272015 335461 272027 335464
rect 271969 335455 272027 335461
rect 282733 335427 282791 335433
rect 282733 335424 282745 335427
rect 271892 335396 282745 335424
rect 282733 335393 282745 335396
rect 282779 335393 282791 335427
rect 282733 335387 282791 335393
rect 282825 335427 282883 335433
rect 282825 335393 282837 335427
rect 282871 335424 282883 335427
rect 284297 335427 284355 335433
rect 284297 335424 284309 335427
rect 282871 335396 284309 335424
rect 282871 335393 282883 335396
rect 282825 335387 282883 335393
rect 284297 335393 284309 335396
rect 284343 335393 284355 335427
rect 284297 335387 284355 335393
rect 284386 335384 284392 335436
rect 284444 335424 284450 335436
rect 285306 335424 285312 335436
rect 284444 335396 285312 335424
rect 284444 335384 284450 335396
rect 285306 335384 285312 335396
rect 285364 335384 285370 335436
rect 285401 335427 285459 335433
rect 285401 335393 285413 335427
rect 285447 335424 285459 335427
rect 291930 335424 291936 335436
rect 285447 335396 291936 335424
rect 285447 335393 285459 335396
rect 285401 335387 285459 335393
rect 291930 335384 291936 335396
rect 291988 335384 291994 335436
rect 268488 335328 268700 335356
rect 267366 335288 267372 335300
rect 267016 335260 267372 335288
rect 259880 335248 259886 335260
rect 267366 335248 267372 335260
rect 267424 335248 267430 335300
rect 201402 335180 201408 335232
rect 201460 335220 201466 335232
rect 251910 335220 251916 335232
rect 201460 335192 251916 335220
rect 201460 335180 201466 335192
rect 251910 335180 251916 335192
rect 251968 335180 251974 335232
rect 268672 335220 268700 335328
rect 268746 335316 268752 335368
rect 268804 335356 268810 335368
rect 268930 335356 268936 335368
rect 268804 335328 268936 335356
rect 268804 335316 268810 335328
rect 268930 335316 268936 335328
rect 268988 335316 268994 335368
rect 269390 335316 269396 335368
rect 269448 335356 269454 335368
rect 269666 335356 269672 335368
rect 269448 335328 269672 335356
rect 269448 335316 269454 335328
rect 269666 335316 269672 335328
rect 269724 335316 269730 335368
rect 270313 335359 270371 335365
rect 270313 335325 270325 335359
rect 270359 335356 270371 335359
rect 270359 335328 271000 335356
rect 270359 335325 270371 335328
rect 270313 335319 270371 335325
rect 269853 335291 269911 335297
rect 269853 335288 269865 335291
rect 269776 335260 269865 335288
rect 269776 335220 269804 335260
rect 269853 335257 269865 335260
rect 269899 335257 269911 335291
rect 270972 335288 271000 335328
rect 271046 335316 271052 335368
rect 271104 335356 271110 335368
rect 271690 335356 271696 335368
rect 271104 335328 271696 335356
rect 271104 335316 271110 335328
rect 271690 335316 271696 335328
rect 271748 335316 271754 335368
rect 271966 335316 271972 335368
rect 272024 335356 272030 335368
rect 272334 335356 272340 335368
rect 272024 335328 272340 335356
rect 272024 335316 272030 335328
rect 272334 335316 272340 335328
rect 272392 335316 272398 335368
rect 272610 335316 272616 335368
rect 272668 335356 272674 335368
rect 273070 335356 273076 335368
rect 272668 335328 273076 335356
rect 272668 335316 272674 335328
rect 273070 335316 273076 335328
rect 273128 335316 273134 335368
rect 273530 335316 273536 335368
rect 273588 335356 273594 335368
rect 273588 335328 273944 335356
rect 273588 335316 273594 335328
rect 271598 335288 271604 335300
rect 270972 335260 271604 335288
rect 269853 335251 269911 335257
rect 271598 335248 271604 335260
rect 271656 335248 271662 335300
rect 273916 335288 273944 335328
rect 273990 335316 273996 335368
rect 274048 335356 274054 335368
rect 274266 335356 274272 335368
rect 274048 335328 274272 335356
rect 274048 335316 274054 335328
rect 274266 335316 274272 335328
rect 274324 335316 274330 335368
rect 275462 335316 275468 335368
rect 275520 335356 275526 335368
rect 275922 335356 275928 335368
rect 275520 335328 275928 335356
rect 275520 335316 275526 335328
rect 275922 335316 275928 335328
rect 275980 335316 275986 335368
rect 276934 335356 276940 335368
rect 276895 335328 276940 335356
rect 276934 335316 276940 335328
rect 276992 335316 276998 335368
rect 277026 335316 277032 335368
rect 277084 335356 277090 335368
rect 277302 335356 277308 335368
rect 277084 335328 277308 335356
rect 277084 335316 277090 335328
rect 277302 335316 277308 335328
rect 277360 335316 277366 335368
rect 277486 335316 277492 335368
rect 277544 335356 277550 335368
rect 277946 335356 277952 335368
rect 277544 335328 277952 335356
rect 277544 335316 277550 335328
rect 277946 335316 277952 335328
rect 278004 335316 278010 335368
rect 279418 335316 279424 335368
rect 279476 335356 279482 335368
rect 279878 335356 279884 335368
rect 279476 335328 279884 335356
rect 279476 335316 279482 335328
rect 279878 335316 279884 335328
rect 279936 335316 279942 335368
rect 280154 335316 280160 335368
rect 280212 335356 280218 335368
rect 280212 335328 280568 335356
rect 280212 335316 280218 335328
rect 274174 335288 274180 335300
rect 273916 335260 274180 335288
rect 274174 335248 274180 335260
rect 274232 335248 274238 335300
rect 274726 335248 274732 335300
rect 274784 335288 274790 335300
rect 275281 335291 275339 335297
rect 275281 335288 275293 335291
rect 274784 335260 275293 335288
rect 274784 335248 274790 335260
rect 275281 335257 275293 335260
rect 275327 335257 275339 335291
rect 280540 335288 280568 335328
rect 281718 335316 281724 335368
rect 281776 335356 281782 335368
rect 282178 335356 282184 335368
rect 281776 335328 282184 335356
rect 281776 335316 281782 335328
rect 282178 335316 282184 335328
rect 282236 335316 282242 335368
rect 282917 335359 282975 335365
rect 282917 335356 282929 335359
rect 282288 335328 282929 335356
rect 281350 335288 281356 335300
rect 280540 335260 281356 335288
rect 275281 335251 275339 335257
rect 281350 335248 281356 335260
rect 281408 335248 281414 335300
rect 269942 335220 269948 335232
rect 268672 335192 269804 335220
rect 269903 335192 269948 335220
rect 269942 335180 269948 335192
rect 270000 335180 270006 335232
rect 277302 335220 277308 335232
rect 277263 335192 277308 335220
rect 277302 335180 277308 335192
rect 277360 335180 277366 335232
rect 277397 335223 277455 335229
rect 277397 335189 277409 335223
rect 277443 335220 277455 335223
rect 282288 335220 282316 335328
rect 282917 335325 282929 335328
rect 282963 335325 282975 335359
rect 282917 335319 282975 335325
rect 283006 335316 283012 335368
rect 283064 335356 283070 335368
rect 283558 335356 283564 335368
rect 283064 335328 283564 335356
rect 283064 335316 283070 335328
rect 283558 335316 283564 335328
rect 283616 335316 283622 335368
rect 284018 335316 284024 335368
rect 284076 335356 284082 335368
rect 284202 335356 284208 335368
rect 284076 335328 284208 335356
rect 284076 335316 284082 335328
rect 284202 335316 284208 335328
rect 284260 335316 284266 335368
rect 284478 335316 284484 335368
rect 284536 335356 284542 335368
rect 284846 335356 284852 335368
rect 284536 335328 284852 335356
rect 284536 335316 284542 335328
rect 284846 335316 284852 335328
rect 284904 335316 284910 335368
rect 285030 335316 285036 335368
rect 285088 335356 285094 335368
rect 285490 335356 285496 335368
rect 285088 335328 285496 335356
rect 285088 335316 285094 335328
rect 285490 335316 285496 335328
rect 285548 335316 285554 335368
rect 285585 335359 285643 335365
rect 285585 335325 285597 335359
rect 285631 335356 285643 335359
rect 290458 335356 290464 335368
rect 285631 335328 290464 335356
rect 285631 335325 285643 335328
rect 285585 335319 285643 335325
rect 290458 335316 290464 335328
rect 290516 335316 290522 335368
rect 282365 335291 282423 335297
rect 282365 335257 282377 335291
rect 282411 335288 282423 335291
rect 396718 335288 396724 335300
rect 282411 335260 396724 335288
rect 282411 335257 282423 335260
rect 282365 335251 282423 335257
rect 396718 335248 396724 335260
rect 396776 335248 396782 335300
rect 403618 335220 403624 335232
rect 277443 335192 282316 335220
rect 282380 335192 403624 335220
rect 277443 335189 277455 335192
rect 277397 335183 277455 335189
rect 194410 335112 194416 335164
rect 194468 335152 194474 335164
rect 245102 335152 245108 335164
rect 194468 335124 245108 335152
rect 194468 335112 194474 335124
rect 245102 335112 245108 335124
rect 245160 335112 245166 335164
rect 268930 335152 268936 335164
rect 268891 335124 268936 335152
rect 268930 335112 268936 335124
rect 268988 335112 268994 335164
rect 270037 335155 270095 335161
rect 270037 335121 270049 335155
rect 270083 335152 270095 335155
rect 270218 335152 270224 335164
rect 270083 335124 270224 335152
rect 270083 335121 270095 335124
rect 270037 335115 270095 335121
rect 270218 335112 270224 335124
rect 270276 335112 270282 335164
rect 276658 335112 276664 335164
rect 276716 335152 276722 335164
rect 279418 335152 279424 335164
rect 276716 335124 279424 335152
rect 276716 335112 276722 335124
rect 279418 335112 279424 335124
rect 279476 335112 279482 335164
rect 279513 335155 279571 335161
rect 279513 335121 279525 335155
rect 279559 335152 279571 335155
rect 282380 335152 282408 335192
rect 403618 335180 403624 335192
rect 403676 335180 403682 335232
rect 279559 335124 282408 335152
rect 282457 335155 282515 335161
rect 279559 335121 279571 335124
rect 279513 335115 279571 335121
rect 282457 335121 282469 335155
rect 282503 335152 282515 335155
rect 433978 335152 433984 335164
rect 282503 335124 433984 335152
rect 282503 335121 282515 335124
rect 282457 335115 282515 335121
rect 433978 335112 433984 335124
rect 434036 335112 434042 335164
rect 197262 335044 197268 335096
rect 197320 335084 197326 335096
rect 251542 335084 251548 335096
rect 197320 335056 251548 335084
rect 197320 335044 197326 335056
rect 251542 335044 251548 335056
rect 251600 335044 251606 335096
rect 269482 335044 269488 335096
rect 269540 335084 269546 335096
rect 405734 335084 405740 335096
rect 269540 335056 405740 335084
rect 269540 335044 269546 335056
rect 405734 335044 405740 335056
rect 405792 335044 405798 335096
rect 190362 334976 190368 335028
rect 190420 335016 190426 335028
rect 250898 335016 250904 335028
rect 190420 334988 250904 335016
rect 190420 334976 190426 334988
rect 250898 334976 250904 334988
rect 250956 334976 250962 335028
rect 277854 334976 277860 335028
rect 277912 335016 277918 335028
rect 278314 335016 278320 335028
rect 277912 334988 278320 335016
rect 277912 334976 277918 334988
rect 278314 334976 278320 334988
rect 278372 334976 278378 335028
rect 278682 334976 278688 335028
rect 278740 335016 278746 335028
rect 434070 335016 434076 335028
rect 278740 334988 434076 335016
rect 278740 334976 278746 334988
rect 434070 334976 434076 334988
rect 434128 334976 434134 335028
rect 186130 334908 186136 334960
rect 186188 334948 186194 334960
rect 245838 334948 245844 334960
rect 186188 334920 245844 334948
rect 186188 334908 186194 334920
rect 245838 334908 245844 334920
rect 245896 334908 245902 334960
rect 278777 334951 278835 334957
rect 278777 334917 278789 334951
rect 278823 334948 278835 334951
rect 282457 334951 282515 334957
rect 282457 334948 282469 334951
rect 278823 334920 282469 334948
rect 278823 334917 278835 334920
rect 278777 334911 278835 334917
rect 282457 334917 282469 334920
rect 282503 334917 282515 334951
rect 282457 334911 282515 334917
rect 282549 334951 282607 334957
rect 282549 334917 282561 334951
rect 282595 334948 282607 334951
rect 434162 334948 434168 334960
rect 282595 334920 434168 334948
rect 282595 334917 282607 334920
rect 282549 334911 282607 334917
rect 434162 334908 434168 334920
rect 434220 334908 434226 334960
rect 183462 334840 183468 334892
rect 183520 334880 183526 334892
rect 250349 334883 250407 334889
rect 250349 334880 250361 334883
rect 183520 334852 250361 334880
rect 183520 334840 183526 334852
rect 250349 334849 250361 334852
rect 250395 334849 250407 334883
rect 250349 334843 250407 334849
rect 272058 334840 272064 334892
rect 272116 334880 272122 334892
rect 437474 334880 437480 334892
rect 272116 334852 437480 334880
rect 272116 334840 272122 334852
rect 437474 334840 437480 334852
rect 437532 334840 437538 334892
rect 179322 334772 179328 334824
rect 179380 334812 179386 334824
rect 250073 334815 250131 334821
rect 250073 334812 250085 334815
rect 179380 334784 250085 334812
rect 179380 334772 179386 334784
rect 250073 334781 250085 334784
rect 250119 334781 250131 334815
rect 250073 334775 250131 334781
rect 251358 334772 251364 334824
rect 251416 334812 251422 334824
rect 252462 334812 252468 334824
rect 251416 334784 252468 334812
rect 251416 334772 251422 334784
rect 252462 334772 252468 334784
rect 252520 334772 252526 334824
rect 273809 334815 273867 334821
rect 273809 334781 273821 334815
rect 273855 334812 273867 334815
rect 275833 334815 275891 334821
rect 273855 334784 274036 334812
rect 273855 334781 273867 334784
rect 273809 334775 273867 334781
rect 169570 334704 169576 334756
rect 169628 334744 169634 334756
rect 244274 334744 244280 334756
rect 169628 334716 244280 334744
rect 169628 334704 169634 334716
rect 244274 334704 244280 334716
rect 244332 334704 244338 334756
rect 245102 334704 245108 334756
rect 245160 334744 245166 334756
rect 254946 334744 254952 334756
rect 245160 334716 254952 334744
rect 245160 334704 245166 334716
rect 254946 334704 254952 334716
rect 255004 334704 255010 334756
rect 271874 334704 271880 334756
rect 271932 334744 271938 334756
rect 272058 334744 272064 334756
rect 271932 334716 272064 334744
rect 271932 334704 271938 334716
rect 272058 334704 272064 334716
rect 272116 334704 272122 334756
rect 274008 334744 274036 334784
rect 275833 334781 275845 334815
rect 275879 334812 275891 334815
rect 280525 334815 280583 334821
rect 275879 334784 280476 334812
rect 275879 334781 275891 334784
rect 275833 334775 275891 334781
rect 280062 334744 280068 334756
rect 274008 334716 280068 334744
rect 280062 334704 280068 334716
rect 280120 334704 280126 334756
rect 165522 334636 165528 334688
rect 165580 334676 165586 334688
rect 238941 334679 238999 334685
rect 238941 334676 238953 334679
rect 165580 334648 238953 334676
rect 165580 334636 165586 334648
rect 238941 334645 238953 334648
rect 238987 334645 238999 334679
rect 247402 334676 247408 334688
rect 238941 334639 238999 334645
rect 241486 334648 247408 334676
rect 158622 334568 158628 334620
rect 158680 334608 158686 334620
rect 241486 334608 241514 334648
rect 247402 334636 247408 334648
rect 247460 334636 247466 334688
rect 268194 334636 268200 334688
rect 268252 334676 268258 334688
rect 273717 334679 273775 334685
rect 273717 334676 273729 334679
rect 268252 334648 273729 334676
rect 268252 334636 268258 334648
rect 273717 334645 273729 334648
rect 273763 334645 273775 334679
rect 273717 334639 273775 334645
rect 273993 334679 274051 334685
rect 273993 334645 274005 334679
rect 274039 334676 274051 334679
rect 280154 334676 280160 334688
rect 274039 334648 280160 334676
rect 274039 334645 274051 334648
rect 273993 334639 274051 334645
rect 280154 334636 280160 334648
rect 280212 334636 280218 334688
rect 280448 334676 280476 334784
rect 280525 334781 280537 334815
rect 280571 334812 280583 334815
rect 536834 334812 536840 334824
rect 280571 334784 536840 334812
rect 280571 334781 280583 334784
rect 280525 334775 280583 334781
rect 536834 334772 536840 334784
rect 536892 334772 536898 334824
rect 280709 334747 280767 334753
rect 280709 334713 280721 334747
rect 280755 334744 280767 334747
rect 539594 334744 539600 334756
rect 280755 334716 539600 334744
rect 280755 334713 280767 334716
rect 280709 334707 280767 334713
rect 539594 334704 539600 334716
rect 539652 334704 539658 334756
rect 281626 334676 281632 334688
rect 280448 334648 281632 334676
rect 281626 334636 281632 334648
rect 281684 334636 281690 334688
rect 281810 334636 281816 334688
rect 281868 334676 281874 334688
rect 550634 334676 550640 334688
rect 281868 334648 550640 334676
rect 281868 334636 281874 334648
rect 550634 334636 550640 334648
rect 550692 334636 550698 334688
rect 158680 334580 241514 334608
rect 247221 334611 247279 334617
rect 158680 334568 158686 334580
rect 247221 334577 247233 334611
rect 247267 334608 247279 334611
rect 247586 334608 247592 334620
rect 247267 334580 247592 334608
rect 247267 334577 247279 334580
rect 247221 334571 247279 334577
rect 247586 334568 247592 334580
rect 247644 334568 247650 334620
rect 248782 334568 248788 334620
rect 248840 334608 248846 334620
rect 249426 334608 249432 334620
rect 248840 334580 249432 334608
rect 248840 334568 248846 334580
rect 249426 334568 249432 334580
rect 249484 334568 249490 334620
rect 262214 334568 262220 334620
rect 262272 334608 262278 334620
rect 273809 334611 273867 334617
rect 273809 334608 273821 334611
rect 262272 334580 273821 334608
rect 262272 334568 262278 334580
rect 273809 334577 273821 334580
rect 273855 334577 273867 334611
rect 273809 334571 273867 334577
rect 274085 334611 274143 334617
rect 274085 334577 274097 334611
rect 274131 334608 274143 334611
rect 280798 334608 280804 334620
rect 274131 334580 280804 334608
rect 274131 334577 274143 334580
rect 274085 334571 274143 334577
rect 280798 334568 280804 334580
rect 280856 334568 280862 334620
rect 281997 334611 282055 334617
rect 281997 334577 282009 334611
rect 282043 334608 282055 334611
rect 554774 334608 554780 334620
rect 282043 334580 554780 334608
rect 282043 334577 282055 334580
rect 281997 334571 282055 334577
rect 554774 334568 554780 334580
rect 554832 334568 554838 334620
rect 204162 334500 204168 334552
rect 204220 334540 204226 334552
rect 204220 334512 244274 334540
rect 204220 334500 204226 334512
rect 211062 334432 211068 334484
rect 211120 334472 211126 334484
rect 238849 334475 238907 334481
rect 238849 334472 238861 334475
rect 211120 334444 238861 334472
rect 211120 334432 211126 334444
rect 238849 334441 238861 334444
rect 238895 334441 238907 334475
rect 238849 334435 238907 334441
rect 238941 334475 238999 334481
rect 238941 334441 238953 334475
rect 238987 334472 238999 334475
rect 244093 334475 244151 334481
rect 244093 334472 244105 334475
rect 238987 334444 244105 334472
rect 238987 334441 238999 334444
rect 238941 334435 238999 334441
rect 244093 334441 244105 334444
rect 244139 334441 244151 334475
rect 244246 334472 244274 334512
rect 267826 334500 267832 334552
rect 267884 334540 267890 334552
rect 387794 334540 387800 334552
rect 267884 334512 387800 334540
rect 267884 334500 267890 334512
rect 387794 334500 387800 334512
rect 387852 334500 387858 334552
rect 252094 334472 252100 334484
rect 244246 334444 252100 334472
rect 244093 334435 244151 334441
rect 252094 334432 252100 334444
rect 252152 334432 252158 334484
rect 262214 334472 262220 334484
rect 262175 334444 262220 334472
rect 262214 334432 262220 334444
rect 262272 334432 262278 334484
rect 270494 334432 270500 334484
rect 270552 334472 270558 334484
rect 270552 334444 273254 334472
rect 270552 334432 270558 334444
rect 208302 334364 208308 334416
rect 208360 334404 208366 334416
rect 251358 334404 251364 334416
rect 208360 334376 251364 334404
rect 208360 334364 208366 334376
rect 251358 334364 251364 334376
rect 251416 334364 251422 334416
rect 251910 334364 251916 334416
rect 251968 334404 251974 334416
rect 255406 334404 255412 334416
rect 251968 334376 255412 334404
rect 251968 334364 251974 334376
rect 255406 334364 255412 334376
rect 255464 334364 255470 334416
rect 273226 334404 273254 334444
rect 277578 334432 277584 334484
rect 277636 334472 277642 334484
rect 282549 334475 282607 334481
rect 282549 334472 282561 334475
rect 277636 334444 282561 334472
rect 277636 334432 277642 334444
rect 282549 334441 282561 334444
rect 282595 334441 282607 334475
rect 282549 334435 282607 334441
rect 282638 334432 282644 334484
rect 282696 334472 282702 334484
rect 393958 334472 393964 334484
rect 282696 334444 393964 334472
rect 282696 334432 282702 334444
rect 393958 334432 393964 334444
rect 394016 334432 394022 334484
rect 325694 334404 325700 334416
rect 273226 334376 325700 334404
rect 325694 334364 325700 334376
rect 325752 334364 325758 334416
rect 222102 334296 222108 334348
rect 222160 334336 222166 334348
rect 253658 334336 253664 334348
rect 222160 334308 253664 334336
rect 222160 334296 222166 334308
rect 253658 334296 253664 334308
rect 253716 334296 253722 334348
rect 274542 334296 274548 334348
rect 274600 334336 274606 334348
rect 276658 334336 276664 334348
rect 274600 334308 276664 334336
rect 274600 334296 274606 334308
rect 276658 334296 276664 334308
rect 276716 334296 276722 334348
rect 276842 334296 276848 334348
rect 276900 334336 276906 334348
rect 282365 334339 282423 334345
rect 282365 334336 282377 334339
rect 276900 334308 282377 334336
rect 276900 334296 276906 334308
rect 282365 334305 282377 334308
rect 282411 334305 282423 334339
rect 282365 334299 282423 334305
rect 282641 334339 282699 334345
rect 282641 334305 282653 334339
rect 282687 334336 282699 334339
rect 391198 334336 391204 334348
rect 282687 334308 391204 334336
rect 282687 334305 282699 334308
rect 282641 334299 282699 334305
rect 391198 334296 391204 334308
rect 391256 334296 391262 334348
rect 215202 334228 215208 334280
rect 215260 334268 215266 334280
rect 238757 334271 238815 334277
rect 238757 334268 238769 334271
rect 215260 334240 238769 334268
rect 215260 334228 215266 334240
rect 238757 334237 238769 334240
rect 238803 334237 238815 334271
rect 238757 334231 238815 334237
rect 238849 334271 238907 334277
rect 238849 334237 238861 334271
rect 238895 334268 238907 334271
rect 241698 334268 241704 334280
rect 238895 334240 241704 334268
rect 238895 334237 238907 334240
rect 238849 334231 238907 334237
rect 241698 334228 241704 334240
rect 241756 334228 241762 334280
rect 261202 334228 261208 334280
rect 261260 334268 261266 334280
rect 309134 334268 309140 334280
rect 261260 334240 309140 334268
rect 261260 334228 261266 334240
rect 309134 334228 309140 334240
rect 309192 334228 309198 334280
rect 229002 334160 229008 334212
rect 229060 334200 229066 334212
rect 249150 334200 249156 334212
rect 229060 334172 249156 334200
rect 229060 334160 229066 334172
rect 249150 334160 249156 334172
rect 249208 334160 249214 334212
rect 264146 334160 264152 334212
rect 264204 334200 264210 334212
rect 292574 334200 292580 334212
rect 264204 334172 292580 334200
rect 264204 334160 264210 334172
rect 292574 334160 292580 334172
rect 292632 334160 292638 334212
rect 226242 334092 226248 334144
rect 226300 334132 226306 334144
rect 245562 334132 245568 334144
rect 226300 334104 245568 334132
rect 226300 334092 226306 334104
rect 245562 334092 245568 334104
rect 245620 334092 245626 334144
rect 253566 334092 253572 334144
rect 253624 334132 253630 334144
rect 253750 334132 253756 334144
rect 253624 334104 253756 334132
rect 253624 334092 253630 334104
rect 253750 334092 253756 334104
rect 253808 334092 253814 334144
rect 260282 334092 260288 334144
rect 260340 334132 260346 334144
rect 289354 334132 289360 334144
rect 260340 334104 289360 334132
rect 260340 334092 260346 334104
rect 289354 334092 289360 334104
rect 289412 334092 289418 334144
rect 233970 334024 233976 334076
rect 234028 334064 234034 334076
rect 249518 334064 249524 334076
rect 234028 334036 249524 334064
rect 234028 334024 234034 334036
rect 249518 334024 249524 334036
rect 249576 334024 249582 334076
rect 259362 334024 259368 334076
rect 259420 334064 259426 334076
rect 287698 334064 287704 334076
rect 259420 334036 287704 334064
rect 259420 334024 259426 334036
rect 287698 334024 287704 334036
rect 287756 334024 287762 334076
rect 233878 333956 233884 334008
rect 233936 333996 233942 334008
rect 249705 333999 249763 334005
rect 249705 333996 249717 333999
rect 233936 333968 249717 333996
rect 233936 333956 233942 333968
rect 249705 333965 249717 333968
rect 249751 333965 249763 333999
rect 249705 333959 249763 333965
rect 260561 333999 260619 334005
rect 260561 333965 260573 333999
rect 260607 333996 260619 333999
rect 285030 333996 285036 334008
rect 260607 333968 285036 333996
rect 260607 333965 260619 333968
rect 260561 333959 260619 333965
rect 285030 333956 285036 333968
rect 285088 333956 285094 334008
rect 147582 333888 147588 333940
rect 147640 333928 147646 333940
rect 245933 333931 245991 333937
rect 245933 333928 245945 333931
rect 147640 333900 245945 333928
rect 147640 333888 147646 333900
rect 245933 333897 245945 333900
rect 245979 333897 245991 333931
rect 245933 333891 245991 333897
rect 267645 333931 267703 333937
rect 267645 333897 267657 333931
rect 267691 333928 267703 333931
rect 383654 333928 383660 333940
rect 267691 333900 383660 333928
rect 267691 333897 267703 333900
rect 267645 333891 267703 333897
rect 383654 333888 383660 333900
rect 383712 333888 383718 333940
rect 144730 333820 144736 333872
rect 144788 333860 144794 333872
rect 247218 333860 247224 333872
rect 144788 333832 247224 333860
rect 144788 333820 144794 333832
rect 247218 333820 247224 333832
rect 247276 333820 247282 333872
rect 268930 333820 268936 333872
rect 268988 333860 268994 333872
rect 394694 333860 394700 333872
rect 268988 333832 394700 333860
rect 268988 333820 268994 333832
rect 394694 333820 394700 333832
rect 394752 333820 394758 333872
rect 128262 333752 128268 333804
rect 128320 333792 128326 333804
rect 243722 333792 243728 333804
rect 128320 333764 243728 333792
rect 128320 333752 128326 333764
rect 243722 333752 243728 333764
rect 243780 333752 243786 333804
rect 244918 333792 244924 333804
rect 244879 333764 244924 333792
rect 244918 333752 244924 333764
rect 244976 333752 244982 333804
rect 268654 333752 268660 333804
rect 268712 333792 268718 333804
rect 398834 333792 398840 333804
rect 268712 333764 398840 333792
rect 268712 333752 268718 333764
rect 398834 333752 398840 333764
rect 398892 333752 398898 333804
rect 95142 333684 95148 333736
rect 95200 333724 95206 333736
rect 237006 333724 237012 333736
rect 95200 333696 237012 333724
rect 95200 333684 95206 333696
rect 237006 333684 237012 333696
rect 237064 333684 237070 333736
rect 269114 333684 269120 333736
rect 269172 333724 269178 333736
rect 408494 333724 408500 333736
rect 269172 333696 408500 333724
rect 269172 333684 269178 333696
rect 408494 333684 408500 333696
rect 408552 333684 408558 333736
rect 88242 333616 88248 333668
rect 88300 333656 88306 333668
rect 242434 333656 242440 333668
rect 88300 333628 242440 333656
rect 88300 333616 88306 333628
rect 242434 333616 242440 333628
rect 242492 333616 242498 333668
rect 269206 333616 269212 333668
rect 269264 333656 269270 333668
rect 412634 333656 412640 333668
rect 269264 333628 412640 333656
rect 269264 333616 269270 333628
rect 412634 333616 412640 333628
rect 412692 333616 412698 333668
rect 70302 333548 70308 333600
rect 70360 333588 70366 333600
rect 240870 333588 240876 333600
rect 70360 333560 240876 333588
rect 70360 333548 70366 333560
rect 240870 333548 240876 333560
rect 240928 333548 240934 333600
rect 270405 333591 270463 333597
rect 270405 333557 270417 333591
rect 270451 333588 270463 333591
rect 415394 333588 415400 333600
rect 270451 333560 415400 333588
rect 270451 333557 270463 333560
rect 270405 333551 270463 333557
rect 415394 333548 415400 333560
rect 415452 333548 415458 333600
rect 66162 333480 66168 333532
rect 66220 333520 66226 333532
rect 240413 333523 240471 333529
rect 240413 333520 240425 333523
rect 66220 333492 240425 333520
rect 66220 333480 66226 333492
rect 240413 333489 240425 333492
rect 240459 333489 240471 333523
rect 240413 333483 240471 333489
rect 271049 333523 271107 333529
rect 271049 333489 271061 333523
rect 271095 333520 271107 333523
rect 423674 333520 423680 333532
rect 271095 333492 423680 333520
rect 271095 333489 271107 333492
rect 271049 333483 271107 333489
rect 423674 333480 423680 333492
rect 423732 333480 423738 333532
rect 61930 333412 61936 333464
rect 61988 333452 61994 333464
rect 240226 333452 240232 333464
rect 61988 333424 240232 333452
rect 61988 333412 61994 333424
rect 240226 333412 240232 333424
rect 240284 333412 240290 333464
rect 258077 333455 258135 333461
rect 258077 333421 258089 333455
rect 258123 333452 258135 333455
rect 271417 333455 271475 333461
rect 258123 333424 271000 333452
rect 258123 333421 258135 333424
rect 258077 333415 258135 333421
rect 35894 333344 35900 333396
rect 35952 333384 35958 333396
rect 237926 333384 237932 333396
rect 35952 333356 237932 333384
rect 35952 333344 35958 333356
rect 237926 333344 237932 333356
rect 237984 333344 237990 333396
rect 258166 333344 258172 333396
rect 258224 333384 258230 333396
rect 270862 333384 270868 333396
rect 258224 333356 270868 333384
rect 258224 333344 258230 333356
rect 270862 333344 270868 333356
rect 270920 333344 270926 333396
rect 270972 333384 271000 333424
rect 271417 333421 271429 333455
rect 271463 333452 271475 333455
rect 430574 333452 430580 333464
rect 271463 333424 430580 333452
rect 271463 333421 271475 333424
rect 271417 333415 271475 333421
rect 430574 333412 430580 333424
rect 430632 333412 430638 333464
rect 271598 333384 271604 333396
rect 270972 333356 271604 333384
rect 271598 333344 271604 333356
rect 271656 333344 271662 333396
rect 271693 333387 271751 333393
rect 271693 333353 271705 333387
rect 271739 333384 271751 333387
rect 426434 333384 426440 333396
rect 271739 333356 426440 333384
rect 271739 333353 271751 333356
rect 271693 333347 271751 333353
rect 426434 333344 426440 333356
rect 426492 333344 426498 333396
rect 33134 333276 33140 333328
rect 33192 333316 33198 333328
rect 237742 333316 237748 333328
rect 33192 333288 237748 333316
rect 33192 333276 33198 333288
rect 237742 333276 237748 333288
rect 237800 333276 237806 333328
rect 243262 333276 243268 333328
rect 243320 333316 243326 333328
rect 243725 333319 243783 333325
rect 243725 333316 243737 333319
rect 243320 333288 243737 333316
rect 243320 333276 243326 333288
rect 243725 333285 243737 333288
rect 243771 333285 243783 333319
rect 243725 333279 243783 333285
rect 256970 333276 256976 333328
rect 257028 333316 257034 333328
rect 257982 333316 257988 333328
rect 257028 333288 257988 333316
rect 257028 333276 257034 333288
rect 257982 333276 257988 333288
rect 258040 333276 258046 333328
rect 263962 333276 263968 333328
rect 264020 333316 264026 333328
rect 264514 333316 264520 333328
rect 264020 333288 264520 333316
rect 264020 333276 264026 333288
rect 264514 333276 264520 333288
rect 264572 333276 264578 333328
rect 265250 333276 265256 333328
rect 265308 333316 265314 333328
rect 266262 333316 266268 333328
rect 265308 333288 266268 333316
rect 265308 333276 265314 333288
rect 266262 333276 266268 333288
rect 266320 333276 266326 333328
rect 267734 333316 267740 333328
rect 267695 333288 267740 333316
rect 267734 333276 267740 333288
rect 267792 333276 267798 333328
rect 267921 333319 267979 333325
rect 267921 333285 267933 333319
rect 267967 333316 267979 333319
rect 268654 333316 268660 333328
rect 267967 333288 268660 333316
rect 267967 333285 267979 333288
rect 267921 333279 267979 333285
rect 268654 333276 268660 333288
rect 268712 333276 268718 333328
rect 271785 333319 271843 333325
rect 271785 333285 271797 333319
rect 271831 333316 271843 333319
rect 433334 333316 433340 333328
rect 271831 333288 433340 333316
rect 271831 333285 271843 333288
rect 271785 333279 271843 333285
rect 433334 333276 433340 333288
rect 433392 333276 433398 333328
rect 28994 333208 29000 333260
rect 29052 333248 29058 333260
rect 237282 333248 237288 333260
rect 29052 333220 237288 333248
rect 29052 333208 29058 333220
rect 237282 333208 237288 333220
rect 237340 333208 237346 333260
rect 238202 333208 238208 333260
rect 238260 333248 238266 333260
rect 238665 333251 238723 333257
rect 238665 333248 238677 333251
rect 238260 333220 238677 333248
rect 238260 333208 238266 333220
rect 238665 333217 238677 333220
rect 238711 333217 238723 333251
rect 238665 333211 238723 333217
rect 239030 333208 239036 333260
rect 239088 333248 239094 333260
rect 239950 333248 239956 333260
rect 239088 333220 239956 333248
rect 239088 333208 239094 333220
rect 239950 333208 239956 333220
rect 240008 333208 240014 333260
rect 240965 333251 241023 333257
rect 240965 333217 240977 333251
rect 241011 333248 241023 333251
rect 241238 333248 241244 333260
rect 241011 333220 241244 333248
rect 241011 333217 241023 333220
rect 240965 333211 241023 333217
rect 241238 333208 241244 333220
rect 241296 333208 241302 333260
rect 242158 333208 242164 333260
rect 242216 333248 242222 333260
rect 243538 333248 243544 333260
rect 242216 333220 243544 333248
rect 242216 333208 242222 333220
rect 243538 333208 243544 333220
rect 243596 333208 243602 333260
rect 245841 333251 245899 333257
rect 245841 333217 245853 333251
rect 245887 333248 245899 333251
rect 246574 333248 246580 333260
rect 245887 333220 246580 333248
rect 245887 333217 245899 333220
rect 245841 333211 245899 333217
rect 246574 333208 246580 333220
rect 246632 333208 246638 333260
rect 257246 333208 257252 333260
rect 257304 333248 257310 333260
rect 436738 333248 436744 333260
rect 257304 333220 436744 333248
rect 257304 333208 257310 333220
rect 436738 333208 436744 333220
rect 436796 333208 436802 333260
rect 148962 333140 148968 333192
rect 149020 333180 149026 333192
rect 247310 333180 247316 333192
rect 149020 333152 247316 333180
rect 149020 333140 149026 333152
rect 247310 333140 247316 333152
rect 247368 333140 247374 333192
rect 247402 333140 247408 333192
rect 247460 333180 247466 333192
rect 248049 333183 248107 333189
rect 248049 333180 248061 333183
rect 247460 333152 248061 333180
rect 247460 333140 247466 333152
rect 248049 333149 248061 333152
rect 248095 333149 248107 333183
rect 248049 333143 248107 333149
rect 250162 333140 250168 333192
rect 250220 333180 250226 333192
rect 250533 333183 250591 333189
rect 250533 333180 250545 333183
rect 250220 333152 250545 333180
rect 250220 333140 250226 333152
rect 250533 333149 250545 333152
rect 250579 333149 250591 333183
rect 250533 333143 250591 333149
rect 251729 333183 251787 333189
rect 251729 333149 251741 333183
rect 251775 333180 251787 333183
rect 252370 333180 252376 333192
rect 251775 333152 252376 333180
rect 251775 333149 251787 333152
rect 251729 333143 251787 333149
rect 252370 333140 252376 333152
rect 252428 333140 252434 333192
rect 263873 333183 263931 333189
rect 263873 333149 263885 333183
rect 263919 333180 263931 333183
rect 271417 333183 271475 333189
rect 271417 333180 271429 333183
rect 263919 333152 271429 333180
rect 263919 333149 263931 333152
rect 263873 333143 263931 333149
rect 271417 333149 271429 333152
rect 271463 333149 271475 333183
rect 271417 333143 271475 333149
rect 271506 333140 271512 333192
rect 271564 333180 271570 333192
rect 271690 333180 271696 333192
rect 271564 333152 271696 333180
rect 271564 333140 271570 333152
rect 271690 333140 271696 333152
rect 271748 333140 271754 333192
rect 390646 333180 390652 333192
rect 271800 333152 390652 333180
rect 153102 333072 153108 333124
rect 153160 333112 153166 333124
rect 247954 333112 247960 333124
rect 153160 333084 247960 333112
rect 153160 333072 153166 333084
rect 247954 333072 247960 333084
rect 248012 333072 248018 333124
rect 268102 333072 268108 333124
rect 268160 333112 268166 333124
rect 271800 333112 271828 333152
rect 390646 333140 390652 333152
rect 390704 333140 390710 333192
rect 380894 333112 380900 333124
rect 268160 333084 271828 333112
rect 271892 333084 380900 333112
rect 268160 333072 268166 333084
rect 151722 333004 151728 333056
rect 151780 333044 151786 333056
rect 247589 333047 247647 333053
rect 247589 333044 247601 333047
rect 151780 333016 247601 333044
rect 151780 333004 151786 333016
rect 247589 333013 247601 333016
rect 247635 333013 247647 333047
rect 247589 333007 247647 333013
rect 267093 333047 267151 333053
rect 267093 333013 267105 333047
rect 267139 333044 267151 333047
rect 271892 333044 271920 333084
rect 380894 333072 380900 333084
rect 380952 333072 380958 333124
rect 362954 333044 362960 333056
rect 267139 333016 271920 333044
rect 271984 333016 362960 333044
rect 267139 333013 267151 333016
rect 267093 333007 267151 333013
rect 154482 332936 154488 332988
rect 154540 332976 154546 332988
rect 245378 332976 245384 332988
rect 154540 332948 245384 332976
rect 154540 332936 154546 332948
rect 245378 332936 245384 332948
rect 245436 332936 245442 332988
rect 265710 332936 265716 332988
rect 265768 332976 265774 332988
rect 271984 332976 272012 333016
rect 362954 333004 362960 333016
rect 363012 333004 363018 333056
rect 358814 332976 358820 332988
rect 265768 332948 272012 332976
rect 272076 332948 358820 332976
rect 265768 332936 265774 332948
rect 180702 332868 180708 332920
rect 180760 332908 180766 332920
rect 250254 332908 250260 332920
rect 180760 332880 250260 332908
rect 180760 332868 180766 332880
rect 250254 332868 250260 332880
rect 250312 332868 250318 332920
rect 265342 332868 265348 332920
rect 265400 332908 265406 332920
rect 272076 332908 272104 332948
rect 358814 332936 358820 332948
rect 358872 332936 358878 332988
rect 265400 332880 272104 332908
rect 272153 332911 272211 332917
rect 265400 332868 265406 332880
rect 272153 332877 272165 332911
rect 272199 332908 272211 332911
rect 340966 332908 340972 332920
rect 272199 332880 340972 332908
rect 272199 332877 272211 332880
rect 272153 332871 272211 332877
rect 340966 332868 340972 332880
rect 341024 332868 341030 332920
rect 209682 332800 209688 332852
rect 209740 332840 209746 332852
rect 252189 332843 252247 332849
rect 252189 332840 252201 332843
rect 209740 332812 252201 332840
rect 209740 332800 209746 332812
rect 252189 332809 252201 332812
rect 252235 332809 252247 332843
rect 252189 332803 252247 332809
rect 265066 332800 265072 332852
rect 265124 332840 265130 332852
rect 356054 332840 356060 332852
rect 265124 332812 356060 332840
rect 265124 332800 265130 332812
rect 356054 332800 356060 332812
rect 356112 332800 356118 332852
rect 227622 332732 227628 332784
rect 227680 332772 227686 332784
rect 253477 332775 253535 332781
rect 253477 332772 253489 332775
rect 227680 332744 253489 332772
rect 227680 332732 227686 332744
rect 253477 332741 253489 332744
rect 253523 332741 253535 332775
rect 253477 332735 253535 332741
rect 261849 332775 261907 332781
rect 261849 332741 261861 332775
rect 261895 332772 261907 332775
rect 316126 332772 316132 332784
rect 261895 332744 316132 332772
rect 261895 332741 261907 332744
rect 261849 332735 261907 332741
rect 316126 332732 316132 332744
rect 316184 332732 316190 332784
rect 230382 332664 230388 332716
rect 230440 332704 230446 332716
rect 254302 332704 254308 332716
rect 230440 332676 254308 332704
rect 230440 332664 230446 332676
rect 254302 332664 254308 332676
rect 254360 332664 254366 332716
rect 261662 332664 261668 332716
rect 261720 332704 261726 332716
rect 313274 332704 313280 332716
rect 261720 332676 313280 332704
rect 261720 332664 261726 332676
rect 313274 332664 313280 332676
rect 313332 332664 313338 332716
rect 233142 332596 233148 332648
rect 233200 332636 233206 332648
rect 251174 332636 251180 332648
rect 233200 332608 251180 332636
rect 233200 332596 233206 332608
rect 251174 332596 251180 332608
rect 251232 332596 251238 332648
rect 252094 332596 252100 332648
rect 252152 332636 252158 332648
rect 255774 332636 255780 332648
rect 252152 332608 255780 332636
rect 252152 332596 252158 332608
rect 255774 332596 255780 332608
rect 255832 332596 255838 332648
rect 263686 332596 263692 332648
rect 263744 332636 263750 332648
rect 306374 332636 306380 332648
rect 263744 332608 306380 332636
rect 263744 332596 263750 332608
rect 306374 332596 306380 332608
rect 306432 332596 306438 332648
rect 261018 332528 261024 332580
rect 261076 332568 261082 332580
rect 307754 332568 307760 332580
rect 261076 332540 307760 332568
rect 261076 332528 261082 332540
rect 307754 332528 307760 332540
rect 307812 332528 307818 332580
rect 263594 332460 263600 332512
rect 263652 332500 263658 332512
rect 311894 332500 311900 332512
rect 263652 332472 311900 332500
rect 263652 332460 263658 332472
rect 311894 332460 311900 332472
rect 311952 332460 311958 332512
rect 177850 332392 177856 332444
rect 177908 332432 177914 332444
rect 249889 332435 249947 332441
rect 249889 332432 249901 332435
rect 177908 332404 249901 332432
rect 177908 332392 177914 332404
rect 249889 332401 249901 332404
rect 249935 332401 249947 332435
rect 249889 332395 249947 332401
rect 263321 332435 263379 332441
rect 263321 332401 263333 332435
rect 263367 332432 263379 332435
rect 318794 332432 318800 332444
rect 263367 332404 318800 332432
rect 263367 332401 263379 332404
rect 263321 332395 263379 332401
rect 318794 332392 318800 332404
rect 318852 332392 318858 332444
rect 161382 332324 161388 332376
rect 161440 332364 161446 332376
rect 248414 332364 248420 332376
rect 161440 332336 248420 332364
rect 161440 332324 161446 332336
rect 248414 332324 248420 332336
rect 248472 332324 248478 332376
rect 262861 332367 262919 332373
rect 262861 332333 262873 332367
rect 262907 332364 262919 332367
rect 329834 332364 329840 332376
rect 262907 332336 329840 332364
rect 262907 332333 262919 332336
rect 262861 332327 262919 332333
rect 329834 332324 329840 332336
rect 329892 332324 329898 332376
rect 140682 332256 140688 332308
rect 140740 332296 140746 332308
rect 246758 332296 246764 332308
rect 140740 332268 246764 332296
rect 140740 332256 140746 332268
rect 246758 332256 246764 332268
rect 246816 332256 246822 332308
rect 270865 332299 270923 332305
rect 270865 332265 270877 332299
rect 270911 332296 270923 332299
rect 280065 332299 280123 332305
rect 280065 332296 280077 332299
rect 270911 332268 280077 332296
rect 270911 332265 270923 332268
rect 270865 332259 270923 332265
rect 280065 332265 280077 332268
rect 280111 332265 280123 332299
rect 280065 332259 280123 332265
rect 280154 332256 280160 332308
rect 280212 332296 280218 332308
rect 280338 332296 280344 332308
rect 280212 332268 280344 332296
rect 280212 332256 280218 332268
rect 280338 332256 280344 332268
rect 280396 332256 280402 332308
rect 280433 332299 280491 332305
rect 280433 332265 280445 332299
rect 280479 332296 280491 332299
rect 357434 332296 357440 332308
rect 280479 332268 357440 332296
rect 280479 332265 280491 332268
rect 280433 332259 280491 332265
rect 357434 332256 357440 332268
rect 357492 332256 357498 332308
rect 126882 332188 126888 332240
rect 126940 332228 126946 332240
rect 245565 332231 245623 332237
rect 245565 332228 245577 332231
rect 126940 332200 245577 332228
rect 126940 332188 126946 332200
rect 245565 332197 245577 332200
rect 245611 332197 245623 332231
rect 245565 332191 245623 332197
rect 275278 332188 275284 332240
rect 275336 332228 275342 332240
rect 423766 332228 423772 332240
rect 275336 332200 423772 332228
rect 275336 332188 275342 332200
rect 423766 332188 423772 332200
rect 423824 332188 423830 332240
rect 97902 332120 97908 332172
rect 97960 332160 97966 332172
rect 243446 332160 243452 332172
rect 97960 332132 243452 332160
rect 97960 332120 97966 332132
rect 243446 332120 243452 332132
rect 243504 332120 243510 332172
rect 259546 332120 259552 332172
rect 259604 332160 259610 332172
rect 437014 332160 437020 332172
rect 259604 332132 437020 332160
rect 259604 332120 259610 332132
rect 437014 332120 437020 332132
rect 437072 332120 437078 332172
rect 85482 332052 85488 332104
rect 85540 332092 85546 332104
rect 240778 332092 240784 332104
rect 85540 332064 240784 332092
rect 85540 332052 85546 332064
rect 240778 332052 240784 332064
rect 240836 332052 240842 332104
rect 258810 332052 258816 332104
rect 258868 332092 258874 332104
rect 436922 332092 436928 332104
rect 258868 332064 436928 332092
rect 258868 332052 258874 332064
rect 436922 332052 436928 332064
rect 436980 332052 436986 332104
rect 81342 331984 81348 332036
rect 81400 332024 81406 332036
rect 241882 332024 241888 332036
rect 81400 331996 241888 332024
rect 81400 331984 81406 331996
rect 241882 331984 241888 331996
rect 241940 331984 241946 332036
rect 255130 331984 255136 332036
rect 255188 332024 255194 332036
rect 436830 332024 436836 332036
rect 255188 331996 436836 332024
rect 255188 331984 255194 331996
rect 436830 331984 436836 331996
rect 436888 331984 436894 332036
rect 59262 331916 59268 331968
rect 59320 331956 59326 331968
rect 239858 331956 239864 331968
rect 59320 331928 239864 331956
rect 59320 331916 59326 331928
rect 239858 331916 239864 331928
rect 239916 331916 239922 331968
rect 240778 331916 240784 331968
rect 240836 331956 240842 331968
rect 240873 331959 240931 331965
rect 240873 331956 240885 331959
rect 240836 331928 240885 331956
rect 240836 331916 240842 331928
rect 240873 331925 240885 331928
rect 240919 331925 240931 331959
rect 240873 331919 240931 331925
rect 252554 331916 252560 331968
rect 252612 331956 252618 331968
rect 519538 331956 519544 331968
rect 252612 331928 519544 331956
rect 252612 331916 252618 331928
rect 519538 331916 519544 331928
rect 519596 331916 519602 331968
rect 19242 331848 19248 331900
rect 19300 331888 19306 331900
rect 236454 331888 236460 331900
rect 19300 331860 236460 331888
rect 19300 331848 19306 331860
rect 236454 331848 236460 331860
rect 236512 331848 236518 331900
rect 259270 331848 259276 331900
rect 259328 331888 259334 331900
rect 285674 331888 285680 331900
rect 259328 331860 285680 331888
rect 259328 331848 259334 331860
rect 285674 331848 285680 331860
rect 285732 331848 285738 331900
rect 285766 331848 285772 331900
rect 285824 331888 285830 331900
rect 580994 331888 581000 331900
rect 285824 331860 581000 331888
rect 285824 331848 285830 331860
rect 580994 331848 581000 331860
rect 581052 331848 581058 331900
rect 262398 331780 262404 331832
rect 262456 331820 262462 331832
rect 300854 331820 300860 331832
rect 262456 331792 300860 331820
rect 262456 331780 262462 331792
rect 300854 331780 300860 331792
rect 300912 331780 300918 331832
rect 266446 331712 266452 331764
rect 266504 331752 266510 331764
rect 298094 331752 298100 331764
rect 266504 331724 298100 331752
rect 266504 331712 266510 331724
rect 298094 331712 298100 331724
rect 298152 331712 298158 331764
rect 248966 331644 248972 331696
rect 249024 331684 249030 331696
rect 249242 331684 249248 331696
rect 249024 331656 249248 331684
rect 249024 331644 249030 331656
rect 249242 331644 249248 331656
rect 249300 331644 249306 331696
rect 259638 331644 259644 331696
rect 259696 331684 259702 331696
rect 284849 331687 284907 331693
rect 284849 331684 284861 331687
rect 259696 331656 284861 331684
rect 259696 331644 259702 331656
rect 284849 331653 284861 331656
rect 284895 331653 284907 331687
rect 284849 331647 284907 331653
rect 284938 331644 284944 331696
rect 284996 331684 285002 331696
rect 292298 331684 292304 331696
rect 284996 331656 292304 331684
rect 284996 331644 285002 331656
rect 292298 331644 292304 331656
rect 292356 331644 292362 331696
rect 248874 331576 248880 331628
rect 248932 331616 248938 331628
rect 249334 331616 249340 331628
rect 248932 331588 249340 331616
rect 248932 331576 248938 331588
rect 249334 331576 249340 331588
rect 249392 331576 249398 331628
rect 276474 331576 276480 331628
rect 276532 331616 276538 331628
rect 289538 331616 289544 331628
rect 276532 331588 289544 331616
rect 276532 331576 276538 331588
rect 289538 331576 289544 331588
rect 289596 331576 289602 331628
rect 274266 331508 274272 331560
rect 274324 331548 274330 331560
rect 290642 331548 290648 331560
rect 274324 331520 290648 331548
rect 274324 331508 274330 331520
rect 290642 331508 290648 331520
rect 290700 331508 290706 331560
rect 275370 331440 275376 331492
rect 275428 331480 275434 331492
rect 290918 331480 290924 331492
rect 275428 331452 290924 331480
rect 275428 331440 275434 331452
rect 290918 331440 290924 331452
rect 290976 331440 290982 331492
rect 273254 331372 273260 331424
rect 273312 331412 273318 331424
rect 289446 331412 289452 331424
rect 273312 331384 289452 331412
rect 273312 331372 273318 331384
rect 289446 331372 289452 331384
rect 289504 331372 289510 331424
rect 274818 331304 274824 331356
rect 274876 331344 274882 331356
rect 290734 331344 290740 331356
rect 274876 331316 290740 331344
rect 274876 331304 274882 331316
rect 290734 331304 290740 331316
rect 290792 331304 290798 331356
rect 40034 331236 40040 331288
rect 40092 331276 40098 331288
rect 238294 331276 238300 331288
rect 40092 331248 238300 331276
rect 40092 331236 40098 331248
rect 238294 331236 238300 331248
rect 238352 331236 238358 331288
rect 280246 331236 280252 331288
rect 280304 331276 280310 331288
rect 280982 331276 280988 331288
rect 280304 331248 280988 331276
rect 280304 331236 280310 331248
rect 280982 331236 280988 331248
rect 281040 331236 281046 331288
rect 284849 331279 284907 331285
rect 284849 331245 284861 331279
rect 284895 331276 284907 331279
rect 291194 331276 291200 331288
rect 284895 331248 291200 331276
rect 284895 331245 284907 331248
rect 284849 331239 284907 331245
rect 291194 331236 291200 331248
rect 291252 331236 291258 331288
rect 279804 330840 282914 330868
rect 272150 330692 272156 330744
rect 272208 330732 272214 330744
rect 272208 330704 277394 330732
rect 272208 330692 272214 330704
rect 273806 330624 273812 330676
rect 273864 330624 273870 330676
rect 275370 330624 275376 330676
rect 275428 330664 275434 330676
rect 275646 330664 275652 330676
rect 275428 330636 275652 330664
rect 275428 330624 275434 330636
rect 275646 330624 275652 330636
rect 275704 330624 275710 330676
rect 277366 330664 277394 330704
rect 277854 330692 277860 330744
rect 277912 330732 277918 330744
rect 278038 330732 278044 330744
rect 277912 330704 278044 330732
rect 277912 330692 277918 330704
rect 278038 330692 278044 330704
rect 278096 330692 278102 330744
rect 279050 330692 279056 330744
rect 279108 330732 279114 330744
rect 279694 330732 279700 330744
rect 279108 330704 279700 330732
rect 279108 330692 279114 330704
rect 279694 330692 279700 330704
rect 279752 330692 279758 330744
rect 279804 330664 279832 330840
rect 277366 330636 279832 330664
rect 282886 330664 282914 330840
rect 422938 330664 422944 330676
rect 282886 330636 422944 330664
rect 422938 330624 422944 330636
rect 422996 330624 423002 330676
rect 23382 330488 23388 330540
rect 23440 330528 23446 330540
rect 236822 330528 236828 330540
rect 23440 330500 236828 330528
rect 23440 330488 23446 330500
rect 236822 330488 236828 330500
rect 236880 330488 236886 330540
rect 273714 330284 273720 330336
rect 273772 330324 273778 330336
rect 273824 330324 273852 330624
rect 277762 330556 277768 330608
rect 277820 330596 277826 330608
rect 278038 330596 278044 330608
rect 277820 330568 278044 330596
rect 277820 330556 277826 330568
rect 278038 330556 278044 330568
rect 278096 330556 278102 330608
rect 280982 330556 280988 330608
rect 281040 330596 281046 330608
rect 281169 330599 281227 330605
rect 281169 330596 281181 330599
rect 281040 330568 281181 330596
rect 281040 330556 281046 330568
rect 281169 330565 281181 330568
rect 281215 330565 281227 330599
rect 281169 330559 281227 330565
rect 285582 330556 285588 330608
rect 285640 330596 285646 330608
rect 538214 330596 538220 330608
rect 285640 330568 538220 330596
rect 285640 330556 285646 330568
rect 538214 330556 538220 330568
rect 538272 330556 538278 330608
rect 275646 330488 275652 330540
rect 275704 330528 275710 330540
rect 275830 330528 275836 330540
rect 275704 330500 275836 330528
rect 275704 330488 275710 330500
rect 275830 330488 275836 330500
rect 275888 330488 275894 330540
rect 281813 330531 281871 330537
rect 281813 330497 281825 330531
rect 281859 330528 281871 330531
rect 282362 330528 282368 330540
rect 281859 330500 282368 330528
rect 281859 330497 281871 330500
rect 281813 330491 281871 330497
rect 282362 330488 282368 330500
rect 282420 330488 282426 330540
rect 282914 330488 282920 330540
rect 282972 330528 282978 330540
rect 574094 330528 574100 330540
rect 282972 330500 574100 330528
rect 282972 330488 282978 330500
rect 574094 330488 574100 330500
rect 574152 330488 574158 330540
rect 278958 330420 278964 330472
rect 279016 330460 279022 330472
rect 279878 330460 279884 330472
rect 279016 330432 279884 330460
rect 279016 330420 279022 330432
rect 279878 330420 279884 330432
rect 279936 330420 279942 330472
rect 280338 330420 280344 330472
rect 280396 330460 280402 330472
rect 280890 330460 280896 330472
rect 280396 330432 280896 330460
rect 280396 330420 280402 330432
rect 280890 330420 280896 330432
rect 280948 330420 280954 330472
rect 281534 330420 281540 330472
rect 281592 330460 281598 330472
rect 282270 330460 282276 330472
rect 281592 330432 282276 330460
rect 281592 330420 281598 330432
rect 282270 330420 282276 330432
rect 282328 330420 282334 330472
rect 273772 330296 273852 330324
rect 273772 330284 273778 330296
rect 272245 330259 272303 330265
rect 272245 330225 272257 330259
rect 272291 330256 272303 330259
rect 273898 330256 273904 330268
rect 272291 330228 273904 330256
rect 272291 330225 272303 330228
rect 272245 330219 272303 330225
rect 273898 330216 273904 330228
rect 273956 330216 273962 330268
rect 272613 330191 272671 330197
rect 272613 330157 272625 330191
rect 272659 330188 272671 330191
rect 274082 330188 274088 330200
rect 272659 330160 274088 330188
rect 272659 330157 272671 330160
rect 272613 330151 272671 330157
rect 274082 330148 274088 330160
rect 274140 330148 274146 330200
rect 266998 329060 267004 329112
rect 267056 329100 267062 329112
rect 267274 329100 267280 329112
rect 267056 329072 267280 329100
rect 267056 329060 267062 329072
rect 267274 329060 267280 329072
rect 267332 329060 267338 329112
rect 238294 327700 238300 327752
rect 238352 327740 238358 327752
rect 437106 327740 437112 327752
rect 238352 327712 437112 327740
rect 238352 327700 238358 327712
rect 437106 327700 437112 327712
rect 437164 327700 437170 327752
rect 265158 327632 265164 327684
rect 265216 327672 265222 327684
rect 265526 327672 265532 327684
rect 265216 327644 265532 327672
rect 265216 327632 265222 327644
rect 265526 327632 265532 327644
rect 265584 327632 265590 327684
rect 244642 326748 244648 326800
rect 244700 326788 244706 326800
rect 244826 326788 244832 326800
rect 244700 326760 244832 326788
rect 244700 326748 244706 326760
rect 244826 326748 244832 326760
rect 244884 326748 244890 326800
rect 244734 326680 244740 326732
rect 244792 326680 244798 326732
rect 245838 326680 245844 326732
rect 245896 326720 245902 326732
rect 246022 326720 246028 326732
rect 245896 326692 246028 326720
rect 245896 326680 245902 326692
rect 246022 326680 246028 326692
rect 246080 326680 246086 326732
rect 241606 326476 241612 326528
rect 241664 326516 241670 326528
rect 242710 326516 242716 326528
rect 241664 326488 242716 326516
rect 241664 326476 241670 326488
rect 242710 326476 242716 326488
rect 242768 326476 242774 326528
rect 244752 326516 244780 326680
rect 248690 326544 248696 326596
rect 248748 326584 248754 326596
rect 249150 326584 249156 326596
rect 248748 326556 249156 326584
rect 248748 326544 248754 326556
rect 249150 326544 249156 326556
rect 249208 326544 249214 326596
rect 255406 326544 255412 326596
rect 255464 326584 255470 326596
rect 256418 326584 256424 326596
rect 255464 326556 256424 326584
rect 255464 326544 255470 326556
rect 256418 326544 256424 326556
rect 256476 326544 256482 326596
rect 270954 326544 270960 326596
rect 271012 326584 271018 326596
rect 271322 326584 271328 326596
rect 271012 326556 271328 326584
rect 271012 326544 271018 326556
rect 271322 326544 271328 326556
rect 271380 326544 271386 326596
rect 244826 326516 244832 326528
rect 244752 326488 244832 326516
rect 244826 326476 244832 326488
rect 244884 326476 244890 326528
rect 255498 326476 255504 326528
rect 255556 326516 255562 326528
rect 255774 326516 255780 326528
rect 255556 326488 255780 326516
rect 255556 326476 255562 326488
rect 255774 326476 255780 326488
rect 255832 326476 255838 326528
rect 255958 326476 255964 326528
rect 256016 326516 256022 326528
rect 256142 326516 256148 326528
rect 256016 326488 256148 326516
rect 256016 326476 256022 326488
rect 256142 326476 256148 326488
rect 256200 326476 256206 326528
rect 257430 326476 257436 326528
rect 257488 326516 257494 326528
rect 257798 326516 257804 326528
rect 257488 326488 257804 326516
rect 257488 326476 257494 326488
rect 257798 326476 257804 326488
rect 257856 326476 257862 326528
rect 270494 326476 270500 326528
rect 270552 326516 270558 326528
rect 271414 326516 271420 326528
rect 270552 326488 271420 326516
rect 270552 326476 270558 326488
rect 271414 326476 271420 326488
rect 271472 326476 271478 326528
rect 235626 326408 235632 326460
rect 235684 326448 235690 326460
rect 240686 326448 240692 326460
rect 235684 326420 235764 326448
rect 240647 326420 240692 326448
rect 235684 326408 235690 326420
rect 235736 326256 235764 326420
rect 240686 326408 240692 326420
rect 240744 326408 240750 326460
rect 241790 326408 241796 326460
rect 241848 326448 241854 326460
rect 242618 326448 242624 326460
rect 241848 326420 242624 326448
rect 241848 326408 241854 326420
rect 242618 326408 242624 326420
rect 242676 326408 242682 326460
rect 243078 326408 243084 326460
rect 243136 326448 243142 326460
rect 243906 326448 243912 326460
rect 243136 326420 243912 326448
rect 243136 326408 243142 326420
rect 243906 326408 243912 326420
rect 243964 326408 243970 326460
rect 244550 326408 244556 326460
rect 244608 326448 244614 326460
rect 245010 326448 245016 326460
rect 244608 326420 245016 326448
rect 244608 326408 244614 326420
rect 245010 326408 245016 326420
rect 245068 326408 245074 326460
rect 246114 326408 246120 326460
rect 246172 326448 246178 326460
rect 246390 326448 246396 326460
rect 246172 326420 246396 326448
rect 246172 326408 246178 326420
rect 246390 326408 246396 326420
rect 246448 326408 246454 326460
rect 247310 326408 247316 326460
rect 247368 326448 247374 326460
rect 248138 326448 248144 326460
rect 247368 326420 248144 326448
rect 247368 326408 247374 326420
rect 248138 326408 248144 326420
rect 248196 326408 248202 326460
rect 250254 326408 250260 326460
rect 250312 326448 250318 326460
rect 250806 326448 250812 326460
rect 250312 326420 250812 326448
rect 250312 326408 250318 326420
rect 250806 326408 250812 326420
rect 250864 326408 250870 326460
rect 252738 326408 252744 326460
rect 252796 326448 252802 326460
rect 253290 326448 253296 326460
rect 252796 326420 253296 326448
rect 252796 326408 252802 326420
rect 253290 326408 253296 326420
rect 253348 326408 253354 326460
rect 269758 326408 269764 326460
rect 269816 326448 269822 326460
rect 269942 326448 269948 326460
rect 269816 326420 269948 326448
rect 269816 326408 269822 326420
rect 269942 326408 269948 326420
rect 270000 326408 270006 326460
rect 270954 326408 270960 326460
rect 271012 326448 271018 326460
rect 271138 326448 271144 326460
rect 271012 326420 271144 326448
rect 271012 326408 271018 326420
rect 271138 326408 271144 326420
rect 271196 326408 271202 326460
rect 236454 326340 236460 326392
rect 236512 326380 236518 326392
rect 236914 326380 236920 326392
rect 236512 326352 236920 326380
rect 236512 326340 236518 326352
rect 236914 326340 236920 326352
rect 236972 326340 236978 326392
rect 237650 326340 237656 326392
rect 237708 326380 237714 326392
rect 238110 326380 238116 326392
rect 237708 326352 238116 326380
rect 237708 326340 237714 326352
rect 238110 326340 238116 326352
rect 238168 326340 238174 326392
rect 240410 326340 240416 326392
rect 240468 326380 240474 326392
rect 240870 326380 240876 326392
rect 240468 326352 240876 326380
rect 240468 326340 240474 326352
rect 240870 326340 240876 326352
rect 240928 326340 240934 326392
rect 241882 326340 241888 326392
rect 241940 326380 241946 326392
rect 242250 326380 242256 326392
rect 241940 326352 242256 326380
rect 241940 326340 241946 326352
rect 242250 326340 242256 326352
rect 242308 326340 242314 326392
rect 243354 326340 243360 326392
rect 243412 326380 243418 326392
rect 243998 326380 244004 326392
rect 243412 326352 244004 326380
rect 243412 326340 243418 326352
rect 243998 326340 244004 326352
rect 244056 326340 244062 326392
rect 247494 326340 247500 326392
rect 247552 326380 247558 326392
rect 248322 326380 248328 326392
rect 247552 326352 248328 326380
rect 247552 326340 247558 326352
rect 248322 326340 248328 326352
rect 248380 326340 248386 326392
rect 248690 326340 248696 326392
rect 248748 326380 248754 326392
rect 249702 326380 249708 326392
rect 248748 326352 249708 326380
rect 248748 326340 248754 326352
rect 249702 326340 249708 326352
rect 249760 326340 249766 326392
rect 250346 326340 250352 326392
rect 250404 326380 250410 326392
rect 250622 326380 250628 326392
rect 250404 326352 250628 326380
rect 250404 326340 250410 326352
rect 250622 326340 250628 326352
rect 250680 326340 250686 326392
rect 251542 326340 251548 326392
rect 251600 326380 251606 326392
rect 252462 326380 252468 326392
rect 251600 326352 252468 326380
rect 251600 326340 251606 326352
rect 252462 326340 252468 326352
rect 252520 326340 252526 326392
rect 252830 326340 252836 326392
rect 252888 326380 252894 326392
rect 253014 326380 253020 326392
rect 252888 326352 253020 326380
rect 252888 326340 252894 326352
rect 253014 326340 253020 326352
rect 253072 326340 253078 326392
rect 254118 326340 254124 326392
rect 254176 326380 254182 326392
rect 254762 326380 254768 326392
rect 254176 326352 254768 326380
rect 254176 326340 254182 326352
rect 254762 326340 254768 326352
rect 254820 326340 254826 326392
rect 258534 326340 258540 326392
rect 258592 326380 258598 326392
rect 258902 326380 258908 326392
rect 258592 326352 258908 326380
rect 258592 326340 258598 326352
rect 258902 326340 258908 326352
rect 258960 326340 258966 326392
rect 260282 326340 260288 326392
rect 260340 326380 260346 326392
rect 260558 326380 260564 326392
rect 260340 326352 260564 326380
rect 260340 326340 260346 326352
rect 260558 326340 260564 326352
rect 260616 326340 260622 326392
rect 263870 326340 263876 326392
rect 263928 326380 263934 326392
rect 264238 326380 264244 326392
rect 263928 326352 264244 326380
rect 263928 326340 263934 326352
rect 264238 326340 264244 326352
rect 264296 326340 264302 326392
rect 271414 326340 271420 326392
rect 271472 326380 271478 326392
rect 271598 326380 271604 326392
rect 271472 326352 271604 326380
rect 271472 326340 271478 326352
rect 271598 326340 271604 326352
rect 271656 326340 271662 326392
rect 283466 326340 283472 326392
rect 283524 326380 283530 326392
rect 283834 326380 283840 326392
rect 283524 326352 283840 326380
rect 283524 326340 283530 326352
rect 283834 326340 283840 326352
rect 283892 326340 283898 326392
rect 241698 326272 241704 326324
rect 241756 326312 241762 326324
rect 242802 326312 242808 326324
rect 241756 326284 242808 326312
rect 241756 326272 241762 326284
rect 242802 326272 242808 326284
rect 242860 326272 242866 326324
rect 243078 326272 243084 326324
rect 243136 326312 243142 326324
rect 244182 326312 244188 326324
rect 243136 326284 244188 326312
rect 243136 326272 243142 326284
rect 244182 326272 244188 326284
rect 244240 326272 244246 326324
rect 235718 326204 235724 326256
rect 235776 326204 235782 326256
rect 240410 326204 240416 326256
rect 240468 326244 240474 326256
rect 241146 326244 241152 326256
rect 240468 326216 241152 326244
rect 240468 326204 240474 326216
rect 241146 326204 241152 326216
rect 241204 326204 241210 326256
rect 244458 326204 244464 326256
rect 244516 326244 244522 326256
rect 244734 326244 244740 326256
rect 244516 326216 244740 326244
rect 244516 326204 244522 326216
rect 244734 326204 244740 326216
rect 244792 326204 244798 326256
rect 246022 326204 246028 326256
rect 246080 326244 246086 326256
rect 246942 326244 246948 326256
rect 246080 326216 246948 326244
rect 246080 326204 246086 326216
rect 246942 326204 246948 326216
rect 247000 326204 247006 326256
rect 248874 326204 248880 326256
rect 248932 326244 248938 326256
rect 249058 326244 249064 326256
rect 248932 326216 249064 326244
rect 248932 326204 248938 326216
rect 249058 326204 249064 326216
rect 249116 326204 249122 326256
rect 250346 326204 250352 326256
rect 250404 326244 250410 326256
rect 251082 326244 251088 326256
rect 250404 326216 251088 326244
rect 250404 326204 250410 326216
rect 251082 326204 251088 326216
rect 251140 326204 251146 326256
rect 252646 326204 252652 326256
rect 252704 326244 252710 326256
rect 253290 326244 253296 326256
rect 252704 326216 253296 326244
rect 252704 326204 252710 326216
rect 253290 326204 253296 326216
rect 253348 326204 253354 326256
rect 256050 326204 256056 326256
rect 256108 326244 256114 326256
rect 256418 326244 256424 326256
rect 256108 326216 256424 326244
rect 256108 326204 256114 326216
rect 256418 326204 256424 326216
rect 256476 326204 256482 326256
rect 256878 326204 256884 326256
rect 256936 326244 256942 326256
rect 257798 326244 257804 326256
rect 256936 326216 257804 326244
rect 256936 326204 256942 326216
rect 257798 326204 257804 326216
rect 257856 326204 257862 326256
rect 260190 326204 260196 326256
rect 260248 326244 260254 326256
rect 260558 326244 260564 326256
rect 260248 326216 260564 326244
rect 260248 326204 260254 326216
rect 260558 326204 260564 326216
rect 260616 326204 260622 326256
rect 245930 326136 245936 326188
rect 245988 326176 245994 326188
rect 246850 326176 246856 326188
rect 245988 326148 246856 326176
rect 245988 326136 245994 326148
rect 246850 326136 246856 326148
rect 246908 326136 246914 326188
rect 255590 326136 255596 326188
rect 255648 326176 255654 326188
rect 256510 326176 256516 326188
rect 255648 326148 256516 326176
rect 255648 326136 255654 326148
rect 256510 326136 256516 326148
rect 256568 326136 256574 326188
rect 259638 326136 259644 326188
rect 259696 326176 259702 326188
rect 259822 326176 259828 326188
rect 259696 326148 259828 326176
rect 259696 326136 259702 326148
rect 259822 326136 259828 326148
rect 259880 326136 259886 326188
rect 244458 326068 244464 326120
rect 244516 326108 244522 326120
rect 245470 326108 245476 326120
rect 244516 326080 245476 326108
rect 244516 326068 244522 326080
rect 245470 326068 245476 326080
rect 245528 326068 245534 326120
rect 246206 326068 246212 326120
rect 246264 326108 246270 326120
rect 246666 326108 246672 326120
rect 246264 326080 246672 326108
rect 246264 326068 246270 326080
rect 246666 326068 246672 326080
rect 246724 326068 246730 326120
rect 248506 326068 248512 326120
rect 248564 326108 248570 326120
rect 249058 326108 249064 326120
rect 248564 326080 249064 326108
rect 248564 326068 248570 326080
rect 249058 326068 249064 326080
rect 249116 326068 249122 326120
rect 252738 326068 252744 326120
rect 252796 326108 252802 326120
rect 253658 326108 253664 326120
rect 252796 326080 253664 326108
rect 252796 326068 252802 326080
rect 253658 326068 253664 326080
rect 253716 326068 253722 326120
rect 255314 326068 255320 326120
rect 255372 326108 255378 326120
rect 256234 326108 256240 326120
rect 255372 326080 256240 326108
rect 255372 326068 255378 326080
rect 256234 326068 256240 326080
rect 256292 326068 256298 326120
rect 269114 326068 269120 326120
rect 269172 326108 269178 326120
rect 269758 326108 269764 326120
rect 269172 326080 269764 326108
rect 269172 326068 269178 326080
rect 269758 326068 269764 326080
rect 269816 326068 269822 326120
rect 270862 326068 270868 326120
rect 270920 326108 270926 326120
rect 271322 326108 271328 326120
rect 270920 326080 271328 326108
rect 270920 326068 270926 326080
rect 271322 326068 271328 326080
rect 271380 326068 271386 326120
rect 244918 326000 244924 326052
rect 244976 326040 244982 326052
rect 245286 326040 245292 326052
rect 244976 326012 245292 326040
rect 244976 326000 244982 326012
rect 245286 326000 245292 326012
rect 245344 326000 245350 326052
rect 254670 325932 254676 325984
rect 254728 325972 254734 325984
rect 255222 325972 255228 325984
rect 254728 325944 255228 325972
rect 254728 325932 254734 325944
rect 255222 325932 255228 325944
rect 255280 325932 255286 325984
rect 247218 324368 247224 324420
rect 247276 324408 247282 324420
rect 247862 324408 247868 324420
rect 247276 324380 247868 324408
rect 247276 324368 247282 324380
rect 247862 324368 247868 324380
rect 247920 324368 247926 324420
rect 238938 323824 238944 323876
rect 238996 323864 239002 323876
rect 239674 323864 239680 323876
rect 238996 323836 239680 323864
rect 238996 323824 239002 323836
rect 239674 323824 239680 323836
rect 239732 323824 239738 323876
rect 262858 323416 262864 323468
rect 262916 323456 262922 323468
rect 263134 323456 263140 323468
rect 262916 323428 263140 323456
rect 262916 323416 262922 323428
rect 263134 323416 263140 323428
rect 263192 323416 263198 323468
rect 449158 322872 449164 322924
rect 449216 322912 449222 322924
rect 469398 322912 469404 322924
rect 449216 322884 469404 322912
rect 449216 322872 449222 322884
rect 469398 322872 469404 322884
rect 469456 322872 469462 322924
rect 485038 322872 485044 322924
rect 485096 322912 485102 322924
rect 486326 322912 486332 322924
rect 485096 322884 486332 322912
rect 485096 322872 485102 322884
rect 486326 322872 486332 322884
rect 486384 322872 486390 322924
rect 338758 322804 338764 322856
rect 338816 322844 338822 322856
rect 498194 322844 498200 322856
rect 338816 322816 498200 322844
rect 338816 322804 338822 322816
rect 498194 322804 498200 322816
rect 498252 322804 498258 322856
rect 340138 322736 340144 322788
rect 340196 322776 340202 322788
rect 499206 322776 499212 322788
rect 340196 322748 499212 322776
rect 340196 322736 340202 322748
rect 499206 322736 499212 322748
rect 499264 322736 499270 322788
rect 342898 322668 342904 322720
rect 342956 322708 342962 322720
rect 500678 322708 500684 322720
rect 342956 322680 500684 322708
rect 342956 322668 342962 322680
rect 500678 322668 500684 322680
rect 500736 322668 500742 322720
rect 345658 322600 345664 322652
rect 345716 322640 345722 322652
rect 501230 322640 501236 322652
rect 345716 322612 501236 322640
rect 345716 322600 345722 322612
rect 501230 322600 501236 322612
rect 501288 322600 501294 322652
rect 349798 322532 349804 322584
rect 349856 322572 349862 322584
rect 503254 322572 503260 322584
rect 349856 322544 503260 322572
rect 349856 322532 349862 322544
rect 503254 322532 503260 322544
rect 503312 322532 503318 322584
rect 353938 322464 353944 322516
rect 353996 322504 354002 322516
rect 505462 322504 505468 322516
rect 353996 322476 505468 322504
rect 353996 322464 354002 322476
rect 505462 322464 505468 322476
rect 505520 322464 505526 322516
rect 352650 322396 352656 322448
rect 352708 322436 352714 322448
rect 503806 322436 503812 322448
rect 352708 322408 503812 322436
rect 352708 322396 352714 322408
rect 503806 322396 503812 322408
rect 503864 322396 503870 322448
rect 356698 322328 356704 322380
rect 356756 322368 356762 322380
rect 506934 322368 506940 322380
rect 356756 322340 506940 322368
rect 356756 322328 356762 322340
rect 506934 322328 506940 322340
rect 506992 322328 506998 322380
rect 360838 322260 360844 322312
rect 360896 322300 360902 322312
rect 474550 322300 474556 322312
rect 360896 322272 474556 322300
rect 360896 322260 360902 322272
rect 474550 322260 474556 322272
rect 474608 322260 474614 322312
rect 359458 322192 359464 322244
rect 359516 322232 359522 322244
rect 471974 322232 471980 322244
rect 359516 322204 471980 322232
rect 359516 322192 359522 322204
rect 471974 322192 471980 322204
rect 472032 322192 472038 322244
rect 519538 322192 519544 322244
rect 519596 322232 519602 322244
rect 536926 322232 536932 322244
rect 519596 322204 536932 322232
rect 519596 322192 519602 322204
rect 536926 322192 536932 322204
rect 536984 322192 536990 322244
rect 363598 322124 363604 322176
rect 363656 322164 363662 322176
rect 476758 322164 476764 322176
rect 363656 322136 476764 322164
rect 363656 322124 363662 322136
rect 476758 322124 476764 322136
rect 476816 322124 476822 322176
rect 240778 322056 240784 322108
rect 240836 322096 240842 322108
rect 241422 322096 241428 322108
rect 240836 322068 241428 322096
rect 240836 322056 240842 322068
rect 241422 322056 241428 322068
rect 241480 322056 241486 322108
rect 367738 322056 367744 322108
rect 367796 322096 367802 322108
rect 478230 322096 478236 322108
rect 367796 322068 478236 322096
rect 367796 322056 367802 322068
rect 478230 322056 478236 322068
rect 478288 322056 478294 322108
rect 440878 321988 440884 322040
rect 440936 322028 440942 322040
rect 485406 322028 485412 322040
rect 440936 322000 485412 322028
rect 440936 321988 440942 322000
rect 485406 321988 485412 322000
rect 485464 321988 485470 322040
rect 440970 321920 440976 321972
rect 441028 321960 441034 321972
rect 484394 321960 484400 321972
rect 441028 321932 484400 321960
rect 441028 321920 441034 321932
rect 484394 321920 484400 321932
rect 484452 321920 484458 321972
rect 450538 321852 450544 321904
rect 450596 321892 450602 321904
rect 492766 321892 492772 321904
rect 450596 321864 492772 321892
rect 450596 321852 450602 321864
rect 492766 321852 492772 321864
rect 492824 321852 492830 321904
rect 237742 321784 237748 321836
rect 237800 321824 237806 321836
rect 238662 321824 238668 321836
rect 237800 321796 238668 321824
rect 237800 321784 237806 321796
rect 238662 321784 238668 321796
rect 238720 321784 238726 321836
rect 454678 321784 454684 321836
rect 454736 321824 454742 321836
rect 495526 321824 495532 321836
rect 454736 321796 495532 321824
rect 454736 321784 454742 321796
rect 495526 321784 495532 321796
rect 495584 321784 495590 321836
rect 453298 321716 453304 321768
rect 453356 321756 453362 321768
rect 494238 321756 494244 321768
rect 453356 321728 494244 321756
rect 453356 321716 453362 321728
rect 494238 321716 494244 321728
rect 494296 321716 494302 321768
rect 268378 321648 268384 321700
rect 268436 321688 268442 321700
rect 268436 321660 528554 321688
rect 268436 321648 268442 321660
rect 486418 321580 486424 321632
rect 486476 321620 486482 321632
rect 488166 321620 488172 321632
rect 486476 321592 488172 321620
rect 486476 321580 486482 321592
rect 488166 321580 488172 321592
rect 488224 321580 488230 321632
rect 528526 321620 528554 321660
rect 530026 321620 530032 321632
rect 528526 321592 530032 321620
rect 530026 321580 530032 321592
rect 530084 321620 530090 321632
rect 537018 321620 537024 321632
rect 530084 321592 537024 321620
rect 530084 321580 530090 321592
rect 537018 321580 537024 321592
rect 537076 321580 537082 321632
rect 240686 321076 240692 321088
rect 240647 321048 240692 321076
rect 240686 321036 240692 321048
rect 240744 321036 240750 321088
rect 288986 320832 288992 320884
rect 289044 320872 289050 320884
rect 580902 320872 580908 320884
rect 289044 320844 580908 320872
rect 289044 320832 289050 320844
rect 580902 320832 580908 320844
rect 580960 320832 580966 320884
rect 3326 306212 3332 306264
rect 3384 306252 3390 306264
rect 6638 306252 6644 306264
rect 3384 306224 6644 306252
rect 3384 306212 3390 306224
rect 6638 306212 6644 306224
rect 6696 306212 6702 306264
rect 284846 300092 284852 300144
rect 284904 300132 284910 300144
rect 292390 300132 292396 300144
rect 284904 300104 292396 300132
rect 284904 300092 284910 300104
rect 292390 300092 292396 300104
rect 292448 300092 292454 300144
rect 237742 278740 237748 278792
rect 237800 278780 237806 278792
rect 238110 278780 238116 278792
rect 237800 278752 238116 278780
rect 237800 278740 237806 278752
rect 238110 278740 238116 278752
rect 238168 278780 238174 278792
rect 437382 278780 437388 278792
rect 238168 278752 437388 278780
rect 238168 278740 238174 278752
rect 437382 278740 437388 278752
rect 437440 278740 437446 278792
rect 537570 273164 537576 273216
rect 537628 273204 537634 273216
rect 580166 273204 580172 273216
rect 537628 273176 580172 273204
rect 537628 273164 537634 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 436922 271940 436928 271992
rect 436980 271980 436986 271992
rect 437106 271980 437112 271992
rect 436980 271952 437112 271980
rect 436980 271940 436986 271952
rect 437106 271940 437112 271952
rect 437164 271940 437170 271992
rect 249242 271804 249248 271856
rect 249300 271844 249306 271856
rect 436922 271844 436928 271856
rect 249300 271816 436928 271844
rect 249300 271804 249306 271816
rect 436922 271804 436928 271816
rect 436980 271804 436986 271856
rect 436922 269016 436928 269068
rect 436980 269056 436986 269068
rect 437106 269056 437112 269068
rect 436980 269028 437112 269056
rect 436980 269016 436986 269028
rect 437106 269016 437112 269028
rect 437164 269016 437170 269068
rect 436830 266772 436836 266824
rect 436888 266812 436894 266824
rect 437198 266812 437204 266824
rect 436888 266784 437204 266812
rect 436888 266772 436894 266784
rect 437198 266772 437204 266784
rect 437256 266772 437262 266824
rect 537478 259360 537484 259412
rect 537536 259400 537542 259412
rect 579798 259400 579804 259412
rect 537536 259372 579804 259400
rect 537536 259360 537542 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 2774 254600 2780 254652
rect 2832 254640 2838 254652
rect 5350 254640 5356 254652
rect 2832 254612 5356 254640
rect 2832 254600 2838 254612
rect 5350 254600 5356 254612
rect 5408 254600 5414 254652
rect 370498 248344 370504 248396
rect 370556 248384 370562 248396
rect 436094 248384 436100 248396
rect 370556 248356 436100 248384
rect 370556 248344 370562 248356
rect 436094 248344 436100 248356
rect 436152 248344 436158 248396
rect 290826 245556 290832 245608
rect 290884 245596 290890 245608
rect 436094 245596 436100 245608
rect 290884 245568 436100 245596
rect 290884 245556 290890 245568
rect 436094 245556 436100 245568
rect 436152 245556 436158 245608
rect 2774 241340 2780 241392
rect 2832 241380 2838 241392
rect 5258 241380 5264 241392
rect 2832 241352 5264 241380
rect 2832 241340 2838 241352
rect 5258 241340 5264 241352
rect 5316 241340 5322 241392
rect 232774 240728 232780 240780
rect 232832 240768 232838 240780
rect 439406 240768 439412 240780
rect 232832 240740 439412 240768
rect 232832 240728 232838 240740
rect 439406 240728 439412 240740
rect 439464 240728 439470 240780
rect 284018 240048 284024 240100
rect 284076 240088 284082 240100
rect 438578 240088 438584 240100
rect 284076 240060 438584 240088
rect 284076 240048 284082 240060
rect 438578 240048 438584 240060
rect 438636 240048 438642 240100
rect 271966 239980 271972 240032
rect 272024 240020 272030 240032
rect 272024 239992 431954 240020
rect 272024 239980 272030 239992
rect 285306 239912 285312 239964
rect 285364 239952 285370 239964
rect 364334 239952 364340 239964
rect 285364 239924 364340 239952
rect 285364 239912 285370 239924
rect 364334 239912 364340 239924
rect 364392 239912 364398 239964
rect 431926 239884 431954 239992
rect 437290 239980 437296 240032
rect 437348 240020 437354 240032
rect 439866 240020 439872 240032
rect 437348 239992 439872 240020
rect 437348 239980 437354 239992
rect 439866 239980 439872 239992
rect 439924 239980 439930 240032
rect 437106 239912 437112 239964
rect 437164 239952 437170 239964
rect 538490 239952 538496 239964
rect 437164 239924 538496 239952
rect 437164 239912 437170 239924
rect 538490 239912 538496 239924
rect 538548 239912 538554 239964
rect 441430 239884 441436 239896
rect 431926 239856 441436 239884
rect 441430 239844 441436 239856
rect 441488 239844 441494 239896
rect 441525 239887 441583 239893
rect 441525 239853 441537 239887
rect 441571 239884 441583 239887
rect 538306 239884 538312 239896
rect 441571 239856 538312 239884
rect 441571 239853 441583 239856
rect 441525 239847 441583 239853
rect 538306 239844 538312 239856
rect 538364 239844 538370 239896
rect 258442 239776 258448 239828
rect 258500 239816 258506 239828
rect 284294 239816 284300 239828
rect 258500 239788 284300 239816
rect 258500 239776 258506 239788
rect 284294 239776 284300 239788
rect 284352 239776 284358 239828
rect 439774 239776 439780 239828
rect 439832 239816 439838 239828
rect 467834 239816 467840 239828
rect 439832 239788 467840 239816
rect 439832 239776 439838 239788
rect 467834 239776 467840 239788
rect 467892 239776 467898 239828
rect 437382 239708 437388 239760
rect 437440 239748 437446 239760
rect 472066 239748 472072 239760
rect 437440 239720 472072 239748
rect 437440 239708 437446 239720
rect 472066 239708 472072 239720
rect 472124 239708 472130 239760
rect 274174 239640 274180 239692
rect 274232 239680 274238 239692
rect 456705 239683 456763 239689
rect 456705 239680 456717 239683
rect 274232 239652 456717 239680
rect 274232 239640 274238 239652
rect 456705 239649 456717 239652
rect 456751 239649 456763 239683
rect 456705 239643 456763 239649
rect 459554 239640 459560 239692
rect 459612 239680 459618 239692
rect 536926 239680 536932 239692
rect 459612 239652 536932 239680
rect 459612 239640 459618 239652
rect 536926 239640 536932 239652
rect 536984 239640 536990 239692
rect 273990 239572 273996 239624
rect 274048 239612 274054 239624
rect 465166 239612 465172 239624
rect 274048 239584 465172 239612
rect 274048 239572 274054 239584
rect 465166 239572 465172 239584
rect 465224 239572 465230 239624
rect 275554 239504 275560 239556
rect 275612 239544 275618 239556
rect 473354 239544 473360 239556
rect 275612 239516 473360 239544
rect 275612 239504 275618 239516
rect 473354 239504 473360 239516
rect 473412 239504 473418 239556
rect 274726 239436 274732 239488
rect 274784 239476 274790 239488
rect 476114 239476 476120 239488
rect 274784 239448 476120 239476
rect 274784 239436 274790 239448
rect 476114 239436 476120 239448
rect 476172 239436 476178 239488
rect 275370 239368 275376 239420
rect 275428 239408 275434 239420
rect 481726 239408 481732 239420
rect 275428 239380 481732 239408
rect 275428 239368 275434 239380
rect 481726 239368 481732 239380
rect 481784 239368 481790 239420
rect 437014 239300 437020 239352
rect 437072 239340 437078 239352
rect 441341 239343 441399 239349
rect 441341 239340 441353 239343
rect 437072 239312 441353 239340
rect 437072 239300 437078 239312
rect 441341 239309 441353 239312
rect 441387 239309 441399 239343
rect 441341 239303 441399 239309
rect 441525 239343 441583 239349
rect 441525 239309 441537 239343
rect 441571 239340 441583 239343
rect 522850 239340 522856 239352
rect 441571 239312 522856 239340
rect 441571 239309 441583 239312
rect 441525 239303 441583 239309
rect 522850 239300 522856 239312
rect 522908 239300 522914 239352
rect 438762 239232 438768 239284
rect 438820 239272 438826 239284
rect 441249 239275 441307 239281
rect 441249 239272 441261 239275
rect 438820 239244 441261 239272
rect 438820 239232 438826 239244
rect 441249 239241 441261 239244
rect 441295 239241 441307 239275
rect 522666 239272 522672 239284
rect 441249 239235 441307 239241
rect 441448 239244 522672 239272
rect 438670 239164 438676 239216
rect 438728 239204 438734 239216
rect 441448 239204 441476 239244
rect 522666 239232 522672 239244
rect 522724 239232 522730 239284
rect 438728 239176 441476 239204
rect 438728 239164 438734 239176
rect 441522 239164 441528 239216
rect 441580 239204 441586 239216
rect 523126 239204 523132 239216
rect 441580 239176 523132 239204
rect 441580 239164 441586 239176
rect 523126 239164 523132 239176
rect 523184 239164 523190 239216
rect 287790 239096 287796 239148
rect 287848 239136 287854 239148
rect 446398 239136 446404 239148
rect 287848 239108 446404 239136
rect 287848 239096 287854 239108
rect 446398 239096 446404 239108
rect 446456 239096 446462 239148
rect 447042 239096 447048 239148
rect 447100 239136 447106 239148
rect 537018 239136 537024 239148
rect 447100 239108 537024 239136
rect 447100 239096 447106 239108
rect 537018 239096 537024 239108
rect 537076 239096 537082 239148
rect 300578 239028 300584 239080
rect 300636 239068 300642 239080
rect 469214 239068 469220 239080
rect 300636 239040 469220 239068
rect 300636 239028 300642 239040
rect 469214 239028 469220 239040
rect 469272 239028 469278 239080
rect 299290 238960 299296 239012
rect 299348 239000 299354 239012
rect 483014 239000 483020 239012
rect 299348 238972 483020 239000
rect 299348 238960 299354 238972
rect 483014 238960 483020 238972
rect 483072 238960 483078 239012
rect 295150 238892 295156 238944
rect 295208 238932 295214 238944
rect 480438 238932 480444 238944
rect 295208 238904 480444 238932
rect 295208 238892 295214 238904
rect 480438 238892 480444 238904
rect 480496 238892 480502 238944
rect 288158 238824 288164 238876
rect 288216 238864 288222 238876
rect 479150 238864 479156 238876
rect 288216 238836 479156 238864
rect 288216 238824 288222 238836
rect 479150 238824 479156 238836
rect 479208 238824 479214 238876
rect 300394 238756 300400 238808
rect 300452 238796 300458 238808
rect 494238 238796 494244 238808
rect 300452 238768 494244 238796
rect 300452 238756 300458 238768
rect 494238 238756 494244 238768
rect 494296 238756 494302 238808
rect 288250 238688 288256 238740
rect 288308 238728 288314 238740
rect 476758 238728 476764 238740
rect 288308 238700 476764 238728
rect 288308 238688 288314 238700
rect 476758 238688 476764 238700
rect 476816 238688 476822 238740
rect 299106 238620 299112 238672
rect 299164 238660 299170 238672
rect 487798 238660 487804 238672
rect 299164 238632 487804 238660
rect 299164 238620 299170 238632
rect 487798 238620 487804 238632
rect 487856 238620 487862 238672
rect 300486 238552 300492 238604
rect 300544 238592 300550 238604
rect 490558 238592 490564 238604
rect 300544 238564 490564 238592
rect 300544 238552 300550 238564
rect 490558 238552 490564 238564
rect 490616 238552 490622 238604
rect 295058 238484 295064 238536
rect 295116 238524 295122 238536
rect 485406 238524 485412 238536
rect 295116 238496 485412 238524
rect 295116 238484 295122 238496
rect 485406 238484 485412 238496
rect 485464 238484 485470 238536
rect 292114 238416 292120 238468
rect 292172 238456 292178 238468
rect 484854 238456 484860 238468
rect 292172 238428 484860 238456
rect 292172 238416 292178 238428
rect 484854 238416 484860 238428
rect 484912 238416 484918 238468
rect 293586 238348 293592 238400
rect 293644 238388 293650 238400
rect 491662 238388 491668 238400
rect 293644 238360 491668 238388
rect 293644 238348 293650 238360
rect 491662 238348 491668 238360
rect 491720 238348 491726 238400
rect 293494 238280 293500 238332
rect 293552 238320 293558 238332
rect 492766 238320 492772 238332
rect 293552 238292 492772 238320
rect 293552 238280 293558 238292
rect 492766 238280 492772 238292
rect 492824 238280 492830 238332
rect 288066 238212 288072 238264
rect 288124 238252 288130 238264
rect 496814 238252 496820 238264
rect 288124 238224 496820 238252
rect 288124 238212 288130 238224
rect 496814 238212 496820 238224
rect 496872 238212 496878 238264
rect 260006 238144 260012 238196
rect 260064 238184 260070 238196
rect 287054 238184 287060 238196
rect 260064 238156 287060 238184
rect 260064 238144 260070 238156
rect 287054 238144 287060 238156
rect 287112 238144 287118 238196
rect 287974 238144 287980 238196
rect 288032 238184 288038 238196
rect 499206 238184 499212 238196
rect 288032 238156 499212 238184
rect 288032 238144 288038 238156
rect 499206 238144 499212 238156
rect 499264 238144 499270 238196
rect 232590 238076 232596 238128
rect 232648 238116 232654 238128
rect 465074 238116 465080 238128
rect 232648 238088 465080 238116
rect 232648 238076 232654 238088
rect 465074 238076 465080 238088
rect 465132 238076 465138 238128
rect 232682 238008 232688 238060
rect 232740 238048 232746 238060
rect 468294 238048 468300 238060
rect 232740 238020 468300 238048
rect 232740 238008 232746 238020
rect 468294 238008 468300 238020
rect 468352 238008 468358 238060
rect 288342 237940 288348 237992
rect 288400 237980 288406 237992
rect 475654 237980 475660 237992
rect 288400 237952 475660 237980
rect 288400 237940 288406 237952
rect 475654 237940 475660 237952
rect 475712 237940 475718 237992
rect 294598 237872 294604 237924
rect 294656 237912 294662 237924
rect 471790 237912 471796 237924
rect 294656 237884 471796 237912
rect 294656 237872 294662 237884
rect 471790 237872 471796 237884
rect 471848 237872 471854 237924
rect 294782 237804 294788 237856
rect 294840 237844 294846 237856
rect 467190 237844 467196 237856
rect 294840 237816 467196 237844
rect 294840 237804 294846 237816
rect 467190 237804 467196 237816
rect 467248 237804 467254 237856
rect 294874 237736 294880 237788
rect 294932 237776 294938 237788
rect 470686 237776 470692 237788
rect 294932 237748 470692 237776
rect 294932 237736 294938 237748
rect 470686 237736 470692 237748
rect 470744 237736 470750 237788
rect 293310 237668 293316 237720
rect 293368 237708 293374 237720
rect 463694 237708 463700 237720
rect 293368 237680 463700 237708
rect 293368 237668 293374 237680
rect 463694 237668 463700 237680
rect 463752 237668 463758 237720
rect 352558 237600 352564 237652
rect 352616 237640 352622 237652
rect 481634 237640 481640 237652
rect 352616 237612 481640 237640
rect 352616 237600 352622 237612
rect 481634 237600 481640 237612
rect 481692 237600 481698 237652
rect 438210 237532 438216 237584
rect 438268 237572 438274 237584
rect 500954 237572 500960 237584
rect 438268 237544 500960 237572
rect 438268 237532 438274 237544
rect 500954 237532 500960 237544
rect 501012 237532 501018 237584
rect 439682 237464 439688 237516
rect 439740 237504 439746 237516
rect 492674 237504 492680 237516
rect 439740 237476 492680 237504
rect 439740 237464 439746 237476
rect 492674 237464 492680 237476
rect 492732 237464 492738 237516
rect 438118 237396 438124 237448
rect 438176 237436 438182 237448
rect 481910 237436 481916 237448
rect 438176 237408 481916 237436
rect 438176 237396 438182 237408
rect 481910 237396 481916 237408
rect 481968 237396 481974 237448
rect 438578 237328 438584 237380
rect 438636 237368 438642 237380
rect 471974 237368 471980 237380
rect 438636 237340 471980 237368
rect 438636 237328 438642 237340
rect 471974 237328 471980 237340
rect 472032 237328 472038 237380
rect 472066 237328 472072 237380
rect 472124 237368 472130 237380
rect 523034 237368 523040 237380
rect 472124 237340 523040 237368
rect 472124 237328 472130 237340
rect 523034 237328 523040 237340
rect 523092 237328 523098 237380
rect 287882 237260 287888 237312
rect 287940 237300 287946 237312
rect 495434 237300 495440 237312
rect 287940 237272 495440 237300
rect 287940 237260 287946 237272
rect 495434 237260 495440 237272
rect 495492 237260 495498 237312
rect 285490 237192 285496 237244
rect 285548 237232 285554 237244
rect 493318 237232 493324 237244
rect 285548 237204 493324 237232
rect 285548 237192 285554 237204
rect 493318 237192 493324 237204
rect 493376 237192 493382 237244
rect 285398 237124 285404 237176
rect 285456 237164 285462 237176
rect 487154 237164 487160 237176
rect 285456 237136 487160 237164
rect 285456 237124 285462 237136
rect 487154 237124 487160 237136
rect 487212 237124 487218 237176
rect 296346 237056 296352 237108
rect 296404 237096 296410 237108
rect 496814 237096 496820 237108
rect 296404 237068 496820 237096
rect 296404 237056 296410 237068
rect 496814 237056 496820 237068
rect 496872 237056 496878 237108
rect 300210 236988 300216 237040
rect 300268 237028 300274 237040
rect 499850 237028 499856 237040
rect 300268 237000 499856 237028
rect 300268 236988 300274 237000
rect 499850 236988 499856 237000
rect 499908 236988 499914 237040
rect 284754 236920 284760 236972
rect 284812 236960 284818 236972
rect 483014 236960 483020 236972
rect 284812 236932 483020 236960
rect 284812 236920 284818 236932
rect 483014 236920 483020 236932
rect 483072 236920 483078 236972
rect 296438 236852 296444 236904
rect 296496 236892 296502 236904
rect 488534 236892 488540 236904
rect 296496 236864 488540 236892
rect 296496 236852 296502 236864
rect 488534 236852 488540 236864
rect 488592 236852 488598 236904
rect 300302 236784 300308 236836
rect 300360 236824 300366 236836
rect 491294 236824 491300 236836
rect 300360 236796 491300 236824
rect 300360 236784 300366 236796
rect 491294 236784 491300 236796
rect 491352 236784 491358 236836
rect 294966 236716 294972 236768
rect 295024 236756 295030 236768
rect 484394 236756 484400 236768
rect 295024 236728 484400 236756
rect 295024 236716 295030 236728
rect 484394 236716 484400 236728
rect 484452 236716 484458 236768
rect 296530 236648 296536 236700
rect 296588 236688 296594 236700
rect 485774 236688 485780 236700
rect 296588 236660 485780 236688
rect 296588 236648 296594 236660
rect 485774 236648 485780 236660
rect 485832 236648 485838 236700
rect 292298 236580 292304 236632
rect 292356 236620 292362 236632
rect 480254 236620 480260 236632
rect 292356 236592 480260 236620
rect 292356 236580 292362 236592
rect 480254 236580 480260 236592
rect 480312 236580 480318 236632
rect 292390 236512 292396 236564
rect 292448 236552 292454 236564
rect 480530 236552 480536 236564
rect 292448 236524 480536 236552
rect 292448 236512 292454 236524
rect 480530 236512 480536 236524
rect 480588 236512 480594 236564
rect 299198 236444 299204 236496
rect 299256 236484 299262 236496
rect 477494 236484 477500 236496
rect 299256 236456 477500 236484
rect 299256 236444 299262 236456
rect 477494 236444 477500 236456
rect 477552 236444 477558 236496
rect 297542 236376 297548 236428
rect 297600 236416 297606 236428
rect 473446 236416 473452 236428
rect 297600 236388 473452 236416
rect 297600 236376 297606 236388
rect 473446 236376 473452 236388
rect 473504 236376 473510 236428
rect 297634 236308 297640 236360
rect 297692 236348 297698 236360
rect 472066 236348 472072 236360
rect 297692 236320 472072 236348
rect 297692 236308 297698 236320
rect 472066 236308 472072 236320
rect 472124 236308 472130 236360
rect 297726 236240 297732 236292
rect 297784 236280 297790 236292
rect 471974 236280 471980 236292
rect 297784 236252 471980 236280
rect 297784 236240 297790 236252
rect 471974 236240 471980 236252
rect 472032 236240 472038 236292
rect 298922 236172 298928 236224
rect 298980 236212 298986 236224
rect 460934 236212 460940 236224
rect 298980 236184 460940 236212
rect 298980 236172 298986 236184
rect 460934 236172 460940 236184
rect 460992 236172 460998 236224
rect 461578 236172 461584 236224
rect 461636 236212 461642 236224
rect 485774 236212 485780 236224
rect 461636 236184 485780 236212
rect 461636 236172 461642 236184
rect 485774 236172 485780 236184
rect 485832 236172 485838 236224
rect 364334 236104 364340 236156
rect 364392 236144 364398 236156
rect 477586 236144 477592 236156
rect 364392 236116 477592 236144
rect 364392 236104 364398 236116
rect 477586 236104 477592 236116
rect 477644 236104 477650 236156
rect 232498 236036 232504 236088
rect 232556 236076 232562 236088
rect 456705 236079 456763 236085
rect 232556 236048 447134 236076
rect 232556 236036 232562 236048
rect 447106 236008 447134 236048
rect 456705 236045 456717 236079
rect 456751 236076 456763 236079
rect 462314 236076 462320 236088
rect 456751 236048 462320 236076
rect 456751 236045 456763 236048
rect 456705 236039 456763 236045
rect 462314 236036 462320 236048
rect 462372 236036 462378 236088
rect 462406 236008 462412 236020
rect 447106 235980 462412 236008
rect 462406 235968 462412 235980
rect 462464 235968 462470 236020
rect 297358 235900 297364 235952
rect 297416 235940 297422 235952
rect 505094 235940 505100 235952
rect 297416 235912 505100 235940
rect 297416 235900 297422 235912
rect 505094 235900 505100 235912
rect 505152 235900 505158 235952
rect 296254 235832 296260 235884
rect 296312 235872 296318 235884
rect 503714 235872 503720 235884
rect 296312 235844 503720 235872
rect 296312 235832 296318 235844
rect 503714 235832 503720 235844
rect 503772 235832 503778 235884
rect 296162 235764 296168 235816
rect 296220 235804 296226 235816
rect 502426 235804 502432 235816
rect 296220 235776 502432 235804
rect 296220 235764 296226 235776
rect 502426 235764 502432 235776
rect 502484 235764 502490 235816
rect 296622 235696 296628 235748
rect 296680 235736 296686 235748
rect 469214 235736 469220 235748
rect 296680 235708 469220 235736
rect 296680 235696 296686 235708
rect 469214 235696 469220 235708
rect 469272 235696 469278 235748
rect 276382 235356 276388 235408
rect 276440 235396 276446 235408
rect 440234 235396 440240 235408
rect 276440 235368 440240 235396
rect 276440 235356 276446 235368
rect 440234 235356 440240 235368
rect 440292 235356 440298 235408
rect 272794 235288 272800 235340
rect 272852 235328 272858 235340
rect 445754 235328 445760 235340
rect 272852 235300 445760 235328
rect 272852 235288 272858 235300
rect 445754 235288 445760 235300
rect 445812 235288 445818 235340
rect 280522 235220 280528 235272
rect 280580 235260 280586 235272
rect 505094 235260 505100 235272
rect 280580 235232 505100 235260
rect 280580 235220 280586 235232
rect 505094 235220 505100 235232
rect 505152 235220 505158 235272
rect 286962 233180 286968 233232
rect 287020 233220 287026 233232
rect 579982 233220 579988 233232
rect 287020 233192 579988 233220
rect 287020 233180 287026 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 289722 219376 289728 219428
rect 289780 219416 289786 219428
rect 579982 219416 579988 219428
rect 289780 219388 579988 219416
rect 289780 219376 289786 219388
rect 579982 219376 579988 219388
rect 580040 219376 580046 219428
rect 2958 202784 2964 202836
rect 3016 202824 3022 202836
rect 6546 202824 6552 202836
rect 3016 202796 6552 202824
rect 3016 202784 3022 202796
rect 6546 202784 6552 202796
rect 6604 202784 6610 202836
rect 298738 193128 298744 193180
rect 298796 193168 298802 193180
rect 579614 193168 579620 193180
rect 298796 193140 579620 193168
rect 298796 193128 298802 193140
rect 579614 193128 579620 193140
rect 579672 193128 579678 193180
rect 2774 188912 2780 188964
rect 2832 188952 2838 188964
rect 5166 188952 5172 188964
rect 2832 188924 5172 188952
rect 2832 188912 2838 188924
rect 5166 188912 5172 188924
rect 5224 188912 5230 188964
rect 289630 179324 289636 179376
rect 289688 179364 289694 179376
rect 579614 179364 579620 179376
rect 289688 179336 579620 179364
rect 289688 179324 289694 179336
rect 579614 179324 579620 179336
rect 579672 179324 579678 179376
rect 108942 177624 108948 177676
rect 109000 177664 109006 177676
rect 243354 177664 243360 177676
rect 109000 177636 243360 177664
rect 109000 177624 109006 177636
rect 243354 177624 243360 177636
rect 243412 177624 243418 177676
rect 104802 177556 104808 177608
rect 104860 177596 104866 177608
rect 243262 177596 243268 177608
rect 104860 177568 243268 177596
rect 104860 177556 104866 177568
rect 243262 177556 243268 177568
rect 243320 177556 243326 177608
rect 268562 177556 268568 177608
rect 268620 177596 268626 177608
rect 402974 177596 402980 177608
rect 268620 177568 402980 177596
rect 268620 177556 268626 177568
rect 402974 177556 402980 177568
rect 403032 177556 403038 177608
rect 64782 177488 64788 177540
rect 64840 177528 64846 177540
rect 240870 177528 240876 177540
rect 64840 177500 240876 177528
rect 64840 177488 64846 177500
rect 240870 177488 240876 177500
rect 240928 177488 240934 177540
rect 269666 177488 269672 177540
rect 269724 177528 269730 177540
rect 416774 177528 416780 177540
rect 269724 177500 416780 177528
rect 269724 177488 269730 177500
rect 416774 177488 416780 177500
rect 416832 177488 416838 177540
rect 53650 177420 53656 177472
rect 53708 177460 53714 177472
rect 239214 177460 239220 177472
rect 53708 177432 239220 177460
rect 53708 177420 53714 177432
rect 239214 177420 239220 177432
rect 239272 177420 239278 177472
rect 271046 177420 271052 177472
rect 271104 177460 271110 177472
rect 434714 177460 434720 177472
rect 271104 177432 434720 177460
rect 271104 177420 271110 177432
rect 434714 177420 434720 177432
rect 434772 177420 434778 177472
rect 9582 177352 9588 177404
rect 9640 177392 9646 177404
rect 234890 177392 234896 177404
rect 9640 177364 234896 177392
rect 9640 177352 9646 177364
rect 234890 177352 234896 177364
rect 234948 177352 234954 177404
rect 280706 177352 280712 177404
rect 280764 177392 280770 177404
rect 540974 177392 540980 177404
rect 280764 177364 540980 177392
rect 280764 177352 280770 177364
rect 540974 177352 540980 177364
rect 541032 177352 541038 177404
rect 4062 177284 4068 177336
rect 4120 177324 4126 177336
rect 234982 177324 234988 177336
rect 4120 177296 234988 177324
rect 4120 177284 4126 177296
rect 234982 177284 234988 177296
rect 235040 177284 235046 177336
rect 280614 177284 280620 177336
rect 280672 177324 280678 177336
rect 549254 177324 549260 177336
rect 280672 177296 549260 177324
rect 280672 177284 280678 177296
rect 549254 177284 549260 177296
rect 549312 177284 549318 177336
rect 274082 162120 274088 162172
rect 274140 162160 274146 162172
rect 444374 162160 444380 162172
rect 274140 162132 444380 162160
rect 274140 162120 274146 162132
rect 444374 162120 444380 162132
rect 444432 162120 444438 162172
rect 286870 153144 286876 153196
rect 286928 153184 286934 153196
rect 580166 153184 580172 153196
rect 286928 153156 580172 153184
rect 286928 153144 286934 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3142 150356 3148 150408
rect 3200 150396 3206 150408
rect 6454 150396 6460 150408
rect 3200 150368 6460 150396
rect 3200 150356 3206 150368
rect 6454 150356 6460 150368
rect 6512 150356 6518 150408
rect 286778 139340 286784 139392
rect 286836 139380 286842 139392
rect 580166 139380 580172 139392
rect 286836 139352 580172 139380
rect 286836 139340 286842 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 2774 137232 2780 137284
rect 2832 137272 2838 137284
rect 5074 137272 5080 137284
rect 2832 137244 5080 137272
rect 2832 137232 2838 137244
rect 5074 137232 5080 137244
rect 5132 137232 5138 137284
rect 286686 126896 286692 126948
rect 286744 126936 286750 126948
rect 579614 126936 579620 126948
rect 286744 126908 579620 126936
rect 286744 126896 286750 126908
rect 579614 126896 579620 126908
rect 579672 126896 579678 126948
rect 286594 100648 286600 100700
rect 286652 100688 286658 100700
rect 580166 100688 580172 100700
rect 286652 100660 580172 100688
rect 286652 100648 286658 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3234 97860 3240 97912
rect 3292 97900 3298 97912
rect 6362 97900 6368 97912
rect 3292 97872 6368 97900
rect 3292 97860 3298 97872
rect 6362 97860 6368 97872
rect 6420 97860 6426 97912
rect 219250 89088 219256 89140
rect 219308 89128 219314 89140
rect 253198 89128 253204 89140
rect 219308 89100 253204 89128
rect 219308 89088 219314 89100
rect 253198 89088 253204 89100
rect 253256 89088 253262 89140
rect 210970 89020 210976 89072
rect 211028 89060 211034 89072
rect 253290 89060 253296 89072
rect 211028 89032 253296 89060
rect 211028 89020 211034 89032
rect 253290 89020 253296 89032
rect 253348 89020 253354 89072
rect 258810 89020 258816 89072
rect 258868 89060 258874 89072
rect 284386 89060 284392 89072
rect 258868 89032 284392 89060
rect 258868 89020 258874 89032
rect 284386 89020 284392 89032
rect 284444 89020 284450 89072
rect 202690 88952 202696 89004
rect 202748 88992 202754 89004
rect 251818 88992 251824 89004
rect 202748 88964 251824 88992
rect 202748 88952 202754 88964
rect 251818 88952 251824 88964
rect 251876 88952 251882 89004
rect 270770 88952 270776 89004
rect 270828 88992 270834 89004
rect 420914 88992 420920 89004
rect 270828 88964 420920 88992
rect 270828 88952 270834 88964
rect 420914 88952 420920 88964
rect 420972 88952 420978 89004
rect 253382 88680 253388 88732
rect 253440 88720 253446 88732
rect 256142 88720 256148 88732
rect 253440 88692 256148 88720
rect 253440 88680 253446 88692
rect 256142 88680 256148 88692
rect 256200 88680 256206 88732
rect 253198 88272 253204 88324
rect 253256 88312 253262 88324
rect 254486 88312 254492 88324
rect 253256 88284 254492 88312
rect 253256 88272 253262 88284
rect 254486 88272 254492 88284
rect 254544 88272 254550 88324
rect 260282 87796 260288 87848
rect 260340 87836 260346 87848
rect 302234 87836 302240 87848
rect 260340 87808 302240 87836
rect 260340 87796 260346 87808
rect 302234 87796 302240 87808
rect 302292 87796 302298 87848
rect 200022 87728 200028 87780
rect 200080 87768 200086 87780
rect 251726 87768 251732 87780
rect 200080 87740 251732 87768
rect 200080 87728 200086 87740
rect 251726 87728 251732 87740
rect 251784 87728 251790 87780
rect 268654 87728 268660 87780
rect 268712 87768 268718 87780
rect 389174 87768 389180 87780
rect 268712 87740 389180 87768
rect 268712 87728 268718 87740
rect 389174 87728 389180 87740
rect 389232 87728 389238 87780
rect 115842 87660 115848 87712
rect 115900 87700 115906 87712
rect 244826 87700 244832 87712
rect 115900 87672 244832 87700
rect 115900 87660 115906 87672
rect 244826 87660 244832 87672
rect 244884 87660 244890 87712
rect 269942 87660 269948 87712
rect 270000 87700 270006 87712
rect 407206 87700 407212 87712
rect 270000 87672 407212 87700
rect 270000 87660 270006 87672
rect 407206 87660 407212 87672
rect 407264 87660 407270 87712
rect 84102 87592 84108 87644
rect 84160 87632 84166 87644
rect 242066 87632 242072 87644
rect 84160 87604 242072 87632
rect 84160 87592 84166 87604
rect 242066 87592 242072 87604
rect 242124 87592 242130 87644
rect 274266 87592 274272 87644
rect 274324 87632 274330 87644
rect 456794 87632 456800 87644
rect 274324 87604 456800 87632
rect 274324 87592 274330 87604
rect 456794 87592 456800 87604
rect 456852 87592 456858 87644
rect 285122 86912 285128 86964
rect 285180 86952 285186 86964
rect 579614 86952 579620 86964
rect 285180 86924 579620 86952
rect 285180 86912 285186 86924
rect 579614 86912 579620 86924
rect 579672 86912 579678 86964
rect 216582 86436 216588 86488
rect 216640 86476 216646 86488
rect 253106 86476 253112 86488
rect 216640 86448 253112 86476
rect 216640 86436 216646 86448
rect 253106 86436 253112 86448
rect 253164 86436 253170 86488
rect 195882 86368 195888 86420
rect 195940 86408 195946 86420
rect 251634 86408 251640 86420
rect 195940 86380 251640 86408
rect 195940 86368 195946 86380
rect 251634 86368 251640 86380
rect 251692 86368 251698 86420
rect 102042 86300 102048 86352
rect 102100 86340 102106 86352
rect 243170 86340 243176 86352
rect 102100 86312 243176 86340
rect 102100 86300 102106 86312
rect 243170 86300 243176 86312
rect 243228 86300 243234 86352
rect 49602 86232 49608 86284
rect 49660 86272 49666 86284
rect 239122 86272 239128 86284
rect 49660 86244 239128 86272
rect 49660 86232 49666 86244
rect 239122 86232 239128 86244
rect 239180 86232 239186 86284
rect 2774 85212 2780 85264
rect 2832 85252 2838 85264
rect 4982 85252 4988 85264
rect 2832 85224 4988 85252
rect 2832 85212 2838 85224
rect 4982 85212 4988 85224
rect 5040 85212 5046 85264
rect 212442 85076 212448 85128
rect 212500 85116 212506 85128
rect 253014 85116 253020 85128
rect 212500 85088 253020 85116
rect 212500 85076 212506 85088
rect 253014 85076 253020 85088
rect 253072 85076 253078 85128
rect 260926 85076 260932 85128
rect 260984 85116 260990 85128
rect 307846 85116 307852 85128
rect 260984 85088 307852 85116
rect 260984 85076 260990 85088
rect 307846 85076 307852 85088
rect 307904 85076 307910 85128
rect 162762 85008 162768 85060
rect 162820 85048 162826 85060
rect 249150 85048 249156 85060
rect 162820 85020 249156 85048
rect 162820 85008 162826 85020
rect 249150 85008 249156 85020
rect 249208 85008 249214 85060
rect 266998 85008 267004 85060
rect 267056 85048 267062 85060
rect 332594 85048 332600 85060
rect 267056 85020 332600 85048
rect 267056 85008 267062 85020
rect 332594 85008 332600 85020
rect 332652 85008 332658 85060
rect 111702 84940 111708 84992
rect 111760 84980 111766 84992
rect 244734 84980 244740 84992
rect 111760 84952 244740 84980
rect 111760 84940 111766 84952
rect 244734 84940 244740 84952
rect 244792 84940 244798 84992
rect 252462 84940 252468 84992
rect 252520 84980 252526 84992
rect 256050 84980 256056 84992
rect 252520 84952 256056 84980
rect 252520 84940 252526 84952
rect 256050 84940 256056 84952
rect 256108 84940 256114 84992
rect 264146 84940 264152 84992
rect 264204 84980 264210 84992
rect 349154 84980 349160 84992
rect 264204 84952 349160 84980
rect 264204 84940 264210 84952
rect 349154 84940 349160 84952
rect 349212 84940 349218 84992
rect 79962 84872 79968 84924
rect 80020 84912 80026 84924
rect 241974 84912 241980 84924
rect 80020 84884 241980 84912
rect 80020 84872 80026 84884
rect 241974 84872 241980 84884
rect 242032 84872 242038 84924
rect 265342 84872 265348 84924
rect 265400 84912 265406 84924
rect 369854 84912 369860 84924
rect 265400 84884 369860 84912
rect 265400 84872 265406 84884
rect 369854 84872 369860 84884
rect 369912 84872 369918 84924
rect 77202 84804 77208 84856
rect 77260 84844 77266 84856
rect 240778 84844 240784 84856
rect 77260 84816 240784 84844
rect 77260 84804 77266 84816
rect 240778 84804 240784 84816
rect 240836 84804 240842 84856
rect 272058 84804 272064 84856
rect 272116 84844 272122 84856
rect 452654 84844 452660 84856
rect 272116 84816 452660 84844
rect 272116 84804 272122 84816
rect 452654 84804 452660 84816
rect 452712 84804 452718 84856
rect 276474 83580 276480 83632
rect 276532 83620 276538 83632
rect 488534 83620 488540 83632
rect 276532 83592 488540 83620
rect 276532 83580 276538 83592
rect 488534 83580 488540 83592
rect 488592 83580 488598 83632
rect 160002 83512 160008 83564
rect 160060 83552 160066 83564
rect 247494 83552 247500 83564
rect 160060 83524 247500 83552
rect 160060 83512 160066 83524
rect 247494 83512 247500 83524
rect 247552 83512 247558 83564
rect 278038 83512 278044 83564
rect 278096 83552 278102 83564
rect 506474 83552 506480 83564
rect 278096 83524 506480 83552
rect 278096 83512 278102 83524
rect 506474 83512 506480 83524
rect 506532 83512 506538 83564
rect 135162 83444 135168 83496
rect 135220 83484 135226 83496
rect 246390 83484 246396 83496
rect 135220 83456 246396 83484
rect 135220 83444 135226 83456
rect 246390 83444 246396 83456
rect 246448 83444 246454 83496
rect 279602 83444 279608 83496
rect 279660 83484 279666 83496
rect 531314 83484 531320 83496
rect 279660 83456 531320 83484
rect 279660 83444 279666 83456
rect 531314 83444 531320 83456
rect 531372 83444 531378 83496
rect 184842 82084 184848 82136
rect 184900 82124 184906 82136
rect 250438 82124 250444 82136
rect 184900 82096 250444 82124
rect 184900 82084 184906 82096
rect 250438 82084 250444 82096
rect 250496 82084 250502 82136
rect 272978 82084 272984 82136
rect 273036 82124 273042 82136
rect 448606 82124 448612 82136
rect 273036 82096 448612 82124
rect 273036 82084 273042 82096
rect 448606 82084 448612 82096
rect 448664 82084 448670 82136
rect 234522 80860 234528 80912
rect 234580 80900 234586 80912
rect 254394 80900 254400 80912
rect 234580 80872 254400 80900
rect 234580 80860 234586 80872
rect 254394 80860 254400 80872
rect 254452 80860 254458 80912
rect 261754 80860 261760 80912
rect 261812 80900 261818 80912
rect 320174 80900 320180 80912
rect 261812 80872 320180 80900
rect 261812 80860 261818 80872
rect 320174 80860 320180 80872
rect 320232 80860 320238 80912
rect 155862 80792 155868 80844
rect 155920 80832 155926 80844
rect 247402 80832 247408 80844
rect 155920 80804 247408 80832
rect 155920 80792 155926 80804
rect 247402 80792 247408 80804
rect 247460 80792 247466 80844
rect 264054 80792 264060 80844
rect 264112 80832 264118 80844
rect 345014 80832 345020 80844
rect 264112 80804 345020 80832
rect 264112 80792 264118 80804
rect 345014 80792 345020 80804
rect 345072 80792 345078 80844
rect 131022 80724 131028 80776
rect 131080 80764 131086 80776
rect 246298 80764 246304 80776
rect 131080 80736 246304 80764
rect 131080 80724 131086 80736
rect 246298 80724 246304 80736
rect 246356 80724 246362 80776
rect 264974 80724 264980 80776
rect 265032 80764 265038 80776
rect 365714 80764 365720 80776
rect 265032 80736 365720 80764
rect 265032 80724 265038 80736
rect 365714 80724 365720 80736
rect 365772 80724 365778 80776
rect 73062 80656 73068 80708
rect 73120 80696 73126 80708
rect 240686 80696 240692 80708
rect 73120 80668 240692 80696
rect 73120 80656 73126 80668
rect 240686 80656 240692 80668
rect 240744 80656 240750 80708
rect 267090 80656 267096 80708
rect 267148 80696 267154 80708
rect 385034 80696 385040 80708
rect 267148 80668 385040 80696
rect 267148 80656 267154 80668
rect 385034 80656 385040 80668
rect 385092 80656 385098 80708
rect 275646 79296 275652 79348
rect 275704 79336 275710 79348
rect 470594 79336 470600 79348
rect 275704 79308 470600 79336
rect 275704 79296 275710 79308
rect 470594 79296 470600 79308
rect 470652 79296 470658 79348
rect 286502 73108 286508 73160
rect 286560 73148 286566 73160
rect 580166 73148 580172 73160
rect 286560 73120 580172 73148
rect 286560 73108 286566 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 2958 59168 2964 59220
rect 3016 59208 3022 59220
rect 6270 59208 6276 59220
rect 3016 59180 6276 59208
rect 3016 59168 3022 59180
rect 6270 59168 6276 59180
rect 6328 59168 6334 59220
rect 2774 45500 2780 45552
rect 2832 45540 2838 45552
rect 4890 45540 4896 45552
rect 2832 45512 4896 45540
rect 2832 45500 2838 45512
rect 4890 45500 4896 45512
rect 4948 45500 4954 45552
rect 286318 33056 286324 33108
rect 286376 33096 286382 33108
rect 580166 33096 580172 33108
rect 286376 33068 580172 33096
rect 286376 33056 286382 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 311158 20612 311164 20664
rect 311216 20652 311222 20664
rect 579982 20652 579988 20664
rect 311216 20624 579988 20652
rect 311216 20612 311222 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 2958 19456 2964 19508
rect 3016 19496 3022 19508
rect 6178 19496 6184 19508
rect 3016 19468 6184 19496
rect 3016 19456 3022 19468
rect 6178 19456 6184 19468
rect 6236 19456 6242 19508
rect 340966 16532 340972 16584
rect 341024 16572 341030 16584
rect 342162 16572 342168 16584
rect 341024 16544 342168 16572
rect 341024 16532 341030 16544
rect 342162 16532 342168 16544
rect 342220 16532 342226 16584
rect 448606 13268 448612 13320
rect 448664 13308 448670 13320
rect 449802 13308 449808 13320
rect 448664 13280 449808 13308
rect 448664 13268 448670 13280
rect 449802 13268 449808 13280
rect 449860 13268 449866 13320
rect 193214 11704 193220 11756
rect 193272 11744 193278 11756
rect 194410 11744 194416 11756
rect 193272 11716 194416 11744
rect 193272 11704 193278 11716
rect 194410 11704 194416 11716
rect 194468 11704 194474 11756
rect 209774 11704 209780 11756
rect 209832 11744 209838 11756
rect 210970 11744 210976 11756
rect 209832 11716 210976 11744
rect 209832 11704 209838 11716
rect 210970 11704 210976 11716
rect 211028 11704 211034 11756
rect 235810 11704 235816 11756
rect 235868 11744 235874 11756
rect 250530 11744 250536 11756
rect 235868 11716 250536 11744
rect 235868 11704 235874 11716
rect 250530 11704 250536 11716
rect 250588 11704 250594 11756
rect 271230 11704 271236 11756
rect 271288 11744 271294 11756
rect 271506 11744 271512 11756
rect 271288 11716 271512 11744
rect 271288 11704 271294 11716
rect 271506 11704 271512 11716
rect 271564 11704 271570 11756
rect 284294 11704 284300 11756
rect 284352 11744 284358 11756
rect 285398 11744 285404 11756
rect 284352 11716 285404 11744
rect 284352 11704 284358 11716
rect 285398 11704 285404 11716
rect 285456 11704 285462 11756
rect 316126 11704 316132 11756
rect 316184 11744 316190 11756
rect 317322 11744 317328 11756
rect 316184 11716 317328 11744
rect 316184 11704 316190 11716
rect 317322 11704 317328 11716
rect 317380 11704 317386 11756
rect 423766 11704 423772 11756
rect 423824 11744 423830 11756
rect 424962 11744 424968 11756
rect 423824 11716 424968 11744
rect 423824 11704 423830 11716
rect 424962 11704 424968 11716
rect 425020 11704 425026 11756
rect 262674 11636 262680 11688
rect 262732 11676 262738 11688
rect 274818 11676 274824 11688
rect 262732 11648 274824 11676
rect 262732 11636 262738 11648
rect 274818 11636 274824 11648
rect 274876 11636 274882 11688
rect 262950 10752 262956 10804
rect 263008 10792 263014 10804
rect 324314 10792 324320 10804
rect 263008 10764 324320 10792
rect 263008 10752 263014 10764
rect 324314 10752 324320 10764
rect 324372 10752 324378 10804
rect 262766 10684 262772 10736
rect 262824 10724 262830 10736
rect 328730 10724 328736 10736
rect 262824 10696 328736 10724
rect 262824 10684 262830 10696
rect 328730 10684 328736 10696
rect 328788 10684 328794 10736
rect 263042 10616 263048 10668
rect 263100 10656 263106 10668
rect 332686 10656 332692 10668
rect 263100 10628 332692 10656
rect 263100 10616 263106 10628
rect 332686 10616 332692 10628
rect 332744 10616 332750 10668
rect 262858 10548 262864 10600
rect 262916 10588 262922 10600
rect 336274 10588 336280 10600
rect 262916 10560 336280 10588
rect 262916 10548 262922 10560
rect 336274 10548 336280 10560
rect 336332 10548 336338 10600
rect 267366 10480 267372 10532
rect 267424 10520 267430 10532
rect 371234 10520 371240 10532
rect 267424 10492 371240 10520
rect 267424 10480 267430 10492
rect 371234 10480 371240 10492
rect 371292 10480 371298 10532
rect 267182 10412 267188 10464
rect 267240 10452 267246 10464
rect 373994 10452 374000 10464
rect 267240 10424 374000 10452
rect 267240 10412 267246 10424
rect 373994 10412 374000 10424
rect 374052 10412 374058 10464
rect 267274 10344 267280 10396
rect 267332 10384 267338 10396
rect 378410 10384 378416 10396
rect 267332 10356 378416 10384
rect 267332 10344 267338 10356
rect 378410 10344 378416 10356
rect 378468 10344 378474 10396
rect 267458 10276 267464 10328
rect 267516 10316 267522 10328
rect 382366 10316 382372 10328
rect 267516 10288 382372 10316
rect 267516 10276 267522 10288
rect 382366 10276 382372 10288
rect 382424 10276 382430 10328
rect 283558 9596 283564 9648
rect 283616 9636 283622 9648
rect 480530 9636 480536 9648
rect 283616 9608 480536 9636
rect 283616 9596 283622 9608
rect 480530 9596 480536 9608
rect 480588 9596 480594 9648
rect 283742 9528 283748 9580
rect 283800 9568 283806 9580
rect 487614 9568 487620 9580
rect 283800 9540 487620 9568
rect 283800 9528 283806 9540
rect 487614 9528 487620 9540
rect 487672 9528 487678 9580
rect 285214 9460 285220 9512
rect 285272 9500 285278 9512
rect 523034 9500 523040 9512
rect 285272 9472 523040 9500
rect 285272 9460 285278 9472
rect 523034 9460 523040 9472
rect 523092 9460 523098 9512
rect 285030 9392 285036 9444
rect 285088 9432 285094 9444
rect 530118 9432 530124 9444
rect 285088 9404 530124 9432
rect 285088 9392 285094 9404
rect 530118 9392 530124 9404
rect 530176 9392 530182 9444
rect 281074 9324 281080 9376
rect 281132 9364 281138 9376
rect 543182 9364 543188 9376
rect 281132 9336 543188 9364
rect 281132 9324 281138 9336
rect 543182 9324 543188 9336
rect 543240 9324 543246 9376
rect 280982 9256 280988 9308
rect 281040 9296 281046 9308
rect 546678 9296 546684 9308
rect 281040 9268 546684 9296
rect 281040 9256 281046 9268
rect 546678 9256 546684 9268
rect 546736 9256 546742 9308
rect 282362 9188 282368 9240
rect 282420 9228 282426 9240
rect 553762 9228 553768 9240
rect 282420 9200 553768 9228
rect 282420 9188 282426 9200
rect 553762 9188 553768 9200
rect 553820 9188 553826 9240
rect 253474 9120 253480 9172
rect 253532 9160 253538 9172
rect 255958 9160 255964 9172
rect 253532 9132 255964 9160
rect 253532 9120 253538 9132
rect 255958 9120 255964 9132
rect 256016 9120 256022 9172
rect 282086 9120 282092 9172
rect 282144 9160 282150 9172
rect 557350 9160 557356 9172
rect 282144 9132 557356 9160
rect 282144 9120 282150 9132
rect 557350 9120 557356 9132
rect 557408 9120 557414 9172
rect 282454 9052 282460 9104
rect 282512 9092 282518 9104
rect 560846 9092 560852 9104
rect 282512 9064 560852 9092
rect 282512 9052 282518 9064
rect 560846 9052 560852 9064
rect 560904 9052 560910 9104
rect 281994 8984 282000 9036
rect 282052 9024 282058 9036
rect 564434 9024 564440 9036
rect 282052 8996 564440 9024
rect 282052 8984 282058 8996
rect 564434 8984 564440 8996
rect 564492 8984 564498 9036
rect 283834 8916 283840 8968
rect 283892 8956 283898 8968
rect 573910 8956 573916 8968
rect 283892 8928 573916 8956
rect 283892 8916 283898 8928
rect 573910 8916 573916 8928
rect 573968 8916 573974 8968
rect 252462 8848 252468 8900
rect 252520 8888 252526 8900
rect 255866 8888 255872 8900
rect 252520 8860 255872 8888
rect 252520 8848 252526 8860
rect 255866 8848 255872 8860
rect 255924 8848 255930 8900
rect 272610 8848 272616 8900
rect 272668 8888 272674 8900
rect 452102 8888 452108 8900
rect 272668 8860 452108 8888
rect 272668 8848 272674 8860
rect 452102 8848 452108 8860
rect 452160 8848 452166 8900
rect 272518 8780 272524 8832
rect 272576 8820 272582 8832
rect 450906 8820 450912 8832
rect 272576 8792 450912 8820
rect 272576 8780 272582 8792
rect 450906 8780 450912 8792
rect 450964 8780 450970 8832
rect 273898 8712 273904 8764
rect 273956 8752 273962 8764
rect 440326 8752 440332 8764
rect 273956 8724 440332 8752
rect 273956 8712 273962 8724
rect 440326 8712 440332 8724
rect 440384 8712 440390 8764
rect 270034 8644 270040 8696
rect 270092 8684 270098 8696
rect 420178 8684 420184 8696
rect 270092 8656 420184 8684
rect 270092 8644 270098 8656
rect 420178 8644 420184 8656
rect 420236 8644 420242 8696
rect 270126 8576 270132 8628
rect 270184 8616 270190 8628
rect 415486 8616 415492 8628
rect 270184 8588 415492 8616
rect 270184 8576 270190 8588
rect 415486 8576 415492 8588
rect 415544 8576 415550 8628
rect 268746 8508 268752 8560
rect 268804 8548 268810 8560
rect 402514 8548 402520 8560
rect 268804 8520 402520 8548
rect 268804 8508 268810 8520
rect 402514 8508 402520 8520
rect 402572 8508 402578 8560
rect 269850 8440 269856 8492
rect 269908 8480 269914 8492
rect 387150 8480 387156 8492
rect 269908 8452 387156 8480
rect 269908 8440 269914 8452
rect 387150 8440 387156 8452
rect 387208 8440 387214 8492
rect 268378 8372 268384 8424
rect 268436 8412 268442 8424
rect 379974 8412 379980 8424
rect 268436 8384 379980 8412
rect 268436 8372 268442 8384
rect 379974 8372 379980 8384
rect 380032 8372 380038 8424
rect 271598 8304 271604 8356
rect 271656 8344 271662 8356
rect 365806 8344 365812 8356
rect 271656 8316 365812 8344
rect 271656 8304 271662 8316
rect 365806 8304 365812 8316
rect 365864 8304 365870 8356
rect 109310 8236 109316 8288
rect 109368 8276 109374 8288
rect 242250 8276 242256 8288
rect 109368 8248 242256 8276
rect 109368 8236 109374 8248
rect 242250 8236 242256 8248
rect 242308 8236 242314 8288
rect 276566 8236 276572 8288
rect 276624 8276 276630 8288
rect 493502 8276 493508 8288
rect 276624 8248 493508 8276
rect 276624 8236 276630 8248
rect 493502 8236 493508 8248
rect 493560 8236 493566 8288
rect 98638 8168 98644 8220
rect 98696 8208 98702 8220
rect 234338 8208 234344 8220
rect 98696 8180 234344 8208
rect 98696 8168 98702 8180
rect 234338 8168 234344 8180
rect 234396 8168 234402 8220
rect 276014 8168 276020 8220
rect 276072 8208 276078 8220
rect 497090 8208 497096 8220
rect 276072 8180 497096 8208
rect 276072 8168 276078 8180
rect 497090 8168 497096 8180
rect 497148 8168 497154 8220
rect 102226 8100 102232 8152
rect 102284 8140 102290 8152
rect 242158 8140 242164 8152
rect 102284 8112 242164 8140
rect 102284 8100 102290 8112
rect 242158 8100 242164 8112
rect 242216 8100 242222 8152
rect 277026 8100 277032 8152
rect 277084 8140 277090 8152
rect 500586 8140 500592 8152
rect 277084 8112 500592 8140
rect 277084 8100 277090 8112
rect 500586 8100 500592 8112
rect 500644 8100 500650 8152
rect 77386 8032 77392 8084
rect 77444 8072 77450 8084
rect 240502 8072 240508 8084
rect 77444 8044 240508 8072
rect 77444 8032 77450 8044
rect 240502 8032 240508 8044
rect 240560 8032 240566 8084
rect 278406 8032 278412 8084
rect 278464 8072 278470 8084
rect 504174 8072 504180 8084
rect 278464 8044 504180 8072
rect 278464 8032 278470 8044
rect 504174 8032 504180 8044
rect 504232 8032 504238 8084
rect 73798 7964 73804 8016
rect 73856 8004 73862 8016
rect 240410 8004 240416 8016
rect 73856 7976 240416 8004
rect 73856 7964 73862 7976
rect 240410 7964 240416 7976
rect 240468 7964 240474 8016
rect 278314 7964 278320 8016
rect 278372 8004 278378 8016
rect 507670 8004 507676 8016
rect 278372 7976 507676 8004
rect 278372 7964 278378 7976
rect 507670 7964 507676 7976
rect 507728 7964 507734 8016
rect 70210 7896 70216 7948
rect 70268 7936 70274 7948
rect 240594 7936 240600 7948
rect 70268 7908 240600 7936
rect 70268 7896 70274 7908
rect 240594 7896 240600 7908
rect 240652 7896 240658 7948
rect 278222 7896 278228 7948
rect 278280 7936 278286 7948
rect 511258 7936 511264 7948
rect 278280 7908 511264 7936
rect 278280 7896 278286 7908
rect 511258 7896 511264 7908
rect 511316 7896 511322 7948
rect 66714 7828 66720 7880
rect 66772 7868 66778 7880
rect 241238 7868 241244 7880
rect 66772 7840 241244 7868
rect 66772 7828 66778 7840
rect 241238 7828 241244 7840
rect 241296 7828 241302 7880
rect 278130 7828 278136 7880
rect 278188 7868 278194 7880
rect 514754 7868 514760 7880
rect 278188 7840 514760 7868
rect 278188 7828 278194 7840
rect 514754 7828 514760 7840
rect 514812 7828 514818 7880
rect 63218 7760 63224 7812
rect 63276 7800 63282 7812
rect 240318 7800 240324 7812
rect 63276 7772 240324 7800
rect 63276 7760 63282 7772
rect 240318 7760 240324 7772
rect 240376 7760 240382 7812
rect 277578 7760 277584 7812
rect 277636 7800 277642 7812
rect 518342 7800 518348 7812
rect 277636 7772 518348 7800
rect 277636 7760 277642 7772
rect 518342 7760 518348 7772
rect 518400 7760 518406 7812
rect 59630 7692 59636 7744
rect 59688 7732 59694 7744
rect 239030 7732 239036 7744
rect 59688 7704 239036 7732
rect 59688 7692 59694 7704
rect 239030 7692 239036 7704
rect 239088 7692 239094 7744
rect 279694 7692 279700 7744
rect 279752 7732 279758 7744
rect 521838 7732 521844 7744
rect 279752 7704 521844 7732
rect 279752 7692 279758 7704
rect 521838 7692 521844 7704
rect 521896 7692 521902 7744
rect 21818 7624 21824 7676
rect 21876 7664 21882 7676
rect 235350 7664 235356 7676
rect 21876 7636 235356 7664
rect 21876 7624 21882 7636
rect 235350 7624 235356 7636
rect 235408 7624 235414 7676
rect 279786 7624 279792 7676
rect 279844 7664 279850 7676
rect 525426 7664 525432 7676
rect 279844 7636 525432 7664
rect 279844 7624 279850 7636
rect 525426 7624 525432 7636
rect 525484 7624 525490 7676
rect 13538 7556 13544 7608
rect 13596 7596 13602 7608
rect 235258 7596 235264 7608
rect 13596 7568 235264 7596
rect 13596 7556 13602 7568
rect 235258 7556 235264 7568
rect 235316 7556 235322 7608
rect 278774 7556 278780 7608
rect 278832 7596 278838 7608
rect 529014 7596 529020 7608
rect 278832 7568 529020 7596
rect 278832 7556 278838 7568
rect 529014 7556 529020 7568
rect 529072 7556 529078 7608
rect 105722 7488 105728 7540
rect 105780 7528 105786 7540
rect 234154 7528 234160 7540
rect 105780 7500 234160 7528
rect 105780 7488 105786 7500
rect 234154 7488 234160 7500
rect 234212 7488 234218 7540
rect 276750 7488 276756 7540
rect 276808 7528 276814 7540
rect 489914 7528 489920 7540
rect 276808 7500 489920 7528
rect 276808 7488 276814 7500
rect 489914 7488 489920 7500
rect 489972 7488 489978 7540
rect 116394 7420 116400 7472
rect 116452 7460 116458 7472
rect 244642 7460 244648 7472
rect 116452 7432 244648 7460
rect 116452 7420 116458 7432
rect 244642 7420 244648 7432
rect 244700 7420 244706 7472
rect 276934 7420 276940 7472
rect 276992 7460 276998 7472
rect 486418 7460 486424 7472
rect 276992 7432 486424 7460
rect 276992 7420 276998 7432
rect 486418 7420 486424 7432
rect 486476 7420 486482 7472
rect 112806 7352 112812 7404
rect 112864 7392 112870 7404
rect 234246 7392 234252 7404
rect 112864 7364 234252 7392
rect 112864 7352 112870 7364
rect 234246 7352 234252 7364
rect 234304 7352 234310 7404
rect 275094 7352 275100 7404
rect 275152 7392 275158 7404
rect 482830 7392 482836 7404
rect 275152 7364 482836 7392
rect 275152 7352 275158 7364
rect 482830 7352 482836 7364
rect 482888 7352 482894 7404
rect 119890 7284 119896 7336
rect 119948 7324 119954 7336
rect 234062 7324 234068 7336
rect 119948 7296 234068 7324
rect 119948 7284 119954 7296
rect 234062 7284 234068 7296
rect 234120 7284 234126 7336
rect 275186 7284 275192 7336
rect 275244 7324 275250 7336
rect 478138 7324 478144 7336
rect 275244 7296 478144 7324
rect 275244 7284 275250 7296
rect 478138 7284 478144 7296
rect 478196 7284 478202 7336
rect 275738 7216 275744 7268
rect 275796 7256 275802 7268
rect 474550 7256 474556 7268
rect 275796 7228 474556 7256
rect 275796 7216 275802 7228
rect 474550 7216 474556 7228
rect 474608 7216 474614 7268
rect 274358 7148 274364 7200
rect 274416 7188 274422 7200
rect 467466 7188 467472 7200
rect 274416 7160 467472 7188
rect 274416 7148 274422 7160
rect 467466 7148 467472 7160
rect 467524 7148 467530 7200
rect 273622 7080 273628 7132
rect 273680 7120 273686 7132
rect 463970 7120 463976 7132
rect 273680 7092 463976 7120
rect 273680 7080 273686 7092
rect 463970 7080 463976 7092
rect 464028 7080 464034 7132
rect 273714 7012 273720 7064
rect 273772 7052 273778 7064
rect 460382 7052 460388 7064
rect 273772 7024 460388 7052
rect 273772 7012 273778 7024
rect 460382 7012 460388 7024
rect 460440 7012 460446 7064
rect 270494 6944 270500 6996
rect 270552 6984 270558 6996
rect 432046 6984 432052 6996
rect 270552 6956 432052 6984
rect 270552 6944 270558 6956
rect 432046 6944 432052 6956
rect 432104 6944 432110 6996
rect 160094 6808 160100 6860
rect 160152 6848 160158 6860
rect 249058 6848 249064 6860
rect 160152 6820 249064 6848
rect 160152 6808 160158 6820
rect 249058 6808 249064 6820
rect 249116 6808 249122 6860
rect 260374 6808 260380 6860
rect 260432 6848 260438 6860
rect 294874 6848 294880 6860
rect 260432 6820 294880 6848
rect 260432 6808 260438 6820
rect 294874 6808 294880 6820
rect 294932 6808 294938 6860
rect 295978 6808 295984 6860
rect 296036 6848 296042 6860
rect 580166 6848 580172 6860
rect 296036 6820 580172 6848
rect 296036 6808 296042 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 156598 6740 156604 6792
rect 156656 6780 156662 6792
rect 247310 6780 247316 6792
rect 156656 6752 247316 6780
rect 156656 6740 156662 6752
rect 247310 6740 247316 6752
rect 247368 6740 247374 6792
rect 264606 6740 264612 6792
rect 264664 6780 264670 6792
rect 354030 6780 354036 6792
rect 264664 6752 354036 6780
rect 264664 6740 264670 6752
rect 354030 6740 354036 6752
rect 354088 6740 354094 6792
rect 153010 6672 153016 6724
rect 153068 6712 153074 6724
rect 247218 6712 247224 6724
rect 153068 6684 247224 6712
rect 153068 6672 153074 6684
rect 247218 6672 247224 6684
rect 247276 6672 247282 6724
rect 265526 6672 265532 6724
rect 265584 6712 265590 6724
rect 357526 6712 357532 6724
rect 265584 6684 357532 6712
rect 265584 6672 265590 6684
rect 357526 6672 357532 6684
rect 357584 6672 357590 6724
rect 149514 6604 149520 6656
rect 149572 6644 149578 6656
rect 247770 6644 247776 6656
rect 149572 6616 247776 6644
rect 149572 6604 149578 6616
rect 247770 6604 247776 6616
rect 247828 6604 247834 6656
rect 265710 6604 265716 6656
rect 265768 6644 265774 6656
rect 361114 6644 361120 6656
rect 265768 6616 361120 6644
rect 265768 6604 265774 6616
rect 361114 6604 361120 6616
rect 361172 6604 361178 6656
rect 145926 6536 145932 6588
rect 145984 6576 145990 6588
rect 247586 6576 247592 6588
rect 145984 6548 247592 6576
rect 145984 6536 145990 6548
rect 247586 6536 247592 6548
rect 247644 6536 247650 6588
rect 265986 6536 265992 6588
rect 266044 6576 266050 6588
rect 364610 6576 364616 6588
rect 266044 6548 364616 6576
rect 266044 6536 266050 6548
rect 364610 6536 364616 6548
rect 364668 6536 364674 6588
rect 2774 6468 2780 6520
rect 2832 6508 2838 6520
rect 4798 6508 4804 6520
rect 2832 6480 4804 6508
rect 2832 6468 2838 6480
rect 4798 6468 4804 6480
rect 4856 6468 4862 6520
rect 142430 6468 142436 6520
rect 142488 6508 142494 6520
rect 246022 6508 246028 6520
rect 142488 6480 246028 6508
rect 142488 6468 142494 6480
rect 246022 6468 246028 6480
rect 246080 6468 246086 6520
rect 266078 6468 266084 6520
rect 266136 6508 266142 6520
rect 368198 6508 368204 6520
rect 266136 6480 368204 6508
rect 266136 6468 266142 6480
rect 368198 6468 368204 6480
rect 368256 6468 368262 6520
rect 138842 6400 138848 6452
rect 138900 6440 138906 6452
rect 246206 6440 246212 6452
rect 138900 6412 246212 6440
rect 138900 6400 138906 6412
rect 246206 6400 246212 6412
rect 246264 6400 246270 6452
rect 266722 6400 266728 6452
rect 266780 6440 266786 6452
rect 374086 6440 374092 6452
rect 266780 6412 374092 6440
rect 266780 6400 266786 6412
rect 374086 6400 374092 6412
rect 374144 6400 374150 6452
rect 135254 6332 135260 6384
rect 135312 6372 135318 6384
rect 246114 6372 246120 6384
rect 135312 6344 246120 6372
rect 135312 6332 135318 6344
rect 246114 6332 246120 6344
rect 246172 6332 246178 6384
rect 266630 6332 266636 6384
rect 266688 6372 266694 6384
rect 377674 6372 377680 6384
rect 266688 6344 377680 6372
rect 266688 6332 266694 6344
rect 377674 6332 377680 6344
rect 377732 6332 377738 6384
rect 122282 6264 122288 6316
rect 122340 6304 122346 6316
rect 244458 6304 244464 6316
rect 122340 6276 244464 6304
rect 122340 6264 122346 6276
rect 244458 6264 244464 6276
rect 244516 6264 244522 6316
rect 267734 6264 267740 6316
rect 267792 6304 267798 6316
rect 393038 6304 393044 6316
rect 267792 6276 393044 6304
rect 267792 6264 267798 6276
rect 393038 6264 393044 6276
rect 393096 6264 393102 6316
rect 118786 6196 118792 6248
rect 118844 6236 118850 6248
rect 244550 6236 244556 6248
rect 118844 6208 244556 6236
rect 118844 6196 118850 6208
rect 244550 6196 244556 6208
rect 244608 6196 244614 6248
rect 267918 6196 267924 6248
rect 267976 6236 267982 6248
rect 396534 6236 396540 6248
rect 267976 6208 396540 6236
rect 267976 6196 267982 6208
rect 396534 6196 396540 6208
rect 396592 6196 396598 6248
rect 44266 6128 44272 6180
rect 44324 6168 44330 6180
rect 238110 6168 238116 6180
rect 44324 6140 238116 6168
rect 44324 6128 44330 6140
rect 238110 6128 238116 6140
rect 238168 6128 238174 6180
rect 268838 6128 268844 6180
rect 268896 6168 268902 6180
rect 400122 6168 400128 6180
rect 268896 6140 400128 6168
rect 268896 6128 268902 6140
rect 400122 6128 400128 6140
rect 400180 6128 400186 6180
rect 188522 6060 188528 6112
rect 188580 6100 188586 6112
rect 250254 6100 250260 6112
rect 188580 6072 250260 6100
rect 188580 6060 188586 6072
rect 250254 6060 250260 6072
rect 250312 6060 250318 6112
rect 264422 6060 264428 6112
rect 264480 6100 264486 6112
rect 350442 6100 350448 6112
rect 264480 6072 350448 6100
rect 264480 6060 264486 6072
rect 350442 6060 350448 6072
rect 350500 6060 350506 6112
rect 192018 5992 192024 6044
rect 192076 6032 192082 6044
rect 250346 6032 250352 6044
rect 192076 6004 250352 6032
rect 192076 5992 192082 6004
rect 250346 5992 250352 6004
rect 250404 5992 250410 6044
rect 264698 5992 264704 6044
rect 264756 6032 264762 6044
rect 346946 6032 346952 6044
rect 264756 6004 346952 6032
rect 264756 5992 264762 6004
rect 346946 5992 346952 6004
rect 347004 5992 347010 6044
rect 206186 5924 206192 5976
rect 206244 5964 206250 5976
rect 251542 5964 251548 5976
rect 206244 5936 251548 5964
rect 206244 5924 206250 5936
rect 251542 5924 251548 5936
rect 251600 5924 251606 5976
rect 264514 5924 264520 5976
rect 264572 5964 264578 5976
rect 343358 5964 343364 5976
rect 264572 5936 343364 5964
rect 264572 5924 264578 5936
rect 343358 5924 343364 5936
rect 343416 5924 343422 5976
rect 213362 5856 213368 5908
rect 213420 5896 213426 5908
rect 252922 5896 252928 5908
rect 213420 5868 252928 5896
rect 213420 5856 213426 5868
rect 252922 5856 252928 5868
rect 252980 5856 252986 5908
rect 263410 5856 263416 5908
rect 263468 5896 263474 5908
rect 338666 5896 338672 5908
rect 263468 5868 338672 5896
rect 263468 5856 263474 5868
rect 338666 5856 338672 5868
rect 338724 5856 338730 5908
rect 216858 5788 216864 5840
rect 216916 5828 216922 5840
rect 252830 5828 252836 5840
rect 216916 5800 252836 5828
rect 216916 5788 216922 5800
rect 252830 5788 252836 5800
rect 252888 5788 252894 5840
rect 263318 5788 263324 5840
rect 263376 5828 263382 5840
rect 335078 5828 335084 5840
rect 263376 5800 335084 5828
rect 263376 5788 263382 5800
rect 335078 5788 335084 5800
rect 335136 5788 335142 5840
rect 220446 5720 220452 5772
rect 220504 5760 220510 5772
rect 252738 5760 252744 5772
rect 220504 5732 252744 5760
rect 220504 5720 220510 5732
rect 252738 5720 252744 5732
rect 252796 5720 252802 5772
rect 262582 5720 262588 5772
rect 262640 5760 262646 5772
rect 331582 5760 331588 5772
rect 262640 5732 331588 5760
rect 262640 5720 262646 5732
rect 331582 5720 331588 5732
rect 331640 5720 331646 5772
rect 223942 5652 223948 5704
rect 224000 5692 224006 5704
rect 253658 5692 253664 5704
rect 224000 5664 253664 5692
rect 224000 5652 224006 5664
rect 253658 5652 253664 5664
rect 253716 5652 253722 5704
rect 263134 5652 263140 5704
rect 263192 5692 263198 5704
rect 327994 5692 328000 5704
rect 263192 5664 328000 5692
rect 263192 5652 263198 5664
rect 327994 5652 328000 5664
rect 328052 5652 328058 5704
rect 227530 5584 227536 5636
rect 227588 5624 227594 5636
rect 254302 5624 254308 5636
rect 227588 5596 254308 5624
rect 227588 5584 227594 5596
rect 254302 5584 254308 5596
rect 254360 5584 254366 5636
rect 262306 5584 262312 5636
rect 262364 5624 262370 5636
rect 324406 5624 324412 5636
rect 262364 5596 324412 5624
rect 262364 5584 262370 5596
rect 324406 5584 324412 5596
rect 324464 5584 324470 5636
rect 231026 5516 231032 5568
rect 231084 5556 231090 5568
rect 254210 5556 254216 5568
rect 231084 5528 254216 5556
rect 231084 5516 231090 5528
rect 254210 5516 254216 5528
rect 254268 5516 254274 5568
rect 260834 5516 260840 5568
rect 260892 5556 260898 5568
rect 322106 5556 322112 5568
rect 260892 5528 322112 5556
rect 260892 5516 260898 5528
rect 322106 5516 322112 5528
rect 322164 5516 322170 5568
rect 177942 5448 177948 5500
rect 178000 5488 178006 5500
rect 249978 5488 249984 5500
rect 178000 5460 249984 5488
rect 178000 5448 178006 5460
rect 249978 5448 249984 5460
rect 250036 5448 250042 5500
rect 259822 5448 259828 5500
rect 259880 5488 259886 5500
rect 290182 5488 290188 5500
rect 259880 5460 290188 5488
rect 259880 5448 259886 5460
rect 290182 5448 290188 5460
rect 290240 5448 290246 5500
rect 293126 5488 293132 5500
rect 290476 5460 293132 5488
rect 174262 5380 174268 5432
rect 174320 5420 174326 5432
rect 248690 5420 248696 5432
rect 174320 5392 248696 5420
rect 174320 5380 174326 5392
rect 248690 5380 248696 5392
rect 248748 5380 248754 5432
rect 260466 5380 260472 5432
rect 260524 5420 260530 5432
rect 290476 5420 290504 5460
rect 293126 5448 293132 5460
rect 293184 5448 293190 5500
rect 293218 5448 293224 5500
rect 293276 5488 293282 5500
rect 298281 5491 298339 5497
rect 293276 5460 298232 5488
rect 293276 5448 293282 5460
rect 260524 5392 290504 5420
rect 260524 5380 260530 5392
rect 290550 5380 290556 5432
rect 290608 5420 290614 5432
rect 298097 5423 298155 5429
rect 298097 5420 298109 5423
rect 290608 5392 298109 5420
rect 290608 5380 290614 5392
rect 298097 5389 298109 5392
rect 298143 5389 298155 5423
rect 298204 5420 298232 5460
rect 298281 5457 298293 5491
rect 298327 5488 298339 5491
rect 465166 5488 465172 5500
rect 298327 5460 465172 5488
rect 298327 5457 298339 5460
rect 298281 5451 298339 5457
rect 465166 5448 465172 5460
rect 465224 5448 465230 5500
rect 475746 5420 475752 5432
rect 298204 5392 475752 5420
rect 298097 5383 298155 5389
rect 475746 5380 475752 5392
rect 475804 5380 475810 5432
rect 173158 5312 173164 5364
rect 173216 5352 173222 5364
rect 249610 5352 249616 5364
rect 173216 5324 249616 5352
rect 173216 5312 173222 5324
rect 249610 5312 249616 5324
rect 249668 5312 249674 5364
rect 257338 5312 257344 5364
rect 257396 5352 257402 5364
rect 264146 5352 264152 5364
rect 257396 5324 264152 5352
rect 257396 5312 257402 5324
rect 264146 5312 264152 5324
rect 264204 5312 264210 5364
rect 277210 5312 277216 5364
rect 277268 5352 277274 5364
rect 492306 5352 492312 5364
rect 277268 5324 492312 5352
rect 277268 5312 277274 5324
rect 492306 5312 492312 5324
rect 492364 5312 492370 5364
rect 170766 5244 170772 5296
rect 170824 5284 170830 5296
rect 248782 5284 248788 5296
rect 170824 5256 248788 5284
rect 170824 5244 170830 5256
rect 248782 5244 248788 5256
rect 248840 5244 248846 5296
rect 257614 5244 257620 5296
rect 257672 5284 257678 5296
rect 267734 5284 267740 5296
rect 257672 5256 267740 5284
rect 257672 5244 257678 5256
rect 267734 5244 267740 5256
rect 267792 5244 267798 5296
rect 276106 5244 276112 5296
rect 276164 5284 276170 5296
rect 495894 5284 495900 5296
rect 276164 5256 495900 5284
rect 276164 5244 276170 5256
rect 495894 5244 495900 5256
rect 495952 5244 495958 5296
rect 169662 5176 169668 5228
rect 169720 5216 169726 5228
rect 248966 5216 248972 5228
rect 169720 5188 248972 5216
rect 169720 5176 169726 5188
rect 248966 5176 248972 5188
rect 249024 5176 249030 5228
rect 257522 5176 257528 5228
rect 257580 5216 257586 5228
rect 268838 5216 268844 5228
rect 257580 5188 268844 5216
rect 257580 5176 257586 5188
rect 268838 5176 268844 5188
rect 268896 5176 268902 5228
rect 277118 5176 277124 5228
rect 277176 5216 277182 5228
rect 499390 5216 499396 5228
rect 277176 5188 499396 5216
rect 277176 5176 277182 5188
rect 499390 5176 499396 5188
rect 499448 5176 499454 5228
rect 167178 5108 167184 5160
rect 167236 5148 167242 5160
rect 248874 5148 248880 5160
rect 167236 5120 248880 5148
rect 167236 5108 167242 5120
rect 248874 5108 248880 5120
rect 248932 5108 248938 5160
rect 257430 5108 257436 5160
rect 257488 5148 257494 5160
rect 271230 5148 271236 5160
rect 257488 5120 271236 5148
rect 257488 5108 257494 5120
rect 271230 5108 271236 5120
rect 271288 5108 271294 5160
rect 277762 5108 277768 5160
rect 277820 5148 277826 5160
rect 510062 5148 510068 5160
rect 277820 5120 510068 5148
rect 277820 5108 277826 5120
rect 510062 5108 510068 5120
rect 510120 5108 510126 5160
rect 166074 5040 166080 5092
rect 166132 5080 166138 5092
rect 248598 5080 248604 5092
rect 166132 5052 248604 5080
rect 166132 5040 166138 5052
rect 248598 5040 248604 5052
rect 248656 5040 248662 5092
rect 257706 5040 257712 5092
rect 257764 5080 257770 5092
rect 272426 5080 272432 5092
rect 257764 5052 272432 5080
rect 257764 5040 257770 5052
rect 272426 5040 272432 5052
rect 272484 5040 272490 5092
rect 278958 5040 278964 5092
rect 279016 5080 279022 5092
rect 282273 5083 282331 5089
rect 279016 5052 282224 5080
rect 279016 5040 279022 5052
rect 163682 4972 163688 5024
rect 163740 5012 163746 5024
rect 249426 5012 249432 5024
rect 163740 4984 249432 5012
rect 163740 4972 163746 4984
rect 249426 4972 249432 4984
rect 249484 4972 249490 5024
rect 259086 4972 259092 5024
rect 259144 5012 259150 5024
rect 276014 5012 276020 5024
rect 259144 4984 276020 5012
rect 259144 4972 259150 4984
rect 276014 4972 276020 4984
rect 276072 4972 276078 5024
rect 277394 4972 277400 5024
rect 277452 5012 277458 5024
rect 277452 4984 278452 5012
rect 277452 4972 277458 4984
rect 141234 4904 141240 4956
rect 141292 4944 141298 4956
rect 245930 4944 245936 4956
rect 141292 4916 245936 4944
rect 141292 4904 141298 4916
rect 245930 4904 245936 4916
rect 245988 4904 245994 4956
rect 246390 4904 246396 4956
rect 246448 4944 246454 4956
rect 255682 4944 255688 4956
rect 246448 4916 255688 4944
rect 246448 4904 246454 4916
rect 255682 4904 255688 4916
rect 255740 4904 255746 4956
rect 258902 4904 258908 4956
rect 258960 4944 258966 4956
rect 278314 4944 278320 4956
rect 258960 4916 278320 4944
rect 258960 4904 258966 4916
rect 278314 4904 278320 4916
rect 278372 4904 278378 4956
rect 278424 4944 278452 4984
rect 278498 4972 278504 5024
rect 278556 5012 278562 5024
rect 282089 5015 282147 5021
rect 282089 5012 282101 5015
rect 278556 4984 282101 5012
rect 278556 4972 278562 4984
rect 282089 4981 282101 4984
rect 282135 4981 282147 5015
rect 282089 4975 282147 4981
rect 278424 4916 279648 4944
rect 12342 4836 12348 4888
rect 12400 4876 12406 4888
rect 235626 4876 235632 4888
rect 12400 4848 235632 4876
rect 12400 4836 12406 4848
rect 235626 4836 235632 4848
rect 235684 4836 235690 4888
rect 242894 4836 242900 4888
rect 242952 4876 242958 4888
rect 255774 4876 255780 4888
rect 242952 4848 255780 4876
rect 242952 4836 242958 4848
rect 255774 4836 255780 4848
rect 255832 4836 255838 4888
rect 259178 4836 259184 4888
rect 259236 4876 259242 4888
rect 279510 4876 279516 4888
rect 259236 4848 279516 4876
rect 259236 4836 259242 4848
rect 279510 4836 279516 4848
rect 279568 4836 279574 4888
rect 279620 4876 279648 4916
rect 280246 4904 280252 4956
rect 280304 4944 280310 4956
rect 282196 4944 282224 5052
rect 282273 5049 282285 5083
rect 282319 5080 282331 5083
rect 513558 5080 513564 5092
rect 282319 5052 513564 5080
rect 282319 5049 282331 5052
rect 282273 5043 282331 5049
rect 513558 5040 513564 5052
rect 513616 5040 513622 5092
rect 282365 5015 282423 5021
rect 282365 4981 282377 5015
rect 282411 5012 282423 5015
rect 517146 5012 517152 5024
rect 282411 4984 517152 5012
rect 282411 4981 282423 4984
rect 282365 4975 282423 4981
rect 517146 4972 517152 4984
rect 517204 4972 517210 5024
rect 534902 4944 534908 4956
rect 280304 4916 282132 4944
rect 282196 4916 534908 4944
rect 280304 4904 280310 4916
rect 281721 4879 281779 4885
rect 281721 4876 281733 4879
rect 279620 4848 281733 4876
rect 281721 4845 281733 4848
rect 281767 4845 281779 4879
rect 281721 4839 281779 4845
rect 281810 4836 281816 4888
rect 281868 4876 281874 4888
rect 282104 4876 282132 4916
rect 534902 4904 534908 4916
rect 534960 4904 534966 4956
rect 545482 4876 545488 4888
rect 281868 4848 282040 4876
rect 282104 4848 545488 4876
rect 281868 4836 281874 4848
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 234430 4808 234436 4820
rect 7708 4780 234436 4808
rect 7708 4768 7714 4780
rect 234430 4768 234436 4780
rect 234488 4768 234494 4820
rect 234614 4768 234620 4820
rect 234672 4808 234678 4820
rect 254118 4808 254124 4820
rect 234672 4780 254124 4808
rect 234672 4768 234678 4780
rect 254118 4768 254124 4780
rect 254176 4768 254182 4820
rect 258350 4768 258356 4820
rect 258408 4808 258414 4820
rect 281902 4808 281908 4820
rect 258408 4780 281908 4808
rect 258408 4768 258414 4780
rect 281902 4768 281908 4780
rect 281960 4768 281966 4820
rect 282012 4808 282040 4848
rect 545482 4836 545488 4848
rect 545540 4836 545546 4888
rect 556154 4808 556160 4820
rect 282012 4780 556160 4808
rect 556154 4768 556160 4780
rect 556212 4768 556218 4820
rect 181438 4700 181444 4752
rect 181496 4740 181502 4752
rect 250622 4740 250628 4752
rect 181496 4712 250628 4740
rect 181496 4700 181502 4712
rect 250622 4700 250628 4712
rect 250680 4700 250686 4752
rect 258994 4700 259000 4752
rect 259052 4740 259058 4752
rect 283098 4740 283104 4752
rect 259052 4712 283104 4740
rect 259052 4700 259058 4712
rect 283098 4700 283104 4712
rect 283156 4700 283162 4752
rect 291930 4700 291936 4752
rect 291988 4740 291994 4752
rect 293037 4743 293095 4749
rect 293037 4740 293049 4743
rect 291988 4712 293049 4740
rect 291988 4700 291994 4712
rect 293037 4709 293049 4712
rect 293083 4709 293095 4743
rect 293037 4703 293095 4709
rect 293126 4700 293132 4752
rect 293184 4740 293190 4752
rect 293678 4740 293684 4752
rect 293184 4712 293684 4740
rect 293184 4700 293190 4712
rect 293678 4700 293684 4712
rect 293736 4700 293742 4752
rect 293773 4743 293831 4749
rect 293773 4709 293785 4743
rect 293819 4740 293831 4743
rect 458082 4740 458088 4752
rect 293819 4712 458088 4740
rect 293819 4709 293831 4712
rect 293773 4703 293831 4709
rect 458082 4700 458088 4712
rect 458140 4700 458146 4752
rect 184934 4632 184940 4684
rect 184992 4672 184998 4684
rect 250714 4672 250720 4684
rect 184992 4644 250720 4672
rect 184992 4632 184998 4644
rect 250714 4632 250720 4644
rect 250772 4632 250778 4684
rect 264790 4632 264796 4684
rect 264848 4672 264854 4684
rect 352834 4672 352840 4684
rect 264848 4644 352840 4672
rect 264848 4632 264854 4644
rect 352834 4632 352840 4644
rect 352892 4632 352898 4684
rect 187326 4564 187332 4616
rect 187384 4604 187390 4616
rect 250162 4604 250168 4616
rect 187384 4576 250168 4604
rect 187384 4564 187390 4576
rect 250162 4564 250168 4576
rect 250220 4564 250226 4616
rect 263778 4564 263784 4616
rect 263836 4604 263842 4616
rect 339862 4604 339868 4616
rect 263836 4576 339868 4604
rect 263836 4564 263842 4576
rect 339862 4564 339868 4576
rect 339920 4564 339926 4616
rect 190822 4496 190828 4548
rect 190880 4536 190886 4548
rect 250070 4536 250076 4548
rect 190880 4508 250076 4536
rect 190880 4496 190886 4508
rect 250070 4496 250076 4508
rect 250128 4496 250134 4548
rect 261938 4496 261944 4548
rect 261996 4536 262002 4548
rect 318518 4536 318524 4548
rect 261996 4508 318524 4536
rect 261996 4496 262002 4508
rect 318518 4496 318524 4508
rect 318576 4496 318582 4548
rect 194410 4428 194416 4480
rect 194468 4468 194474 4480
rect 251450 4468 251456 4480
rect 194468 4440 251456 4468
rect 194468 4428 194474 4440
rect 251450 4428 251456 4440
rect 251508 4428 251514 4480
rect 261110 4428 261116 4480
rect 261168 4468 261174 4480
rect 315022 4468 315028 4480
rect 261168 4440 315028 4468
rect 261168 4428 261174 4440
rect 315022 4428 315028 4440
rect 315080 4428 315086 4480
rect 197906 4360 197912 4412
rect 197964 4400 197970 4412
rect 252278 4400 252284 4412
rect 197964 4372 252284 4400
rect 197964 4360 197970 4372
rect 252278 4360 252284 4372
rect 252336 4360 252342 4412
rect 261570 4360 261576 4412
rect 261628 4400 261634 4412
rect 311434 4400 311440 4412
rect 261628 4372 311440 4400
rect 261628 4360 261634 4372
rect 311434 4360 311440 4372
rect 311492 4360 311498 4412
rect 201494 4292 201500 4344
rect 201552 4332 201558 4344
rect 251358 4332 251364 4344
rect 201552 4304 251364 4332
rect 201552 4292 201558 4304
rect 251358 4292 251364 4304
rect 251416 4292 251422 4344
rect 259638 4292 259644 4344
rect 259696 4332 259702 4344
rect 304350 4332 304356 4344
rect 259696 4304 304356 4332
rect 259696 4292 259702 4304
rect 304350 4292 304356 4304
rect 304408 4292 304414 4344
rect 205082 4224 205088 4276
rect 205140 4264 205146 4276
rect 252186 4264 252192 4276
rect 205140 4236 252192 4264
rect 205140 4224 205146 4236
rect 252186 4224 252192 4236
rect 252244 4224 252250 4276
rect 259454 4224 259460 4276
rect 259512 4264 259518 4276
rect 300762 4264 300768 4276
rect 259512 4236 300768 4264
rect 259512 4224 259518 4236
rect 300762 4224 300768 4236
rect 300820 4224 300826 4276
rect 218054 4156 218060 4208
rect 218112 4196 218118 4208
rect 219342 4196 219348 4208
rect 218112 4168 219348 4196
rect 218112 4156 218118 4168
rect 219342 4156 219348 4168
rect 219400 4156 219406 4208
rect 222746 4156 222752 4208
rect 222804 4196 222810 4208
rect 226242 4196 226248 4208
rect 222804 4168 226248 4196
rect 222804 4156 222810 4168
rect 226242 4156 226248 4168
rect 226300 4156 226306 4208
rect 226334 4156 226340 4208
rect 226392 4196 226398 4208
rect 227622 4196 227628 4208
rect 226392 4168 227628 4196
rect 226392 4156 226398 4168
rect 227622 4156 227628 4168
rect 227680 4156 227686 4208
rect 227714 4156 227720 4208
rect 227772 4196 227778 4208
rect 253382 4196 253388 4208
rect 227772 4168 253388 4196
rect 227772 4156 227778 4168
rect 253382 4156 253388 4168
rect 253440 4156 253446 4208
rect 260558 4156 260564 4208
rect 260616 4196 260622 4208
rect 297266 4196 297272 4208
rect 260616 4168 297272 4196
rect 260616 4156 260622 4168
rect 297266 4156 297272 4168
rect 297324 4156 297330 4208
rect 440234 4156 440240 4208
rect 440292 4196 440298 4208
rect 441522 4196 441528 4208
rect 440292 4168 441528 4196
rect 440292 4156 440298 4168
rect 441522 4156 441528 4168
rect 441580 4156 441586 4208
rect 57238 4088 57244 4140
rect 57296 4128 57302 4140
rect 57296 4100 64874 4128
rect 57296 4088 57302 4100
rect 60826 4020 60832 4072
rect 60884 4060 60890 4072
rect 61930 4060 61936 4072
rect 60884 4032 61936 4060
rect 60884 4020 60890 4032
rect 61930 4020 61936 4032
rect 61988 4020 61994 4072
rect 64846 4060 64874 4100
rect 69106 4088 69112 4140
rect 69164 4128 69170 4140
rect 70302 4128 70308 4140
rect 69164 4100 70308 4128
rect 69164 4088 69170 4100
rect 70302 4088 70308 4100
rect 70360 4088 70366 4140
rect 71498 4088 71504 4140
rect 71556 4128 71562 4140
rect 233881 4131 233939 4137
rect 233881 4128 233893 4131
rect 71556 4100 233893 4128
rect 71556 4088 71562 4100
rect 233881 4097 233893 4100
rect 233927 4097 233939 4131
rect 233881 4091 233939 4097
rect 234062 4088 234068 4140
rect 234120 4128 234126 4140
rect 238386 4128 238392 4140
rect 234120 4100 238392 4128
rect 234120 4088 234126 4100
rect 238386 4088 238392 4100
rect 238444 4088 238450 4140
rect 284846 4088 284852 4140
rect 284904 4128 284910 4140
rect 299658 4128 299664 4140
rect 284904 4100 299664 4128
rect 284904 4088 284910 4100
rect 299658 4088 299664 4100
rect 299716 4088 299722 4140
rect 300118 4088 300124 4140
rect 300176 4128 300182 4140
rect 433242 4128 433248 4140
rect 300176 4100 433248 4128
rect 300176 4088 300182 4100
rect 433242 4088 433248 4100
rect 433300 4088 433306 4140
rect 434162 4088 434168 4140
rect 434220 4128 434226 4140
rect 508866 4128 508872 4140
rect 434220 4100 508872 4128
rect 434220 4088 434226 4100
rect 508866 4088 508872 4100
rect 508924 4088 508930 4140
rect 239306 4060 239312 4072
rect 64846 4032 239312 4060
rect 239306 4020 239312 4032
rect 239364 4020 239370 4072
rect 290458 4020 290464 4072
rect 290516 4060 290522 4072
rect 422570 4060 422576 4072
rect 290516 4032 422576 4060
rect 290516 4020 290522 4032
rect 422570 4020 422576 4032
rect 422628 4020 422634 4072
rect 422938 4020 422944 4072
rect 422996 4060 423002 4072
rect 422996 4032 431954 4060
rect 422996 4020 423002 4032
rect 50154 3952 50160 4004
rect 50212 3992 50218 4004
rect 238018 3992 238024 4004
rect 50212 3964 238024 3992
rect 50212 3952 50218 3964
rect 238018 3952 238024 3964
rect 238076 3952 238082 4004
rect 289446 3952 289452 4004
rect 289504 3992 289510 4004
rect 296073 3995 296131 4001
rect 296073 3992 296085 3995
rect 289504 3964 296085 3992
rect 289504 3952 289510 3964
rect 296073 3961 296085 3964
rect 296119 3961 296131 3995
rect 296073 3955 296131 3961
rect 296162 3952 296168 4004
rect 296220 3992 296226 4004
rect 429654 3992 429660 4004
rect 296220 3964 429660 3992
rect 296220 3952 296226 3964
rect 429654 3952 429660 3964
rect 429712 3952 429718 4004
rect 431926 3992 431954 4032
rect 433978 4020 433984 4072
rect 434036 4060 434042 4072
rect 512454 4060 512460 4072
rect 434036 4032 512460 4060
rect 434036 4020 434042 4032
rect 512454 4020 512460 4032
rect 512512 4020 512518 4072
rect 439130 3992 439136 4004
rect 431926 3964 439136 3992
rect 439130 3952 439136 3964
rect 439188 3952 439194 4004
rect 439498 3952 439504 4004
rect 439556 3992 439562 4004
rect 519538 3992 519544 4004
rect 439556 3964 519544 3992
rect 439556 3952 439562 3964
rect 519538 3952 519544 3964
rect 519596 3952 519602 4004
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 238846 3924 238852 3936
rect 46716 3896 238852 3924
rect 46716 3884 46722 3896
rect 238846 3884 238852 3896
rect 238904 3884 238910 3936
rect 291838 3884 291844 3936
rect 291896 3924 291902 3936
rect 426158 3924 426164 3936
rect 291896 3896 426164 3924
rect 291896 3884 291902 3896
rect 426158 3884 426164 3896
rect 426216 3884 426222 3936
rect 434070 3884 434076 3936
rect 434128 3924 434134 3936
rect 515950 3924 515956 3936
rect 434128 3896 515956 3924
rect 434128 3884 434134 3896
rect 515950 3884 515956 3896
rect 516008 3884 516014 3936
rect 45462 3816 45468 3868
rect 45520 3856 45526 3868
rect 238202 3856 238208 3868
rect 45520 3828 238208 3856
rect 45520 3816 45526 3828
rect 238202 3816 238208 3828
rect 238260 3816 238266 3868
rect 269574 3816 269580 3868
rect 269632 3856 269638 3868
rect 408402 3856 408408 3868
rect 269632 3828 408408 3856
rect 269632 3816 269638 3828
rect 408402 3816 408408 3828
rect 408460 3816 408466 3868
rect 408494 3816 408500 3868
rect 408552 3856 408558 3868
rect 533706 3856 533712 3868
rect 408552 3828 533712 3856
rect 408552 3816 408558 3828
rect 533706 3816 533712 3828
rect 533764 3816 533770 3868
rect 39574 3748 39580 3800
rect 39632 3788 39638 3800
rect 237466 3788 237472 3800
rect 39632 3760 237472 3788
rect 39632 3748 39638 3760
rect 237466 3748 237472 3760
rect 237524 3748 237530 3800
rect 247586 3748 247592 3800
rect 247644 3788 247650 3800
rect 255498 3788 255504 3800
rect 247644 3760 255504 3788
rect 247644 3748 247650 3760
rect 255498 3748 255504 3760
rect 255556 3748 255562 3800
rect 289538 3748 289544 3800
rect 289596 3788 289602 3800
rect 447410 3788 447416 3800
rect 289596 3760 447416 3788
rect 289596 3748 289602 3760
rect 447410 3748 447416 3760
rect 447468 3748 447474 3800
rect 38378 3680 38384 3732
rect 38436 3720 38442 3732
rect 237650 3720 237656 3732
rect 38436 3692 237656 3720
rect 38436 3680 38442 3692
rect 237650 3680 237656 3692
rect 237708 3680 237714 3732
rect 239125 3723 239183 3729
rect 239125 3689 239137 3723
rect 239171 3720 239183 3723
rect 242710 3720 242716 3732
rect 239171 3692 242716 3720
rect 239171 3689 239183 3692
rect 239125 3683 239183 3689
rect 242710 3680 242716 3692
rect 242768 3680 242774 3732
rect 244090 3680 244096 3732
rect 244148 3720 244154 3732
rect 251910 3720 251916 3732
rect 244148 3692 251916 3720
rect 244148 3680 244154 3692
rect 251910 3680 251916 3692
rect 251968 3680 251974 3732
rect 280798 3680 280804 3732
rect 280856 3720 280862 3732
rect 443822 3720 443828 3732
rect 280856 3692 443828 3720
rect 280856 3680 280862 3692
rect 443822 3680 443828 3692
rect 443880 3680 443886 3732
rect 32398 3612 32404 3664
rect 32456 3652 32462 3664
rect 237558 3652 237564 3664
rect 32456 3624 237564 3652
rect 32456 3612 32462 3624
rect 237558 3612 237564 3624
rect 237616 3612 237622 3664
rect 241698 3612 241704 3664
rect 241756 3652 241762 3664
rect 252002 3652 252008 3664
rect 241756 3624 252008 3652
rect 241756 3612 241762 3624
rect 252002 3612 252008 3624
rect 252060 3612 252066 3664
rect 254670 3612 254676 3664
rect 254728 3612 254734 3664
rect 258534 3612 258540 3664
rect 258592 3652 258598 3664
rect 258592 3624 267734 3652
rect 258592 3612 258598 3624
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 28810 3584 28816 3596
rect 27764 3556 28816 3584
rect 27764 3544 27770 3556
rect 28810 3544 28816 3556
rect 28868 3544 28874 3596
rect 31294 3544 31300 3596
rect 31352 3584 31358 3596
rect 232038 3584 232044 3596
rect 31352 3556 232044 3584
rect 31352 3544 31358 3556
rect 232038 3544 232044 3556
rect 232096 3544 232102 3596
rect 236454 3584 236460 3596
rect 232148 3556 236460 3584
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 20622 3516 20628 3528
rect 19484 3488 20628 3516
rect 19484 3476 19490 3488
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 232148 3516 232176 3556
rect 236454 3544 236460 3556
rect 236512 3544 236518 3596
rect 238726 3556 239352 3584
rect 24268 3488 232176 3516
rect 24268 3476 24274 3488
rect 232222 3476 232228 3528
rect 232280 3516 232286 3528
rect 233142 3516 233148 3528
rect 232280 3488 233148 3516
rect 232280 3476 232286 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233418 3476 233424 3528
rect 233476 3516 233482 3528
rect 234522 3516 234528 3528
rect 233476 3488 234528 3516
rect 233476 3476 233482 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 238110 3476 238116 3528
rect 238168 3516 238174 3528
rect 238726 3516 238754 3556
rect 238168 3488 238754 3516
rect 238168 3476 238174 3488
rect 14734 3408 14740 3460
rect 14792 3448 14798 3460
rect 237098 3448 237104 3460
rect 14792 3420 237104 3448
rect 14792 3408 14798 3420
rect 237098 3408 237104 3420
rect 237156 3408 237162 3460
rect 239324 3448 239352 3556
rect 240502 3544 240508 3596
rect 240560 3584 240566 3596
rect 254688 3584 254716 3612
rect 240560 3556 254716 3584
rect 240560 3544 240566 3556
rect 257890 3544 257896 3596
rect 257948 3584 257954 3596
rect 260650 3584 260656 3596
rect 257948 3556 260656 3584
rect 257948 3544 257954 3556
rect 260650 3544 260656 3556
rect 260708 3544 260714 3596
rect 267706 3584 267734 3624
rect 290642 3612 290648 3664
rect 290700 3652 290706 3664
rect 296257 3655 296315 3661
rect 290700 3624 296208 3652
rect 290700 3612 290706 3624
rect 280706 3584 280712 3596
rect 267706 3556 280712 3584
rect 280706 3544 280712 3556
rect 280764 3544 280770 3596
rect 287698 3544 287704 3596
rect 287756 3584 287762 3596
rect 288986 3584 288992 3596
rect 287756 3556 288992 3584
rect 287756 3544 287762 3556
rect 288986 3544 288992 3556
rect 289044 3544 289050 3596
rect 289354 3544 289360 3596
rect 289412 3584 289418 3596
rect 296070 3584 296076 3596
rect 289412 3556 296076 3584
rect 289412 3544 289418 3556
rect 296070 3544 296076 3556
rect 296128 3544 296134 3596
rect 296180 3584 296208 3624
rect 296257 3621 296269 3655
rect 296303 3652 296315 3655
rect 454494 3652 454500 3664
rect 296303 3624 454500 3652
rect 296303 3621 296315 3624
rect 296257 3615 296315 3621
rect 454494 3612 454500 3624
rect 454552 3612 454558 3664
rect 461578 3584 461584 3596
rect 296180 3556 461584 3584
rect 461578 3544 461584 3556
rect 461636 3544 461642 3596
rect 244366 3476 244372 3528
rect 244424 3516 244430 3528
rect 245194 3516 245200 3528
rect 244424 3488 245200 3516
rect 244424 3476 244430 3488
rect 245194 3476 245200 3488
rect 245252 3476 245258 3528
rect 254670 3476 254676 3528
rect 254728 3516 254734 3528
rect 255406 3516 255412 3528
rect 254728 3488 255412 3516
rect 254728 3476 254734 3488
rect 255406 3476 255412 3488
rect 255464 3476 255470 3528
rect 257798 3476 257804 3528
rect 257856 3516 257862 3528
rect 259454 3516 259460 3528
rect 257856 3488 259460 3516
rect 257856 3476 257862 3488
rect 259454 3476 259460 3488
rect 259512 3476 259518 3528
rect 260098 3476 260104 3528
rect 260156 3516 260162 3528
rect 261754 3516 261760 3528
rect 260156 3488 261760 3516
rect 260156 3476 260162 3488
rect 261754 3476 261760 3488
rect 261812 3476 261818 3528
rect 276658 3476 276664 3528
rect 276716 3516 276722 3528
rect 468662 3516 468668 3528
rect 276716 3488 468668 3516
rect 276716 3476 276722 3488
rect 468662 3476 468668 3488
rect 468720 3476 468726 3528
rect 254854 3448 254860 3460
rect 239324 3420 254860 3448
rect 254854 3408 254860 3420
rect 254912 3408 254918 3460
rect 257154 3408 257160 3460
rect 257212 3448 257218 3460
rect 265342 3448 265348 3460
rect 257212 3420 265348 3448
rect 257212 3408 257218 3420
rect 265342 3408 265348 3420
rect 265400 3408 265406 3460
rect 271138 3408 271144 3460
rect 271196 3448 271202 3460
rect 316218 3448 316224 3460
rect 271196 3420 316224 3448
rect 271196 3408 271202 3420
rect 316218 3408 316224 3420
rect 316276 3408 316282 3460
rect 319438 3408 319444 3460
rect 319496 3448 319502 3460
rect 583386 3448 583392 3460
rect 319496 3420 583392 3448
rect 319496 3408 319502 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 35802 3380 35808 3392
rect 34848 3352 35808 3380
rect 34848 3340 34854 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 35986 3340 35992 3392
rect 36044 3380 36050 3392
rect 37182 3380 37188 3392
rect 36044 3352 37188 3380
rect 36044 3340 36050 3352
rect 37182 3340 37188 3352
rect 37240 3340 37246 3392
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 42702 3380 42708 3392
rect 41932 3352 42708 3380
rect 41932 3340 41938 3352
rect 42702 3340 42708 3352
rect 42760 3340 42766 3392
rect 43070 3340 43076 3392
rect 43128 3380 43134 3392
rect 44082 3380 44088 3392
rect 43128 3352 44088 3380
rect 43128 3340 43134 3352
rect 44082 3340 44088 3352
rect 44140 3340 44146 3392
rect 48958 3340 48964 3392
rect 49016 3380 49022 3392
rect 49602 3380 49608 3392
rect 49016 3352 49608 3380
rect 49016 3340 49022 3352
rect 49602 3340 49608 3352
rect 49660 3340 49666 3392
rect 51350 3340 51356 3392
rect 51408 3380 51414 3392
rect 52362 3380 52368 3392
rect 51408 3352 52368 3380
rect 51408 3340 51414 3352
rect 52362 3340 52368 3352
rect 52420 3340 52426 3392
rect 52546 3340 52552 3392
rect 52604 3380 52610 3392
rect 53650 3380 53656 3392
rect 52604 3352 53656 3380
rect 52604 3340 52610 3352
rect 53650 3340 53656 3352
rect 53708 3340 53714 3392
rect 58434 3340 58440 3392
rect 58492 3380 58498 3392
rect 59262 3380 59268 3392
rect 58492 3352 59268 3380
rect 58492 3340 58498 3352
rect 59262 3340 59268 3352
rect 59320 3340 59326 3392
rect 64322 3340 64328 3392
rect 64380 3380 64386 3392
rect 64782 3380 64788 3392
rect 64380 3352 64788 3380
rect 64380 3340 64386 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 65518 3340 65524 3392
rect 65576 3380 65582 3392
rect 66162 3380 66168 3392
rect 65576 3352 66168 3380
rect 65576 3340 65582 3352
rect 66162 3340 66168 3352
rect 66220 3340 66226 3392
rect 67910 3340 67916 3392
rect 67968 3380 67974 3392
rect 68922 3380 68928 3392
rect 67968 3352 68928 3380
rect 67968 3340 67974 3352
rect 68922 3340 68928 3352
rect 68980 3340 68986 3392
rect 72602 3340 72608 3392
rect 72660 3380 72666 3392
rect 73062 3380 73068 3392
rect 72660 3352 73068 3380
rect 72660 3340 72666 3352
rect 73062 3340 73068 3352
rect 73120 3340 73126 3392
rect 74994 3340 75000 3392
rect 75052 3380 75058 3392
rect 75822 3380 75828 3392
rect 75052 3352 75828 3380
rect 75052 3340 75058 3352
rect 75822 3340 75828 3352
rect 75880 3340 75886 3392
rect 76190 3340 76196 3392
rect 76248 3380 76254 3392
rect 77202 3380 77208 3392
rect 76248 3352 77208 3380
rect 76248 3340 76254 3352
rect 77202 3340 77208 3352
rect 77260 3340 77266 3392
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 81342 3380 81348 3392
rect 80940 3352 81348 3380
rect 80940 3340 80946 3352
rect 81342 3340 81348 3352
rect 81400 3340 81406 3392
rect 82078 3340 82084 3392
rect 82136 3380 82142 3392
rect 82722 3380 82728 3392
rect 82136 3352 82728 3380
rect 82136 3340 82142 3352
rect 82722 3340 82728 3352
rect 82780 3340 82786 3392
rect 83274 3340 83280 3392
rect 83332 3380 83338 3392
rect 84102 3380 84108 3392
rect 83332 3352 84108 3380
rect 83332 3340 83338 3352
rect 84102 3340 84108 3352
rect 84160 3340 84166 3392
rect 84470 3340 84476 3392
rect 84528 3380 84534 3392
rect 85482 3380 85488 3392
rect 84528 3352 85488 3380
rect 84528 3340 84534 3352
rect 85482 3340 85488 3352
rect 85540 3340 85546 3392
rect 85666 3340 85672 3392
rect 85724 3380 85730 3392
rect 86678 3380 86684 3392
rect 85724 3352 86684 3380
rect 85724 3340 85730 3352
rect 86678 3340 86684 3352
rect 86736 3340 86742 3392
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 92382 3380 92388 3392
rect 91612 3352 92388 3380
rect 91612 3340 91618 3352
rect 92382 3340 92388 3352
rect 92440 3340 92446 3392
rect 239125 3383 239183 3389
rect 239125 3380 239137 3383
rect 92492 3352 239137 3380
rect 6454 3272 6460 3324
rect 6512 3312 6518 3324
rect 7558 3312 7564 3324
rect 6512 3284 7564 3312
rect 6512 3272 6518 3284
rect 7558 3272 7564 3284
rect 7616 3272 7622 3324
rect 78582 3272 78588 3324
rect 78640 3312 78646 3324
rect 92492 3312 92520 3352
rect 239125 3349 239137 3352
rect 239171 3349 239183 3383
rect 242618 3380 242624 3392
rect 239125 3343 239183 3349
rect 239232 3352 242624 3380
rect 78640 3284 92520 3312
rect 78640 3272 78646 3284
rect 92750 3272 92756 3324
rect 92808 3312 92814 3324
rect 93762 3312 93768 3324
rect 92808 3284 93768 3312
rect 92808 3272 92814 3284
rect 93762 3272 93768 3284
rect 93820 3272 93826 3324
rect 97442 3272 97448 3324
rect 97500 3312 97506 3324
rect 97902 3312 97908 3324
rect 97500 3284 97908 3312
rect 97500 3272 97506 3284
rect 97902 3272 97908 3284
rect 97960 3272 97966 3324
rect 99834 3272 99840 3324
rect 99892 3312 99898 3324
rect 100662 3312 100668 3324
rect 99892 3284 100668 3312
rect 99892 3272 99898 3284
rect 100662 3272 100668 3284
rect 100720 3272 100726 3324
rect 101030 3272 101036 3324
rect 101088 3312 101094 3324
rect 102042 3312 102048 3324
rect 101088 3284 102048 3312
rect 101088 3272 101094 3284
rect 102042 3272 102048 3284
rect 102100 3272 102106 3324
rect 239232 3312 239260 3352
rect 242618 3340 242624 3352
rect 242676 3340 242682 3392
rect 251174 3340 251180 3392
rect 251232 3380 251238 3392
rect 256418 3380 256424 3392
rect 251232 3352 256424 3380
rect 251232 3340 251238 3352
rect 256418 3340 256424 3352
rect 256476 3340 256482 3392
rect 268194 3340 268200 3392
rect 268252 3380 268258 3392
rect 401318 3380 401324 3392
rect 268252 3352 401324 3380
rect 268252 3340 268258 3352
rect 401318 3340 401324 3352
rect 401376 3340 401382 3392
rect 403618 3340 403624 3392
rect 403676 3380 403682 3392
rect 526622 3380 526628 3392
rect 403676 3352 526628 3380
rect 403676 3340 403682 3352
rect 526622 3340 526628 3352
rect 526680 3340 526686 3392
rect 102152 3284 239260 3312
rect 89162 3204 89168 3256
rect 89220 3244 89226 3256
rect 102152 3244 102180 3284
rect 239306 3272 239312 3324
rect 239364 3312 239370 3324
rect 244918 3312 244924 3324
rect 239364 3284 244924 3312
rect 239364 3272 239370 3284
rect 244918 3272 244924 3284
rect 244976 3272 244982 3324
rect 264238 3272 264244 3324
rect 264296 3312 264302 3324
rect 270034 3312 270040 3324
rect 264296 3284 270040 3312
rect 264296 3272 264302 3284
rect 270034 3272 270040 3284
rect 270092 3272 270098 3324
rect 271506 3272 271512 3324
rect 271564 3312 271570 3324
rect 305546 3312 305552 3324
rect 271564 3284 305552 3312
rect 271564 3272 271570 3284
rect 305546 3272 305552 3284
rect 305604 3272 305610 3324
rect 307754 3272 307760 3324
rect 307812 3312 307818 3324
rect 309042 3312 309048 3324
rect 307812 3284 309048 3312
rect 307812 3272 307818 3284
rect 309042 3272 309048 3284
rect 309100 3272 309106 3324
rect 309134 3272 309140 3324
rect 309192 3312 309198 3324
rect 436738 3312 436744 3324
rect 309192 3284 436744 3312
rect 309192 3272 309198 3284
rect 436738 3272 436744 3284
rect 436796 3272 436802 3324
rect 439590 3272 439596 3324
rect 439648 3312 439654 3324
rect 448606 3312 448612 3324
rect 439648 3284 448612 3312
rect 439648 3272 439654 3284
rect 448606 3272 448612 3284
rect 448664 3272 448670 3324
rect 243906 3244 243912 3256
rect 89220 3216 102180 3244
rect 102244 3216 243912 3244
rect 89220 3204 89226 3216
rect 96246 3136 96252 3188
rect 96304 3176 96310 3188
rect 102244 3176 102272 3216
rect 243906 3204 243912 3216
rect 243964 3204 243970 3256
rect 280890 3204 280896 3256
rect 280948 3244 280954 3256
rect 394234 3244 394240 3256
rect 280948 3216 394240 3244
rect 280948 3204 280954 3216
rect 394234 3204 394240 3216
rect 394292 3204 394298 3256
rect 396718 3204 396724 3256
rect 396776 3244 396782 3256
rect 498194 3244 498200 3256
rect 396776 3216 498200 3244
rect 396776 3204 396782 3216
rect 498194 3204 498200 3216
rect 498252 3204 498258 3256
rect 96304 3148 102272 3176
rect 96304 3136 96310 3148
rect 103330 3136 103336 3188
rect 103388 3176 103394 3188
rect 243446 3176 243452 3188
rect 103388 3148 243452 3176
rect 103388 3136 103394 3148
rect 243446 3136 243452 3148
rect 243504 3136 243510 3188
rect 271414 3136 271420 3188
rect 271472 3176 271478 3188
rect 273622 3176 273628 3188
rect 271472 3148 273628 3176
rect 271472 3136 271478 3148
rect 273622 3136 273628 3148
rect 273680 3136 273686 3188
rect 289262 3136 289268 3188
rect 289320 3176 289326 3188
rect 390646 3176 390652 3188
rect 289320 3148 390652 3176
rect 289320 3136 289326 3148
rect 390646 3136 390652 3148
rect 390704 3136 390710 3188
rect 393958 3136 393964 3188
rect 394016 3176 394022 3188
rect 494698 3176 494704 3188
rect 394016 3148 494704 3176
rect 394016 3136 394022 3148
rect 494698 3136 494704 3148
rect 494756 3136 494762 3188
rect 106918 3068 106924 3120
rect 106976 3108 106982 3120
rect 107562 3108 107568 3120
rect 106976 3080 107568 3108
rect 106976 3068 106982 3080
rect 107562 3068 107568 3080
rect 107620 3068 107626 3120
rect 108114 3068 108120 3120
rect 108172 3108 108178 3120
rect 108942 3108 108948 3120
rect 108172 3080 108948 3108
rect 108172 3068 108178 3080
rect 108942 3068 108948 3080
rect 109000 3068 109006 3120
rect 110506 3068 110512 3120
rect 110564 3108 110570 3120
rect 243078 3108 243084 3120
rect 110564 3080 243084 3108
rect 110564 3068 110570 3080
rect 243078 3068 243084 3080
rect 243136 3068 243142 3120
rect 269758 3068 269764 3120
rect 269816 3108 269822 3120
rect 340966 3108 340972 3120
rect 269816 3080 340972 3108
rect 269816 3068 269822 3080
rect 340966 3068 340972 3080
rect 341024 3068 341030 3120
rect 357434 3068 357440 3120
rect 357492 3108 357498 3120
rect 358722 3108 358728 3120
rect 357492 3080 358728 3108
rect 357492 3068 357498 3080
rect 358722 3068 358728 3080
rect 358780 3068 358786 3120
rect 365714 3068 365720 3120
rect 365772 3108 365778 3120
rect 367002 3108 367008 3120
rect 365772 3080 367008 3108
rect 365772 3068 365778 3080
rect 367002 3068 367008 3080
rect 367060 3068 367066 3120
rect 373994 3068 374000 3120
rect 374052 3108 374058 3120
rect 375282 3108 375288 3120
rect 374052 3080 375288 3108
rect 374052 3068 374058 3080
rect 375282 3068 375288 3080
rect 375340 3068 375346 3120
rect 382274 3068 382280 3120
rect 382332 3108 382338 3120
rect 383562 3108 383568 3120
rect 382332 3080 383568 3108
rect 382332 3068 382338 3080
rect 383562 3068 383568 3080
rect 383620 3068 383626 3120
rect 400858 3068 400864 3120
rect 400916 3108 400922 3120
rect 501782 3108 501788 3120
rect 400916 3080 501788 3108
rect 400916 3068 400922 3080
rect 501782 3068 501788 3080
rect 501840 3068 501846 3120
rect 114002 3000 114008 3052
rect 114060 3040 114066 3052
rect 114462 3040 114468 3052
rect 114060 3012 114468 3040
rect 114060 3000 114066 3012
rect 114462 3000 114468 3012
rect 114520 3000 114526 3052
rect 115198 3000 115204 3052
rect 115256 3040 115262 3052
rect 115842 3040 115848 3052
rect 115256 3012 115848 3040
rect 115256 3000 115262 3012
rect 115842 3000 115848 3012
rect 115900 3000 115906 3052
rect 123478 3000 123484 3052
rect 123536 3040 123542 3052
rect 124122 3040 124128 3052
rect 123536 3012 124128 3040
rect 123536 3000 123542 3012
rect 124122 3000 124128 3012
rect 124180 3000 124186 3052
rect 124674 3000 124680 3052
rect 124732 3040 124738 3052
rect 125502 3040 125508 3052
rect 124732 3012 125508 3040
rect 124732 3000 124738 3012
rect 125502 3000 125508 3012
rect 125560 3000 125566 3052
rect 125870 3000 125876 3052
rect 125928 3040 125934 3052
rect 126882 3040 126888 3052
rect 125928 3012 126888 3040
rect 125928 3000 125934 3012
rect 126882 3000 126888 3012
rect 126940 3000 126946 3052
rect 126974 3000 126980 3052
rect 127032 3040 127038 3052
rect 128262 3040 128268 3052
rect 127032 3012 128268 3040
rect 127032 3000 127038 3012
rect 128262 3000 128268 3012
rect 128320 3000 128326 3052
rect 128357 3043 128415 3049
rect 128357 3009 128369 3043
rect 128403 3040 128415 3043
rect 245286 3040 245292 3052
rect 128403 3012 245292 3040
rect 128403 3009 128415 3012
rect 128357 3003 128415 3009
rect 245286 3000 245292 3012
rect 245344 3000 245350 3052
rect 249978 3000 249984 3052
rect 250036 3040 250042 3052
rect 252462 3040 252468 3052
rect 250036 3012 252468 3040
rect 250036 3000 250042 3012
rect 252462 3000 252468 3012
rect 252520 3000 252526 3052
rect 271322 3000 271328 3052
rect 271380 3040 271386 3052
rect 277118 3040 277124 3052
rect 271380 3012 277124 3040
rect 271380 3000 271386 3012
rect 277118 3000 277124 3012
rect 277176 3000 277182 3052
rect 289078 3000 289084 3052
rect 289136 3040 289142 3052
rect 351638 3040 351644 3052
rect 289136 3012 351644 3040
rect 289136 3000 289142 3012
rect 351638 3000 351644 3012
rect 351696 3000 351702 3052
rect 391198 3000 391204 3052
rect 391256 3040 391262 3052
rect 491110 3040 491116 3052
rect 391256 3012 491116 3040
rect 391256 3000 391262 3012
rect 491110 3000 491116 3012
rect 491168 3000 491174 3052
rect 121086 2932 121092 2984
rect 121144 2972 121150 2984
rect 245378 2972 245384 2984
rect 121144 2944 245384 2972
rect 121144 2932 121150 2944
rect 245378 2932 245384 2944
rect 245436 2932 245442 2984
rect 253198 2972 253204 2984
rect 248386 2944 253204 2972
rect 117590 2864 117596 2916
rect 117648 2904 117654 2916
rect 128357 2907 128415 2913
rect 128357 2904 128369 2907
rect 117648 2876 128369 2904
rect 117648 2864 117654 2876
rect 128357 2873 128369 2876
rect 128403 2873 128415 2907
rect 128357 2867 128415 2873
rect 130562 2864 130568 2916
rect 130620 2904 130626 2916
rect 131022 2904 131028 2916
rect 130620 2876 131028 2904
rect 130620 2864 130626 2876
rect 131022 2864 131028 2876
rect 131080 2864 131086 2916
rect 132954 2864 132960 2916
rect 133012 2904 133018 2916
rect 133782 2904 133788 2916
rect 133012 2876 133788 2904
rect 133012 2864 133018 2876
rect 133782 2864 133788 2876
rect 133840 2864 133846 2916
rect 134150 2864 134156 2916
rect 134208 2904 134214 2916
rect 135162 2904 135168 2916
rect 134208 2876 135168 2904
rect 134208 2864 134214 2876
rect 135162 2864 135168 2876
rect 135220 2864 135226 2916
rect 140038 2864 140044 2916
rect 140096 2904 140102 2916
rect 140682 2904 140688 2916
rect 140096 2876 140688 2904
rect 140096 2864 140102 2876
rect 140682 2864 140688 2876
rect 140740 2864 140746 2916
rect 143534 2864 143540 2916
rect 143592 2904 143598 2916
rect 144822 2904 144828 2916
rect 143592 2876 144828 2904
rect 143592 2864 143598 2876
rect 144822 2864 144828 2876
rect 144880 2864 144886 2916
rect 147122 2864 147128 2916
rect 147180 2904 147186 2916
rect 147582 2904 147588 2916
rect 147180 2876 147588 2904
rect 147180 2864 147186 2876
rect 147582 2864 147588 2876
rect 147640 2864 147646 2916
rect 148318 2864 148324 2916
rect 148376 2904 148382 2916
rect 148962 2904 148968 2916
rect 148376 2876 148968 2904
rect 148376 2864 148382 2876
rect 148962 2864 148968 2876
rect 149020 2864 149026 2916
rect 150618 2864 150624 2916
rect 150676 2904 150682 2916
rect 151722 2904 151728 2916
rect 150676 2876 151728 2904
rect 150676 2864 150682 2876
rect 151722 2864 151728 2876
rect 151780 2864 151786 2916
rect 151814 2864 151820 2916
rect 151872 2904 151878 2916
rect 153102 2904 153108 2916
rect 151872 2876 153108 2904
rect 151872 2864 151878 2876
rect 153102 2864 153108 2876
rect 153160 2864 153166 2916
rect 155402 2864 155408 2916
rect 155460 2904 155466 2916
rect 155862 2904 155868 2916
rect 155460 2876 155868 2904
rect 155460 2864 155466 2876
rect 155862 2864 155868 2876
rect 155920 2864 155926 2916
rect 157794 2864 157800 2916
rect 157852 2904 157858 2916
rect 158622 2904 158628 2916
rect 157852 2876 158628 2904
rect 157852 2864 157858 2876
rect 158622 2864 158628 2876
rect 158680 2864 158686 2916
rect 158898 2864 158904 2916
rect 158956 2904 158962 2916
rect 160002 2904 160008 2916
rect 158956 2876 160008 2904
rect 158956 2864 158962 2876
rect 160002 2864 160008 2876
rect 160060 2864 160066 2916
rect 164878 2864 164884 2916
rect 164936 2904 164942 2916
rect 165522 2904 165528 2916
rect 164936 2876 165528 2904
rect 164936 2864 164942 2876
rect 165522 2864 165528 2876
rect 165580 2864 165586 2916
rect 168374 2864 168380 2916
rect 168432 2904 168438 2916
rect 169570 2904 169576 2916
rect 168432 2876 169576 2904
rect 168432 2864 168438 2876
rect 169570 2864 169576 2876
rect 169628 2864 169634 2916
rect 171962 2864 171968 2916
rect 172020 2904 172026 2916
rect 172020 2876 176608 2904
rect 172020 2864 172026 2876
rect 175458 2796 175464 2848
rect 175516 2836 175522 2848
rect 175516 2808 176516 2836
rect 175516 2796 175522 2808
rect 176488 2700 176516 2808
rect 176580 2768 176608 2876
rect 176654 2864 176660 2916
rect 176712 2904 176718 2916
rect 177850 2904 177856 2916
rect 176712 2876 177856 2904
rect 176712 2864 176718 2876
rect 177850 2864 177856 2876
rect 177908 2864 177914 2916
rect 233970 2904 233976 2916
rect 177960 2876 233976 2904
rect 177960 2768 177988 2876
rect 233970 2864 233976 2876
rect 234028 2864 234034 2916
rect 237006 2864 237012 2916
rect 237064 2904 237070 2916
rect 248386 2904 248414 2944
rect 253198 2932 253204 2944
rect 253256 2932 253262 2984
rect 289170 2932 289176 2984
rect 289228 2972 289234 2984
rect 344554 2972 344560 2984
rect 289228 2944 344560 2972
rect 289228 2932 289234 2944
rect 344554 2932 344560 2944
rect 344612 2932 344618 2984
rect 415394 2932 415400 2984
rect 415452 2972 415458 2984
rect 416682 2972 416688 2984
rect 415452 2944 416688 2972
rect 415452 2932 415458 2944
rect 416682 2932 416688 2944
rect 416740 2932 416746 2984
rect 417510 2932 417516 2984
rect 417568 2972 417574 2984
rect 469858 2972 469864 2984
rect 417568 2944 469864 2972
rect 417568 2932 417574 2944
rect 469858 2932 469864 2944
rect 469916 2932 469922 2984
rect 237064 2876 248414 2904
rect 237064 2864 237070 2876
rect 248782 2864 248788 2916
rect 248840 2904 248846 2916
rect 253290 2904 253296 2916
rect 248840 2876 253296 2904
rect 248840 2864 248846 2876
rect 253290 2864 253296 2876
rect 253348 2864 253354 2916
rect 286410 2864 286416 2916
rect 286468 2904 286474 2916
rect 337470 2904 337476 2916
rect 286468 2876 337476 2904
rect 286468 2864 286474 2876
rect 337470 2864 337476 2876
rect 337528 2864 337534 2916
rect 409230 2864 409236 2916
rect 409288 2904 409294 2916
rect 455690 2904 455696 2916
rect 409288 2876 455696 2904
rect 409288 2864 409294 2876
rect 455690 2864 455696 2876
rect 455748 2864 455754 2916
rect 233786 2836 233792 2848
rect 176580 2740 177988 2768
rect 178052 2808 233792 2836
rect 178052 2700 178080 2808
rect 233786 2796 233792 2808
rect 233844 2796 233850 2848
rect 233881 2839 233939 2845
rect 233881 2805 233893 2839
rect 233927 2836 233939 2839
rect 241054 2836 241060 2848
rect 233927 2808 241060 2836
rect 233927 2805 233939 2808
rect 233881 2799 233939 2805
rect 241054 2796 241060 2808
rect 241112 2796 241118 2848
rect 282178 2796 282184 2848
rect 282236 2836 282242 2848
rect 323302 2836 323308 2848
rect 282236 2808 323308 2836
rect 282236 2796 282242 2808
rect 323302 2796 323308 2808
rect 323360 2796 323366 2848
rect 324314 2796 324320 2848
rect 324372 2836 324378 2848
rect 325602 2836 325608 2848
rect 324372 2808 325608 2836
rect 324372 2796 324378 2808
rect 325602 2796 325608 2808
rect 325660 2796 325666 2848
rect 332594 2796 332600 2848
rect 332652 2836 332658 2848
rect 333882 2836 333888 2848
rect 332652 2808 333888 2836
rect 332652 2796 332658 2808
rect 333882 2796 333888 2808
rect 333940 2796 333946 2848
rect 414658 2796 414664 2848
rect 414716 2836 414722 2848
rect 459186 2836 459192 2848
rect 414716 2808 459192 2836
rect 414716 2796 414722 2808
rect 459186 2796 459192 2808
rect 459244 2796 459250 2848
rect 176488 2672 178080 2700
<< via1 >>
rect 105452 700952 105504 701004
rect 262220 700952 262272 701004
rect 256516 700884 256568 700936
rect 429844 700884 429896 700936
rect 89168 700816 89220 700868
rect 262312 700816 262364 700868
rect 72976 700748 73028 700800
rect 262496 700748 262548 700800
rect 256424 700680 256476 700732
rect 462320 700680 462372 700732
rect 256608 700612 256660 700664
rect 478512 700612 478564 700664
rect 40500 700544 40552 700596
rect 263692 700544 263744 700596
rect 24308 700476 24360 700528
rect 263600 700476 263652 700528
rect 283656 700476 283708 700528
rect 300124 700476 300176 700528
rect 8116 700408 8168 700460
rect 263784 700408 263836 700460
rect 269764 700408 269816 700460
rect 283840 700408 283892 700460
rect 283932 700408 283984 700460
rect 364984 700408 365036 700460
rect 255136 700340 255188 700392
rect 527180 700340 527232 700392
rect 255044 700272 255096 700324
rect 543464 700272 543516 700324
rect 257712 700204 257764 700256
rect 413652 700204 413704 700256
rect 257804 700136 257856 700188
rect 397460 700136 397512 700188
rect 137836 700068 137888 700120
rect 260932 700068 260984 700120
rect 154120 700000 154172 700052
rect 262404 700000 262456 700052
rect 170312 699932 170364 699984
rect 260840 699932 260892 699984
rect 259184 699864 259236 699916
rect 348792 699864 348844 699916
rect 235172 699796 235224 699848
rect 235908 699796 235960 699848
rect 257896 699796 257948 699848
rect 332508 699796 332560 699848
rect 202788 699728 202840 699780
rect 259644 699728 259696 699780
rect 218980 699660 219032 699712
rect 261024 699660 261076 699712
rect 261484 699660 261536 699712
rect 267648 699660 267700 699712
rect 283564 699660 283616 699712
rect 283932 699660 283984 699712
rect 253572 696940 253624 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 264980 683204 265032 683256
rect 253756 683136 253808 683188
rect 580172 683136 580224 683188
rect 3424 670760 3476 670812
rect 265072 670760 265124 670812
rect 253664 670692 253716 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 265164 656888 265216 656940
rect 252468 643084 252520 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 266360 632068 266412 632120
rect 252376 630640 252428 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 266452 618264 266504 618316
rect 252284 616836 252336 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 266544 605820 266596 605872
rect 251088 590656 251140 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 266636 579640 266688 579692
rect 250996 576852 251048 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 267740 565836 267792 565888
rect 250904 563048 250956 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 267832 553392 267884 553444
rect 249708 536800 249760 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 267924 527144 267976 527196
rect 249616 524424 249668 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 269120 514768 269172 514820
rect 249524 510620 249576 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 269212 500964 269264 501016
rect 248328 484372 248380 484424
rect 580172 484372 580224 484424
rect 3424 474716 3476 474768
rect 269304 474716 269356 474768
rect 249432 470568 249484 470620
rect 579988 470568 580040 470620
rect 3240 462340 3292 462392
rect 270776 462340 270828 462392
rect 248236 456764 248288 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 270592 448536 270644 448588
rect 259276 434664 259328 434716
rect 261484 434664 261536 434716
rect 246948 430584 247000 430636
rect 580172 430584 580224 430636
rect 3424 422288 3476 422340
rect 270684 422288 270736 422340
rect 248144 418140 248196 418192
rect 580172 418140 580224 418192
rect 3148 409844 3200 409896
rect 271880 409844 271932 409896
rect 246856 404336 246908 404388
rect 580172 404336 580224 404388
rect 3424 397468 3476 397520
rect 270500 397468 270552 397520
rect 260840 391620 260892 391672
rect 261116 391620 261168 391672
rect 235908 391484 235960 391536
rect 259828 391552 259880 391604
rect 259644 391484 259696 391536
rect 269764 391484 269816 391536
rect 259184 391416 259236 391468
rect 283656 391416 283708 391468
rect 257896 391348 257948 391400
rect 283564 391348 283616 391400
rect 255228 391280 255280 391332
rect 494060 391280 494112 391332
rect 253848 391212 253900 391264
rect 558920 391212 558972 391264
rect 242072 390464 242124 390516
rect 262312 390600 262364 390652
rect 263232 390600 263284 390652
rect 249340 390532 249392 390584
rect 249708 390532 249760 390584
rect 250812 390532 250864 390584
rect 251088 390532 251140 390584
rect 260932 390532 260984 390584
rect 261576 390532 261628 390584
rect 262220 390532 262272 390584
rect 262496 390532 262548 390584
rect 263600 390532 263652 390584
rect 264428 390532 264480 390584
rect 265072 390532 265124 390584
rect 265716 390532 265768 390584
rect 266452 390532 266504 390584
rect 266912 390532 266964 390584
rect 267740 390532 267792 390584
rect 268200 390532 268252 390584
rect 269120 390532 269172 390584
rect 269488 390532 269540 390584
rect 270684 390532 270736 390584
rect 271144 390532 271196 390584
rect 246304 390396 246356 390448
rect 289084 390464 289136 390516
rect 245016 390328 245068 390380
rect 288992 390396 289044 390448
rect 240048 390260 240100 390312
rect 247500 390260 247552 390312
rect 248144 390260 248196 390312
rect 537484 390328 537536 390380
rect 243820 390192 243872 390244
rect 248972 390260 249024 390312
rect 249432 390260 249484 390312
rect 250444 390260 250496 390312
rect 250904 390260 250956 390312
rect 252100 390260 252152 390312
rect 252468 390260 252520 390312
rect 252928 390260 252980 390312
rect 253664 390260 253716 390312
rect 254584 390260 254636 390312
rect 255136 390260 255188 390312
rect 256240 390260 256292 390312
rect 256608 390260 256660 390312
rect 257068 390260 257120 390312
rect 257804 390260 257856 390312
rect 286968 390260 287020 390312
rect 286784 390192 286836 390244
rect 242532 390124 242584 390176
rect 289728 390124 289780 390176
rect 238668 390056 238720 390108
rect 286600 390056 286652 390108
rect 241152 389988 241204 390040
rect 289636 389988 289688 390040
rect 4712 389920 4764 389972
rect 5356 389852 5408 389904
rect 270500 389920 270552 389972
rect 271512 389920 271564 389972
rect 271604 389920 271656 389972
rect 276940 389920 276992 389972
rect 6552 389784 6604 389836
rect 270224 389784 270276 389836
rect 273260 389852 273312 389904
rect 275652 389784 275704 389836
rect 5172 389716 5224 389768
rect 276480 389716 276532 389768
rect 6460 389648 6512 389700
rect 278228 389648 278280 389700
rect 5080 389580 5132 389632
rect 277768 389580 277820 389632
rect 284208 389580 284260 389632
rect 292212 389580 292264 389632
rect 6368 389512 6420 389564
rect 279424 389512 279476 389564
rect 284116 389512 284168 389564
rect 292120 389512 292172 389564
rect 4988 389444 5040 389496
rect 279056 389444 279108 389496
rect 283748 389444 283800 389496
rect 298836 389444 298888 389496
rect 6276 389376 6328 389428
rect 280712 389376 280764 389428
rect 285036 389376 285088 389428
rect 292028 389376 292080 389428
rect 4896 389308 4948 389360
rect 280252 389308 280304 389360
rect 283288 389308 283340 389360
rect 294604 389308 294656 389360
rect 243360 389240 243412 389292
rect 537576 389240 537628 389292
rect 6644 389172 6696 389224
rect 274640 389172 274692 389224
rect 282828 389172 282880 389224
rect 293316 389172 293368 389224
rect 5448 389104 5500 389156
rect 272800 389104 272852 389156
rect 3332 389036 3384 389088
rect 272340 389036 272392 389088
rect 4068 388968 4120 389020
rect 273628 388968 273680 389020
rect 245476 388900 245528 388952
rect 286416 388900 286468 388952
rect 239588 388832 239640 388884
rect 286876 388832 286928 388884
rect 239220 388764 239272 388816
rect 286692 388764 286744 388816
rect 3976 388696 4028 388748
rect 273996 388696 274048 388748
rect 5264 388628 5316 388680
rect 275284 388628 275336 388680
rect 3884 388560 3936 388612
rect 274824 388560 274876 388612
rect 3792 388492 3844 388544
rect 276112 388492 276164 388544
rect 3700 388424 3752 388476
rect 277492 388424 277544 388476
rect 3608 388356 3660 388408
rect 278780 388356 278832 388408
rect 3516 388288 3568 388340
rect 279884 388288 279936 388340
rect 245568 388220 245620 388272
rect 580172 388220 580224 388272
rect 244326 388152 244378 388204
rect 249156 388152 249208 388204
rect 249524 388152 249576 388204
rect 580908 388152 580960 388204
rect 243958 388084 244010 388136
rect 580816 388084 580868 388136
rect 242808 388016 242860 388068
rect 580724 388016 580776 388068
rect 240416 387948 240468 388000
rect 240876 387923 240928 387932
rect 240876 387889 240885 387923
rect 240885 387889 240919 387923
rect 240919 387889 240928 387923
rect 240876 387880 240928 387889
rect 241244 387948 241296 388000
rect 580632 387948 580684 388000
rect 580540 387880 580592 387932
rect 236736 387855 236788 387864
rect 236736 387821 236745 387855
rect 236745 387821 236779 387855
rect 236779 387821 236788 387855
rect 236736 387812 236788 387821
rect 238392 387812 238444 387864
rect 580448 387812 580500 387864
rect 287612 387132 287664 387184
rect 294696 387132 294748 387184
rect 298744 386656 298796 386708
rect 234896 386452 234948 386504
rect 295984 386588 296036 386640
rect 287612 386452 287664 386504
rect 293408 386452 293460 386504
rect 580264 386384 580316 386436
rect 287520 385636 287572 385688
rect 293500 385636 293552 385688
rect 287612 385364 287664 385416
rect 293592 385364 293644 385416
rect 288348 385024 288400 385076
rect 438124 385024 438176 385076
rect 288348 383664 288400 383716
rect 299020 383664 299072 383716
rect 287612 382372 287664 382424
rect 294880 382372 294932 382424
rect 288348 382304 288400 382356
rect 294788 382304 294840 382356
rect 288164 380944 288216 380996
rect 298928 380944 298980 380996
rect 288348 380876 288400 380928
rect 537116 380876 537168 380928
rect 288348 379720 288400 379772
rect 290832 379720 290884 379772
rect 288256 379516 288308 379568
rect 370504 379516 370556 379568
rect 288348 378224 288400 378276
rect 353944 378224 353996 378276
rect 288256 378156 288308 378208
rect 356704 378156 356756 378208
rect 288348 376796 288400 376848
rect 349804 376796 349856 376848
rect 288256 376728 288308 376780
rect 352656 376728 352708 376780
rect 288164 375436 288216 375488
rect 342904 375436 342956 375488
rect 288348 375368 288400 375420
rect 345664 375368 345716 375420
rect 288164 374076 288216 374128
rect 338764 374076 338816 374128
rect 288348 374008 288400 374060
rect 340144 374008 340196 374060
rect 288348 372716 288400 372768
rect 453304 372716 453356 372768
rect 288164 372648 288216 372700
rect 454684 372648 454736 372700
rect 288256 372580 288308 372632
rect 496820 372580 496872 372632
rect 288256 371220 288308 371272
rect 450544 371220 450596 371272
rect 287612 369928 287664 369980
rect 488540 369928 488592 369980
rect 288348 369860 288400 369912
rect 489920 369860 489972 369912
rect 287612 368568 287664 368620
rect 485044 368568 485096 368620
rect 288256 368500 288308 368552
rect 486424 368500 486476 368552
rect 287980 367140 288032 367192
rect 440976 367140 441028 367192
rect 288348 367072 288400 367124
rect 440884 367072 440936 367124
rect 289084 365644 289136 365696
rect 580172 365644 580224 365696
rect 288348 364352 288400 364404
rect 478880 364352 478932 364404
rect 288164 362992 288216 363044
rect 363604 362992 363656 363044
rect 287152 362924 287204 362976
rect 367744 362924 367796 362976
rect 288256 361700 288308 361752
rect 360844 361700 360896 361752
rect 288348 361632 288400 361684
rect 472072 361632 472124 361684
rect 288164 361564 288216 361616
rect 474740 361564 474792 361616
rect 288164 360272 288216 360324
rect 359464 360272 359516 360324
rect 288348 360204 288400 360256
rect 470600 360204 470652 360256
rect 288348 358776 288400 358828
rect 449164 358776 449216 358828
rect 2780 358436 2832 358488
rect 4712 358436 4764 358488
rect 288164 358300 288216 358352
rect 467840 358300 467892 358352
rect 287336 358232 287388 358284
rect 480260 358232 480312 358284
rect 287428 358164 287480 358216
rect 481640 358164 481692 358216
rect 287520 358096 287572 358148
rect 483020 358096 483072 358148
rect 287704 358028 287756 358080
rect 491300 358028 491352 358080
rect 288256 357484 288308 357536
rect 297456 357484 297508 357536
rect 288348 357416 288400 357468
rect 297364 357416 297416 357468
rect 287612 356260 287664 356312
rect 296260 356260 296312 356312
rect 287428 356056 287480 356108
rect 296168 356056 296220 356108
rect 287980 354764 288032 354816
rect 300216 354764 300268 354816
rect 288348 354696 288400 354748
rect 438216 354696 438268 354748
rect 287612 353744 287664 353796
rect 296352 353744 296404 353796
rect 286416 353200 286468 353252
rect 580172 353200 580224 353252
rect 288348 351908 288400 351960
rect 300400 351908 300452 351960
rect 288348 350616 288400 350668
rect 300308 350616 300360 350668
rect 288072 350548 288124 350600
rect 439688 350548 439740 350600
rect 287704 350276 287756 350328
rect 287980 350276 288032 350328
rect 288256 349256 288308 349308
rect 296444 349256 296496 349308
rect 288348 349120 288400 349172
rect 300492 349120 300544 349172
rect 288256 347896 288308 347948
rect 296536 347896 296588 347948
rect 288348 347760 288400 347812
rect 299112 347760 299164 347812
rect 288348 346672 288400 346724
rect 294972 346672 295024 346724
rect 287612 346400 287664 346452
rect 295064 346400 295116 346452
rect 2780 345856 2832 345908
rect 5448 345856 5500 345908
rect 287336 345108 287388 345160
rect 299296 345108 299348 345160
rect 288348 345040 288400 345092
rect 352564 345040 352616 345092
rect 288164 343680 288216 343732
rect 295156 343680 295208 343732
rect 288348 342252 288400 342304
rect 299204 342252 299256 342304
rect 288348 340960 288400 341012
rect 297640 340960 297692 341012
rect 287704 340892 287756 340944
rect 297548 340892 297600 340944
rect 288348 339532 288400 339584
rect 296628 339532 296680 339584
rect 288256 339464 288308 339516
rect 297732 339464 297784 339516
rect 288256 338172 288308 338224
rect 300584 338172 300636 338224
rect 269718 338104 269770 338156
rect 288348 338104 288400 338156
rect 439780 338104 439832 338156
rect 234804 337900 234856 337952
rect 235218 337900 235270 337952
rect 235678 337900 235730 337952
rect 235954 337900 236006 337952
rect 236506 337900 236558 337952
rect 237518 337900 237570 337952
rect 237610 337900 237662 337952
rect 234988 337832 235040 337884
rect 235816 337628 235868 337680
rect 236782 337832 236834 337884
rect 236966 337832 237018 337884
rect 237886 337832 237938 337884
rect 237978 337764 238030 337816
rect 236920 337628 236972 337680
rect 237656 337628 237708 337680
rect 238622 337900 238674 337952
rect 238806 337900 238858 337952
rect 238898 337900 238950 337952
rect 239450 337900 239502 337952
rect 240462 337900 240514 337952
rect 241750 337900 241802 337952
rect 242118 337900 242170 337952
rect 242670 337900 242722 337952
rect 242854 337900 242906 337952
rect 243314 337900 243366 337952
rect 243498 337900 243550 337952
rect 243774 337900 243826 337952
rect 244510 337900 244562 337952
rect 245062 337900 245114 337952
rect 245154 337900 245206 337952
rect 245338 337900 245390 337952
rect 247362 337900 247414 337952
rect 248190 337900 248242 337952
rect 249754 337900 249806 337952
rect 249846 337900 249898 337952
rect 250766 337900 250818 337952
rect 250858 337900 250910 337952
rect 251502 337900 251554 337952
rect 252606 337900 252658 337952
rect 254262 337900 254314 337952
rect 254906 337900 254958 337952
rect 255090 337900 255142 337952
rect 256194 337900 256246 337952
rect 257390 337900 257442 337952
rect 257574 337900 257626 337952
rect 257758 337900 257810 337952
rect 257850 337900 257902 337952
rect 258862 337900 258914 337952
rect 259138 337900 259190 337952
rect 260150 337900 260202 337952
rect 260242 337900 260294 337952
rect 261806 337900 261858 337952
rect 261990 337900 262042 337952
rect 263646 337900 263698 337952
rect 264934 337900 264986 337952
rect 267234 337900 267286 337952
rect 267326 337900 267378 337952
rect 268246 337900 268298 337952
rect 269994 337900 270046 337952
rect 270178 337900 270230 337952
rect 270638 337900 270690 337952
rect 270730 337900 270782 337952
rect 271282 337900 271334 337952
rect 271374 337900 271426 337952
rect 272662 337900 272714 337952
rect 239174 337832 239226 337884
rect 238852 337764 238904 337816
rect 238392 337628 238444 337680
rect 239036 337628 239088 337680
rect 241106 337832 241158 337884
rect 241474 337832 241526 337884
rect 239496 337764 239548 337816
rect 240554 337764 240606 337816
rect 240876 337739 240928 337748
rect 240876 337705 240885 337739
rect 240885 337705 240919 337739
rect 240919 337705 240928 337739
rect 240876 337696 240928 337705
rect 240508 337628 240560 337680
rect 241704 337628 241756 337680
rect 237932 337560 237984 337612
rect 236460 337492 236512 337544
rect 240692 337535 240744 337544
rect 240692 337501 240701 337535
rect 240701 337501 240735 337535
rect 240735 337501 240744 337535
rect 240692 337492 240744 337501
rect 241520 337492 241572 337544
rect 242486 337832 242538 337884
rect 243176 337832 243228 337884
rect 243958 337832 244010 337884
rect 244234 337832 244286 337884
rect 242302 337764 242354 337816
rect 242946 337764 242998 337816
rect 243406 337764 243458 337816
rect 242256 337628 242308 337680
rect 242532 337628 242584 337680
rect 243452 337628 243504 337680
rect 243912 337628 243964 337680
rect 244096 337628 244148 337680
rect 244694 337832 244746 337884
rect 244878 337832 244930 337884
rect 246350 337832 246402 337884
rect 246534 337832 246586 337884
rect 247270 337832 247322 337884
rect 247454 337832 247506 337884
rect 247776 337832 247828 337884
rect 248098 337832 248150 337884
rect 244786 337764 244838 337816
rect 245476 337807 245528 337816
rect 245476 337773 245485 337807
rect 245485 337773 245519 337807
rect 245519 337773 245528 337807
rect 245476 337764 245528 337773
rect 245614 337764 245666 337816
rect 245798 337764 245850 337816
rect 247086 337764 247138 337816
rect 244556 337628 244608 337680
rect 244740 337628 244792 337680
rect 244832 337628 244884 337680
rect 246396 337628 246448 337680
rect 246488 337628 246540 337680
rect 247040 337628 247092 337680
rect 247316 337628 247368 337680
rect 247638 337764 247690 337816
rect 248374 337832 248426 337884
rect 248558 337832 248610 337884
rect 250398 337832 250450 337884
rect 247960 337628 248012 337680
rect 248328 337696 248380 337748
rect 251042 337832 251094 337884
rect 251686 337832 251738 337884
rect 250214 337764 250266 337816
rect 250812 337764 250864 337816
rect 250076 337739 250128 337748
rect 250076 337705 250085 337739
rect 250085 337705 250119 337739
rect 250119 337705 250128 337739
rect 250076 337696 250128 337705
rect 248420 337628 248472 337680
rect 250260 337628 250312 337680
rect 242808 337603 242860 337612
rect 242808 337569 242817 337603
rect 242817 337569 242851 337603
rect 242851 337569 242860 337603
rect 242808 337560 242860 337569
rect 245200 337603 245252 337612
rect 245200 337569 245209 337603
rect 245209 337569 245243 337603
rect 245243 337569 245252 337603
rect 245200 337560 245252 337569
rect 248144 337560 248196 337612
rect 250076 337560 250128 337612
rect 251272 337739 251324 337748
rect 251272 337705 251281 337739
rect 251281 337705 251315 337739
rect 251315 337705 251324 337739
rect 251272 337696 251324 337705
rect 252054 337832 252106 337884
rect 252790 337832 252842 337884
rect 253066 337832 253118 337884
rect 253342 337832 253394 337884
rect 254446 337832 254498 337884
rect 253204 337628 253256 337680
rect 254078 337764 254130 337816
rect 255366 337832 255418 337884
rect 255458 337832 255510 337884
rect 255826 337832 255878 337884
rect 256102 337832 256154 337884
rect 254400 337628 254452 337680
rect 254952 337628 255004 337680
rect 255044 337628 255096 337680
rect 251824 337560 251876 337612
rect 255780 337560 255832 337612
rect 251640 337492 251692 337544
rect 255596 337535 255648 337544
rect 255596 337501 255605 337535
rect 255605 337501 255639 337535
rect 255639 337501 255648 337535
rect 255596 337492 255648 337501
rect 255872 337492 255924 337544
rect 257482 337764 257534 337816
rect 258034 337832 258086 337884
rect 258586 337832 258638 337884
rect 257804 337696 257856 337748
rect 257620 337628 257672 337680
rect 257160 337603 257212 337612
rect 257160 337569 257169 337603
rect 257169 337569 257203 337603
rect 257203 337569 257212 337603
rect 257160 337560 257212 337569
rect 259874 337832 259926 337884
rect 260058 337832 260110 337884
rect 260886 337832 260938 337884
rect 261438 337832 261490 337884
rect 262174 337832 262226 337884
rect 262634 337832 262686 337884
rect 263462 337832 263514 337884
rect 259000 337628 259052 337680
rect 259184 337560 259236 337612
rect 259920 337560 259972 337612
rect 256240 337492 256292 337544
rect 261760 337764 261812 337816
rect 262082 337764 262134 337816
rect 262542 337764 262594 337816
rect 261576 337628 261628 337680
rect 262128 337628 262180 337680
rect 263830 337764 263882 337816
rect 263784 337628 263836 337680
rect 264198 337832 264250 337884
rect 264566 337832 264618 337884
rect 265670 337832 265722 337884
rect 265854 337832 265906 337884
rect 266866 337832 266918 337884
rect 266958 337832 267010 337884
rect 267142 337832 267194 337884
rect 260840 337560 260892 337612
rect 264060 337560 264112 337612
rect 264428 337560 264480 337612
rect 265716 337628 265768 337680
rect 265992 337628 266044 337680
rect 266820 337628 266872 337680
rect 267464 337832 267516 337884
rect 267878 337832 267930 337884
rect 268890 337832 268942 337884
rect 269258 337832 269310 337884
rect 269442 337832 269494 337884
rect 269764 337832 269816 337884
rect 270270 337832 270322 337884
rect 270546 337832 270598 337884
rect 272110 337832 272162 337884
rect 272294 337832 272346 337884
rect 272478 337832 272530 337884
rect 276342 337900 276394 337952
rect 276526 337900 276578 337952
rect 278274 337900 278326 337952
rect 279470 337900 279522 337952
rect 279654 337900 279706 337952
rect 280666 337900 280718 337952
rect 281862 337900 281914 337952
rect 283150 337900 283202 337952
rect 283334 337900 283386 337952
rect 283426 337900 283478 337952
rect 284070 337900 284122 337952
rect 286416 337900 286468 337952
rect 273030 337832 273082 337884
rect 273766 337832 273818 337884
rect 274226 337832 274278 337884
rect 274870 337832 274922 337884
rect 275146 337832 275198 337884
rect 275238 337832 275290 337884
rect 277354 337832 277406 337884
rect 277906 337832 277958 337884
rect 267464 337696 267516 337748
rect 268292 337696 268344 337748
rect 267004 337628 267056 337680
rect 268292 337560 268344 337612
rect 269396 337628 269448 337680
rect 269580 337560 269632 337612
rect 260196 337492 260248 337544
rect 271650 337764 271702 337816
rect 272570 337764 272622 337816
rect 272846 337764 272898 337816
rect 272892 337628 272944 337680
rect 272432 337560 272484 337612
rect 274042 337764 274094 337816
rect 274456 337764 274508 337816
rect 274456 337628 274508 337680
rect 274364 337603 274416 337612
rect 274364 337569 274373 337603
rect 274373 337569 274407 337603
rect 274407 337569 274416 337603
rect 274364 337560 274416 337569
rect 274732 337560 274784 337612
rect 270776 337492 270828 337544
rect 272524 337492 272576 337544
rect 272800 337535 272852 337544
rect 272800 337501 272809 337535
rect 272809 337501 272843 337535
rect 272843 337501 272852 337535
rect 272800 337492 272852 337501
rect 274088 337492 274140 337544
rect 277216 337560 277268 337612
rect 278458 337832 278510 337884
rect 279746 337832 279798 337884
rect 280022 337832 280074 337884
rect 280574 337832 280626 337884
rect 280850 337832 280902 337884
rect 280942 337832 280994 337884
rect 281126 337832 281178 337884
rect 281540 337832 281592 337884
rect 282138 337832 282190 337884
rect 282782 337832 282834 337884
rect 279608 337671 279660 337680
rect 279608 337637 279617 337671
rect 279617 337637 279651 337671
rect 279651 337637 279660 337671
rect 279608 337628 279660 337637
rect 279884 337628 279936 337680
rect 278136 337560 278188 337612
rect 280896 337696 280948 337748
rect 281080 337628 281132 337680
rect 275468 337492 275520 337544
rect 276756 337492 276808 337544
rect 279240 337492 279292 337544
rect 281770 337764 281822 337816
rect 281632 337560 281684 337612
rect 284162 337832 284214 337884
rect 284438 337832 284490 337884
rect 284944 337832 284996 337884
rect 282828 337628 282880 337680
rect 283196 337628 283248 337680
rect 283288 337628 283340 337680
rect 283472 337628 283524 337680
rect 281724 337492 281776 337544
rect 255504 337467 255556 337476
rect 255504 337433 255513 337467
rect 255513 337433 255547 337467
rect 255547 337433 255556 337467
rect 255504 337424 255556 337433
rect 273260 337424 273312 337476
rect 283748 337424 283800 337476
rect 268200 337356 268252 337408
rect 271880 337356 271932 337408
rect 278780 337356 278832 337408
rect 273352 337263 273404 337272
rect 273352 337229 273361 337263
rect 273361 337229 273395 337263
rect 273395 337229 273404 337263
rect 273352 337220 273404 337229
rect 270960 337152 271012 337204
rect 273720 337084 273772 337136
rect 236644 337016 236696 337068
rect 237196 337016 237248 337068
rect 278872 337016 278924 337068
rect 237840 336991 237892 337000
rect 237840 336957 237849 336991
rect 237849 336957 237883 336991
rect 237883 336957 237892 336991
rect 237840 336948 237892 336957
rect 439504 336948 439556 337000
rect 271512 336880 271564 336932
rect 282460 336880 282512 336932
rect 235264 336744 235316 336796
rect 236000 336744 236052 336796
rect 236184 336744 236236 336796
rect 237104 336744 237156 336796
rect 237748 336744 237800 336796
rect 261668 336812 261720 336864
rect 283104 336880 283156 336932
rect 568580 336880 568632 336932
rect 283196 336812 283248 336864
rect 569960 336812 570012 336864
rect 86868 336676 86920 336728
rect 242164 336676 242216 336728
rect 264612 336676 264664 336728
rect 266176 336676 266228 336728
rect 100668 336608 100720 336660
rect 235356 336608 235408 336660
rect 82728 336540 82780 336592
rect 241888 336540 241940 336592
rect 265256 336540 265308 336592
rect 269212 336608 269264 336660
rect 282920 336744 282972 336796
rect 283288 336744 283340 336796
rect 572720 336744 572772 336796
rect 347780 336676 347832 336728
rect 354680 336608 354732 336660
rect 268568 336540 268620 336592
rect 361580 336540 361632 336592
rect 44088 336472 44140 336524
rect 244280 336472 244332 336524
rect 249156 336472 249208 336524
rect 251180 336472 251232 336524
rect 254492 336472 254544 336524
rect 260748 336472 260800 336524
rect 270868 336472 270920 336524
rect 368480 336472 368532 336524
rect 75828 336404 75880 336456
rect 42708 336336 42760 336388
rect 241244 336404 241296 336456
rect 242992 336404 243044 336456
rect 260840 336404 260892 336456
rect 266452 336404 266504 336456
rect 372620 336404 372672 336456
rect 245568 336336 245620 336388
rect 253940 336336 253992 336388
rect 266912 336336 266964 336388
rect 375380 336336 375432 336388
rect 28908 336268 28960 336320
rect 237288 336268 237340 336320
rect 241704 336268 241756 336320
rect 241888 336268 241940 336320
rect 248880 336268 248932 336320
rect 266452 336268 266504 336320
rect 266544 336268 266596 336320
rect 266728 336268 266780 336320
rect 382280 336268 382332 336320
rect 20628 336200 20680 336252
rect 236552 336200 236604 336252
rect 237012 336200 237064 336252
rect 243360 336200 243412 336252
rect 258816 336200 258868 336252
rect 276020 336200 276072 336252
rect 276940 336200 276992 336252
rect 238484 336132 238536 336184
rect 7564 336064 7616 336116
rect 235540 336064 235592 336116
rect 250536 336132 250588 336184
rect 254952 336132 255004 336184
rect 263876 336132 263928 336184
rect 277676 336200 277728 336252
rect 278688 336200 278740 336252
rect 397460 336200 397512 336252
rect 241704 336064 241756 336116
rect 257252 336064 257304 336116
rect 272248 336064 272300 336116
rect 274916 336064 274968 336116
rect 275744 336064 275796 336116
rect 275836 336107 275888 336116
rect 275836 336073 275845 336107
rect 275845 336073 275879 336107
rect 275879 336073 275888 336107
rect 275836 336064 275888 336073
rect 276112 336064 276164 336116
rect 277584 336064 277636 336116
rect 278504 336064 278556 336116
rect 404360 336132 404412 336184
rect 280344 336064 280396 336116
rect 281264 336064 281316 336116
rect 411260 336064 411312 336116
rect 5448 335996 5500 336048
rect 235448 335996 235500 336048
rect 238576 335996 238628 336048
rect 252560 335996 252612 336048
rect 261392 335996 261444 336048
rect 263600 335996 263652 336048
rect 265992 335996 266044 336048
rect 270316 335996 270368 336048
rect 418160 335996 418212 336048
rect 93768 335928 93820 335980
rect 241980 335928 242032 335980
rect 243820 335928 243872 335980
rect 244372 335928 244424 335980
rect 253480 335928 253532 335980
rect 264152 335928 264204 335980
rect 264704 335928 264756 335980
rect 265624 335928 265676 335980
rect 274824 335928 274876 335980
rect 275836 335928 275888 335980
rect 300124 335928 300176 335980
rect 107568 335860 107620 335912
rect 243912 335860 243964 335912
rect 257252 335860 257304 335912
rect 260472 335860 260524 335912
rect 262404 335860 262456 335912
rect 270500 335860 270552 335912
rect 275100 335860 275152 335912
rect 275744 335860 275796 335912
rect 276112 335860 276164 335912
rect 276848 335860 276900 335912
rect 277216 335860 277268 335912
rect 277584 335860 277636 335912
rect 280252 335860 280304 335912
rect 287612 335860 287664 335912
rect 288256 335860 288308 335912
rect 114468 335792 114520 335844
rect 125508 335724 125560 335776
rect 124128 335656 124180 335708
rect 240784 335792 240836 335844
rect 241520 335792 241572 335844
rect 242348 335792 242400 335844
rect 244188 335792 244240 335844
rect 259736 335792 259788 335844
rect 266544 335792 266596 335844
rect 268016 335792 268068 335844
rect 249156 335724 249208 335776
rect 258080 335724 258132 335776
rect 263232 335767 263284 335776
rect 244648 335656 244700 335708
rect 245108 335656 245160 335708
rect 258172 335656 258224 335708
rect 258356 335656 258408 335708
rect 259460 335656 259512 335708
rect 259736 335656 259788 335708
rect 260012 335656 260064 335708
rect 260380 335656 260432 335708
rect 263232 335733 263241 335767
rect 263241 335733 263275 335767
rect 263275 335733 263284 335767
rect 263232 335724 263284 335733
rect 266636 335724 266688 335776
rect 267096 335724 267148 335776
rect 269120 335724 269172 335776
rect 262680 335656 262732 335708
rect 234252 335588 234304 335640
rect 244556 335588 244608 335640
rect 245384 335588 245436 335640
rect 247776 335588 247828 335640
rect 254952 335588 255004 335640
rect 255136 335588 255188 335640
rect 257068 335588 257120 335640
rect 260104 335588 260156 335640
rect 264152 335588 264204 335640
rect 264704 335588 264756 335640
rect 267648 335588 267700 335640
rect 234068 335520 234120 335572
rect 234160 335452 234212 335504
rect 256792 335452 256844 335504
rect 258080 335452 258132 335504
rect 258264 335452 258316 335504
rect 259460 335520 259512 335572
rect 260288 335520 260340 335572
rect 262864 335563 262916 335572
rect 262864 335529 262873 335563
rect 262873 335529 262907 335563
rect 262907 335529 262916 335563
rect 262864 335520 262916 335529
rect 263140 335520 263192 335572
rect 10968 335384 11020 335436
rect 235724 335384 235776 335436
rect 236000 335384 236052 335436
rect 236368 335384 236420 335436
rect 234344 335316 234396 335368
rect 236184 335316 236236 335368
rect 237196 335316 237248 335368
rect 242992 335384 243044 335436
rect 243176 335384 243228 335436
rect 255136 335384 255188 335436
rect 258448 335384 258500 335436
rect 259092 335384 259144 335436
rect 256608 335316 256660 335368
rect 257068 335316 257120 335368
rect 258356 335316 258408 335368
rect 258724 335316 258776 335368
rect 259552 335452 259604 335504
rect 259828 335452 259880 335504
rect 260472 335452 260524 335504
rect 259276 335384 259328 335436
rect 260012 335384 260064 335436
rect 260840 335384 260892 335436
rect 262128 335384 262180 335436
rect 262496 335384 262548 335436
rect 262864 335384 262916 335436
rect 264520 335520 264572 335572
rect 266912 335452 266964 335504
rect 264244 335384 264296 335436
rect 264704 335384 264756 335436
rect 266360 335384 266412 335436
rect 267188 335520 267240 335572
rect 268476 335520 268528 335572
rect 268568 335520 268620 335572
rect 269120 335520 269172 335572
rect 269488 335520 269540 335572
rect 269212 335452 269264 335504
rect 269856 335520 269908 335572
rect 259920 335316 259972 335368
rect 260380 335316 260432 335368
rect 219348 335248 219400 335300
rect 253204 335248 253256 335300
rect 259092 335248 259144 335300
rect 259276 335291 259328 335300
rect 259276 335257 259285 335291
rect 259285 335257 259319 335291
rect 259319 335257 259328 335291
rect 259276 335248 259328 335257
rect 259828 335248 259880 335300
rect 260656 335316 260708 335368
rect 261300 335316 261352 335368
rect 261576 335316 261628 335368
rect 262588 335316 262640 335368
rect 262956 335316 263008 335368
rect 263140 335316 263192 335368
rect 263416 335316 263468 335368
rect 263692 335316 263744 335368
rect 264612 335316 264664 335368
rect 264888 335316 264940 335368
rect 264980 335316 265032 335368
rect 265900 335316 265952 335368
rect 266636 335316 266688 335368
rect 266820 335316 266872 335368
rect 267096 335316 267148 335368
rect 267556 335316 267608 335368
rect 267924 335316 267976 335368
rect 268384 335316 268436 335368
rect 268568 335384 268620 335436
rect 269028 335384 269080 335436
rect 269304 335384 269356 335436
rect 269856 335384 269908 335436
rect 270040 335384 270092 335436
rect 270408 335384 270460 335436
rect 271052 335656 271104 335708
rect 271328 335384 271380 335436
rect 277216 335767 277268 335776
rect 277216 335733 277225 335767
rect 277225 335733 277259 335767
rect 277259 335733 277268 335767
rect 277216 335724 277268 335733
rect 278872 335724 278924 335776
rect 280068 335724 280120 335776
rect 280620 335724 280672 335776
rect 281448 335724 281500 335776
rect 282000 335724 282052 335776
rect 282644 335724 282696 335776
rect 273720 335588 273772 335640
rect 273628 335520 273680 335572
rect 274180 335520 274232 335572
rect 275008 335520 275060 335572
rect 275560 335520 275612 335572
rect 277400 335520 277452 335572
rect 278320 335520 278372 335572
rect 281172 335656 281224 335708
rect 287520 335792 287572 335844
rect 288164 335792 288216 335844
rect 289084 335724 289136 335776
rect 289176 335656 289228 335708
rect 279148 335588 279200 335640
rect 282644 335588 282696 335640
rect 283012 335588 283064 335640
rect 286416 335588 286468 335640
rect 289268 335588 289320 335640
rect 284852 335520 284904 335572
rect 285404 335520 285456 335572
rect 291844 335520 291896 335572
rect 296076 335860 296128 335912
rect 284392 335384 284444 335436
rect 285312 335384 285364 335436
rect 291936 335384 291988 335436
rect 267372 335248 267424 335300
rect 201408 335180 201460 335232
rect 251916 335180 251968 335232
rect 268752 335316 268804 335368
rect 268936 335316 268988 335368
rect 269396 335316 269448 335368
rect 269672 335316 269724 335368
rect 271052 335316 271104 335368
rect 271696 335316 271748 335368
rect 271972 335316 272024 335368
rect 272340 335316 272392 335368
rect 272616 335316 272668 335368
rect 273076 335316 273128 335368
rect 273536 335316 273588 335368
rect 271604 335248 271656 335300
rect 273996 335316 274048 335368
rect 274272 335316 274324 335368
rect 275468 335316 275520 335368
rect 275928 335316 275980 335368
rect 276940 335359 276992 335368
rect 276940 335325 276949 335359
rect 276949 335325 276983 335359
rect 276983 335325 276992 335359
rect 276940 335316 276992 335325
rect 277032 335316 277084 335368
rect 277308 335316 277360 335368
rect 277492 335316 277544 335368
rect 277952 335316 278004 335368
rect 279424 335316 279476 335368
rect 279884 335316 279936 335368
rect 280160 335316 280212 335368
rect 274180 335248 274232 335300
rect 274732 335248 274784 335300
rect 281724 335316 281776 335368
rect 282184 335316 282236 335368
rect 281356 335248 281408 335300
rect 269948 335223 270000 335232
rect 269948 335189 269957 335223
rect 269957 335189 269991 335223
rect 269991 335189 270000 335223
rect 269948 335180 270000 335189
rect 277308 335223 277360 335232
rect 277308 335189 277317 335223
rect 277317 335189 277351 335223
rect 277351 335189 277360 335223
rect 277308 335180 277360 335189
rect 283012 335316 283064 335368
rect 283564 335316 283616 335368
rect 284024 335316 284076 335368
rect 284208 335316 284260 335368
rect 284484 335316 284536 335368
rect 284852 335316 284904 335368
rect 285036 335316 285088 335368
rect 285496 335316 285548 335368
rect 290464 335316 290516 335368
rect 396724 335248 396776 335300
rect 194416 335112 194468 335164
rect 245108 335112 245160 335164
rect 268936 335155 268988 335164
rect 268936 335121 268945 335155
rect 268945 335121 268979 335155
rect 268979 335121 268988 335155
rect 268936 335112 268988 335121
rect 270224 335112 270276 335164
rect 276664 335112 276716 335164
rect 279424 335112 279476 335164
rect 403624 335180 403676 335232
rect 433984 335112 434036 335164
rect 197268 335044 197320 335096
rect 251548 335044 251600 335096
rect 269488 335044 269540 335096
rect 405740 335044 405792 335096
rect 190368 334976 190420 335028
rect 250904 334976 250956 335028
rect 277860 334976 277912 335028
rect 278320 334976 278372 335028
rect 278688 334976 278740 335028
rect 434076 334976 434128 335028
rect 186136 334908 186188 334960
rect 245844 334908 245896 334960
rect 434168 334908 434220 334960
rect 183468 334840 183520 334892
rect 272064 334840 272116 334892
rect 437480 334840 437532 334892
rect 179328 334772 179380 334824
rect 251364 334772 251416 334824
rect 252468 334772 252520 334824
rect 169576 334704 169628 334756
rect 244280 334704 244332 334756
rect 245108 334704 245160 334756
rect 254952 334704 255004 334756
rect 271880 334704 271932 334756
rect 272064 334704 272116 334756
rect 280068 334704 280120 334756
rect 165528 334636 165580 334688
rect 158628 334568 158680 334620
rect 247408 334636 247460 334688
rect 268200 334636 268252 334688
rect 280160 334636 280212 334688
rect 536840 334772 536892 334824
rect 539600 334704 539652 334756
rect 281632 334636 281684 334688
rect 281816 334636 281868 334688
rect 550640 334636 550692 334688
rect 247592 334568 247644 334620
rect 248788 334568 248840 334620
rect 249432 334568 249484 334620
rect 262220 334568 262272 334620
rect 280804 334568 280856 334620
rect 554780 334568 554832 334620
rect 204168 334500 204220 334552
rect 211068 334432 211120 334484
rect 267832 334500 267884 334552
rect 387800 334500 387852 334552
rect 252100 334432 252152 334484
rect 262220 334475 262272 334484
rect 262220 334441 262229 334475
rect 262229 334441 262263 334475
rect 262263 334441 262272 334475
rect 262220 334432 262272 334441
rect 270500 334432 270552 334484
rect 208308 334364 208360 334416
rect 251364 334364 251416 334416
rect 251916 334364 251968 334416
rect 255412 334364 255464 334416
rect 277584 334432 277636 334484
rect 282644 334432 282696 334484
rect 393964 334432 394016 334484
rect 325700 334364 325752 334416
rect 222108 334296 222160 334348
rect 253664 334296 253716 334348
rect 274548 334296 274600 334348
rect 276664 334296 276716 334348
rect 276848 334296 276900 334348
rect 391204 334296 391256 334348
rect 215208 334228 215260 334280
rect 241704 334228 241756 334280
rect 261208 334228 261260 334280
rect 309140 334228 309192 334280
rect 229008 334160 229060 334212
rect 249156 334160 249208 334212
rect 264152 334160 264204 334212
rect 292580 334160 292632 334212
rect 226248 334092 226300 334144
rect 245568 334092 245620 334144
rect 253572 334092 253624 334144
rect 253756 334092 253808 334144
rect 260288 334092 260340 334144
rect 289360 334092 289412 334144
rect 233976 334024 234028 334076
rect 249524 334024 249576 334076
rect 259368 334024 259420 334076
rect 287704 334024 287756 334076
rect 233884 333956 233936 334008
rect 285036 333956 285088 334008
rect 147588 333888 147640 333940
rect 383660 333888 383712 333940
rect 144736 333820 144788 333872
rect 247224 333820 247276 333872
rect 268936 333820 268988 333872
rect 394700 333820 394752 333872
rect 128268 333752 128320 333804
rect 243728 333752 243780 333804
rect 244924 333795 244976 333804
rect 244924 333761 244933 333795
rect 244933 333761 244967 333795
rect 244967 333761 244976 333795
rect 244924 333752 244976 333761
rect 268660 333752 268712 333804
rect 398840 333752 398892 333804
rect 95148 333684 95200 333736
rect 237012 333684 237064 333736
rect 269120 333684 269172 333736
rect 408500 333684 408552 333736
rect 88248 333616 88300 333668
rect 242440 333616 242492 333668
rect 269212 333616 269264 333668
rect 412640 333616 412692 333668
rect 70308 333548 70360 333600
rect 240876 333548 240928 333600
rect 415400 333548 415452 333600
rect 66168 333480 66220 333532
rect 423680 333480 423732 333532
rect 61936 333412 61988 333464
rect 240232 333412 240284 333464
rect 35900 333344 35952 333396
rect 237932 333344 237984 333396
rect 258172 333344 258224 333396
rect 270868 333344 270920 333396
rect 430580 333412 430632 333464
rect 271604 333344 271656 333396
rect 426440 333344 426492 333396
rect 33140 333276 33192 333328
rect 237748 333276 237800 333328
rect 243268 333276 243320 333328
rect 256976 333276 257028 333328
rect 257988 333276 258040 333328
rect 263968 333276 264020 333328
rect 264520 333276 264572 333328
rect 265256 333276 265308 333328
rect 266268 333276 266320 333328
rect 267740 333319 267792 333328
rect 267740 333285 267749 333319
rect 267749 333285 267783 333319
rect 267783 333285 267792 333319
rect 267740 333276 267792 333285
rect 268660 333276 268712 333328
rect 433340 333276 433392 333328
rect 29000 333208 29052 333260
rect 237288 333208 237340 333260
rect 238208 333208 238260 333260
rect 239036 333208 239088 333260
rect 239956 333208 240008 333260
rect 241244 333208 241296 333260
rect 242164 333208 242216 333260
rect 243544 333208 243596 333260
rect 246580 333208 246632 333260
rect 257252 333208 257304 333260
rect 436744 333208 436796 333260
rect 148968 333140 149020 333192
rect 247316 333140 247368 333192
rect 247408 333140 247460 333192
rect 250168 333140 250220 333192
rect 252376 333140 252428 333192
rect 271512 333140 271564 333192
rect 271696 333140 271748 333192
rect 153108 333072 153160 333124
rect 247960 333072 248012 333124
rect 268108 333072 268160 333124
rect 390652 333140 390704 333192
rect 151728 333004 151780 333056
rect 380900 333072 380952 333124
rect 154488 332936 154540 332988
rect 245384 332936 245436 332988
rect 265716 332936 265768 332988
rect 362960 333004 363012 333056
rect 180708 332868 180760 332920
rect 250260 332868 250312 332920
rect 265348 332868 265400 332920
rect 358820 332936 358872 332988
rect 340972 332868 341024 332920
rect 209688 332800 209740 332852
rect 265072 332800 265124 332852
rect 356060 332800 356112 332852
rect 227628 332732 227680 332784
rect 316132 332732 316184 332784
rect 230388 332664 230440 332716
rect 254308 332664 254360 332716
rect 261668 332664 261720 332716
rect 313280 332664 313332 332716
rect 233148 332596 233200 332648
rect 251180 332596 251232 332648
rect 252100 332596 252152 332648
rect 255780 332596 255832 332648
rect 263692 332596 263744 332648
rect 306380 332596 306432 332648
rect 261024 332528 261076 332580
rect 307760 332528 307812 332580
rect 263600 332460 263652 332512
rect 311900 332460 311952 332512
rect 177856 332392 177908 332444
rect 318800 332392 318852 332444
rect 161388 332324 161440 332376
rect 248420 332324 248472 332376
rect 329840 332324 329892 332376
rect 140688 332256 140740 332308
rect 246764 332256 246816 332308
rect 280160 332256 280212 332308
rect 280344 332256 280396 332308
rect 357440 332256 357492 332308
rect 126888 332188 126940 332240
rect 275284 332188 275336 332240
rect 423772 332188 423824 332240
rect 97908 332120 97960 332172
rect 243452 332120 243504 332172
rect 259552 332120 259604 332172
rect 437020 332120 437072 332172
rect 85488 332052 85540 332104
rect 240784 332052 240836 332104
rect 258816 332052 258868 332104
rect 436928 332052 436980 332104
rect 81348 331984 81400 332036
rect 241888 331984 241940 332036
rect 255136 331984 255188 332036
rect 436836 331984 436888 332036
rect 59268 331916 59320 331968
rect 239864 331916 239916 331968
rect 240784 331916 240836 331968
rect 252560 331916 252612 331968
rect 519544 331916 519596 331968
rect 19248 331848 19300 331900
rect 236460 331848 236512 331900
rect 259276 331848 259328 331900
rect 285680 331848 285732 331900
rect 285772 331848 285824 331900
rect 581000 331848 581052 331900
rect 262404 331780 262456 331832
rect 300860 331780 300912 331832
rect 266452 331712 266504 331764
rect 298100 331712 298152 331764
rect 248972 331644 249024 331696
rect 249248 331644 249300 331696
rect 259644 331644 259696 331696
rect 284944 331644 284996 331696
rect 292304 331644 292356 331696
rect 248880 331576 248932 331628
rect 249340 331576 249392 331628
rect 276480 331576 276532 331628
rect 289544 331576 289596 331628
rect 274272 331508 274324 331560
rect 290648 331508 290700 331560
rect 275376 331440 275428 331492
rect 290924 331440 290976 331492
rect 273260 331372 273312 331424
rect 289452 331372 289504 331424
rect 274824 331304 274876 331356
rect 290740 331304 290792 331356
rect 40040 331236 40092 331288
rect 238300 331236 238352 331288
rect 280252 331236 280304 331288
rect 280988 331236 281040 331288
rect 291200 331236 291252 331288
rect 272156 330692 272208 330744
rect 273812 330624 273864 330676
rect 275376 330624 275428 330676
rect 275652 330624 275704 330676
rect 277860 330692 277912 330744
rect 278044 330692 278096 330744
rect 279056 330692 279108 330744
rect 279700 330692 279752 330744
rect 422944 330624 422996 330676
rect 23388 330488 23440 330540
rect 236828 330488 236880 330540
rect 273720 330284 273772 330336
rect 277768 330556 277820 330608
rect 278044 330556 278096 330608
rect 280988 330556 281040 330608
rect 285588 330556 285640 330608
rect 538220 330556 538272 330608
rect 275652 330488 275704 330540
rect 275836 330488 275888 330540
rect 282368 330488 282420 330540
rect 282920 330488 282972 330540
rect 574100 330488 574152 330540
rect 278964 330420 279016 330472
rect 279884 330420 279936 330472
rect 280344 330420 280396 330472
rect 280896 330420 280948 330472
rect 281540 330420 281592 330472
rect 282276 330420 282328 330472
rect 273904 330216 273956 330268
rect 274088 330148 274140 330200
rect 267004 329060 267056 329112
rect 267280 329060 267332 329112
rect 238300 327700 238352 327752
rect 437112 327700 437164 327752
rect 265164 327632 265216 327684
rect 265532 327632 265584 327684
rect 244648 326748 244700 326800
rect 244832 326748 244884 326800
rect 244740 326680 244792 326732
rect 245844 326680 245896 326732
rect 246028 326680 246080 326732
rect 241612 326476 241664 326528
rect 242716 326476 242768 326528
rect 248696 326544 248748 326596
rect 249156 326544 249208 326596
rect 255412 326544 255464 326596
rect 256424 326544 256476 326596
rect 270960 326544 271012 326596
rect 271328 326544 271380 326596
rect 244832 326476 244884 326528
rect 255504 326476 255556 326528
rect 255780 326476 255832 326528
rect 255964 326476 256016 326528
rect 256148 326476 256200 326528
rect 257436 326476 257488 326528
rect 257804 326476 257856 326528
rect 270500 326476 270552 326528
rect 271420 326476 271472 326528
rect 235632 326408 235684 326460
rect 240692 326451 240744 326460
rect 240692 326417 240701 326451
rect 240701 326417 240735 326451
rect 240735 326417 240744 326451
rect 240692 326408 240744 326417
rect 241796 326408 241848 326460
rect 242624 326408 242676 326460
rect 243084 326408 243136 326460
rect 243912 326408 243964 326460
rect 244556 326408 244608 326460
rect 245016 326408 245068 326460
rect 246120 326408 246172 326460
rect 246396 326408 246448 326460
rect 247316 326408 247368 326460
rect 248144 326408 248196 326460
rect 250260 326408 250312 326460
rect 250812 326408 250864 326460
rect 252744 326408 252796 326460
rect 253296 326408 253348 326460
rect 269764 326408 269816 326460
rect 269948 326408 270000 326460
rect 270960 326408 271012 326460
rect 271144 326408 271196 326460
rect 236460 326340 236512 326392
rect 236920 326340 236972 326392
rect 237656 326340 237708 326392
rect 238116 326340 238168 326392
rect 240416 326340 240468 326392
rect 240876 326340 240928 326392
rect 241888 326340 241940 326392
rect 242256 326340 242308 326392
rect 243360 326340 243412 326392
rect 244004 326340 244056 326392
rect 247500 326340 247552 326392
rect 248328 326340 248380 326392
rect 248696 326340 248748 326392
rect 249708 326340 249760 326392
rect 250352 326340 250404 326392
rect 250628 326340 250680 326392
rect 251548 326340 251600 326392
rect 252468 326340 252520 326392
rect 252836 326340 252888 326392
rect 253020 326340 253072 326392
rect 254124 326340 254176 326392
rect 254768 326340 254820 326392
rect 258540 326340 258592 326392
rect 258908 326340 258960 326392
rect 260288 326340 260340 326392
rect 260564 326340 260616 326392
rect 263876 326340 263928 326392
rect 264244 326340 264296 326392
rect 271420 326340 271472 326392
rect 271604 326340 271656 326392
rect 283472 326340 283524 326392
rect 283840 326340 283892 326392
rect 241704 326272 241756 326324
rect 242808 326272 242860 326324
rect 243084 326272 243136 326324
rect 244188 326272 244240 326324
rect 235724 326204 235776 326256
rect 240416 326204 240468 326256
rect 241152 326204 241204 326256
rect 244464 326204 244516 326256
rect 244740 326204 244792 326256
rect 246028 326204 246080 326256
rect 246948 326204 247000 326256
rect 248880 326204 248932 326256
rect 249064 326204 249116 326256
rect 250352 326204 250404 326256
rect 251088 326204 251140 326256
rect 252652 326204 252704 326256
rect 253296 326204 253348 326256
rect 256056 326204 256108 326256
rect 256424 326204 256476 326256
rect 256884 326204 256936 326256
rect 257804 326204 257856 326256
rect 260196 326204 260248 326256
rect 260564 326204 260616 326256
rect 245936 326136 245988 326188
rect 246856 326136 246908 326188
rect 255596 326136 255648 326188
rect 256516 326136 256568 326188
rect 259644 326136 259696 326188
rect 259828 326136 259880 326188
rect 244464 326068 244516 326120
rect 245476 326068 245528 326120
rect 246212 326068 246264 326120
rect 246672 326068 246724 326120
rect 248512 326068 248564 326120
rect 249064 326068 249116 326120
rect 252744 326068 252796 326120
rect 253664 326068 253716 326120
rect 255320 326068 255372 326120
rect 256240 326068 256292 326120
rect 269120 326068 269172 326120
rect 269764 326068 269816 326120
rect 270868 326068 270920 326120
rect 271328 326068 271380 326120
rect 244924 326000 244976 326052
rect 245292 326000 245344 326052
rect 254676 325932 254728 325984
rect 255228 325932 255280 325984
rect 247224 324368 247276 324420
rect 247868 324368 247920 324420
rect 238944 323824 238996 323876
rect 239680 323824 239732 323876
rect 262864 323416 262916 323468
rect 263140 323416 263192 323468
rect 449164 322872 449216 322924
rect 469404 322872 469456 322924
rect 485044 322872 485096 322924
rect 486332 322872 486384 322924
rect 338764 322804 338816 322856
rect 498200 322804 498252 322856
rect 340144 322736 340196 322788
rect 499212 322736 499264 322788
rect 342904 322668 342956 322720
rect 500684 322668 500736 322720
rect 345664 322600 345716 322652
rect 501236 322600 501288 322652
rect 349804 322532 349856 322584
rect 503260 322532 503312 322584
rect 353944 322464 353996 322516
rect 505468 322464 505520 322516
rect 352656 322396 352708 322448
rect 503812 322396 503864 322448
rect 356704 322328 356756 322380
rect 506940 322328 506992 322380
rect 360844 322260 360896 322312
rect 474556 322260 474608 322312
rect 359464 322192 359516 322244
rect 471980 322192 472032 322244
rect 519544 322192 519596 322244
rect 536932 322192 536984 322244
rect 363604 322124 363656 322176
rect 476764 322124 476816 322176
rect 240784 322056 240836 322108
rect 241428 322056 241480 322108
rect 367744 322056 367796 322108
rect 478236 322056 478288 322108
rect 440884 321988 440936 322040
rect 485412 321988 485464 322040
rect 440976 321920 441028 321972
rect 484400 321920 484452 321972
rect 450544 321852 450596 321904
rect 492772 321852 492824 321904
rect 237748 321784 237800 321836
rect 238668 321784 238720 321836
rect 454684 321784 454736 321836
rect 495532 321784 495584 321836
rect 453304 321716 453356 321768
rect 494244 321716 494296 321768
rect 268384 321648 268436 321700
rect 486424 321580 486476 321632
rect 488172 321580 488224 321632
rect 530032 321580 530084 321632
rect 537024 321580 537076 321632
rect 240692 321079 240744 321088
rect 240692 321045 240701 321079
rect 240701 321045 240735 321079
rect 240735 321045 240744 321079
rect 240692 321036 240744 321045
rect 288992 320832 289044 320884
rect 580908 320832 580960 320884
rect 3332 306212 3384 306264
rect 6644 306212 6696 306264
rect 284852 300092 284904 300144
rect 292396 300092 292448 300144
rect 237748 278740 237800 278792
rect 238116 278740 238168 278792
rect 437388 278740 437440 278792
rect 537576 273164 537628 273216
rect 580172 273164 580224 273216
rect 436928 271940 436980 271992
rect 437112 271940 437164 271992
rect 249248 271804 249300 271856
rect 436928 271804 436980 271856
rect 436928 269016 436980 269068
rect 437112 269016 437164 269068
rect 436836 266772 436888 266824
rect 437204 266772 437256 266824
rect 537484 259360 537536 259412
rect 579804 259360 579856 259412
rect 2780 254600 2832 254652
rect 5356 254600 5408 254652
rect 370504 248344 370556 248396
rect 436100 248344 436152 248396
rect 290832 245556 290884 245608
rect 436100 245556 436152 245608
rect 2780 241340 2832 241392
rect 5264 241340 5316 241392
rect 232780 240728 232832 240780
rect 439412 240728 439464 240780
rect 284024 240048 284076 240100
rect 438584 240048 438636 240100
rect 271972 239980 272024 240032
rect 285312 239912 285364 239964
rect 364340 239912 364392 239964
rect 437296 239980 437348 240032
rect 439872 239980 439924 240032
rect 437112 239912 437164 239964
rect 538496 239912 538548 239964
rect 441436 239844 441488 239896
rect 538312 239844 538364 239896
rect 258448 239776 258500 239828
rect 284300 239776 284352 239828
rect 439780 239776 439832 239828
rect 467840 239776 467892 239828
rect 437388 239708 437440 239760
rect 472072 239708 472124 239760
rect 274180 239640 274232 239692
rect 459560 239640 459612 239692
rect 536932 239640 536984 239692
rect 273996 239572 274048 239624
rect 465172 239572 465224 239624
rect 275560 239504 275612 239556
rect 473360 239504 473412 239556
rect 274732 239436 274784 239488
rect 476120 239436 476172 239488
rect 275376 239368 275428 239420
rect 481732 239368 481784 239420
rect 437020 239300 437072 239352
rect 522856 239300 522908 239352
rect 438768 239232 438820 239284
rect 438676 239164 438728 239216
rect 522672 239232 522724 239284
rect 441528 239164 441580 239216
rect 523132 239164 523184 239216
rect 287796 239096 287848 239148
rect 446404 239096 446456 239148
rect 447048 239096 447100 239148
rect 537024 239096 537076 239148
rect 300584 239028 300636 239080
rect 469220 239028 469272 239080
rect 299296 238960 299348 239012
rect 483020 238960 483072 239012
rect 295156 238892 295208 238944
rect 480444 238892 480496 238944
rect 288164 238824 288216 238876
rect 479156 238824 479208 238876
rect 300400 238756 300452 238808
rect 494244 238756 494296 238808
rect 288256 238688 288308 238740
rect 476764 238688 476816 238740
rect 299112 238620 299164 238672
rect 487804 238620 487856 238672
rect 300492 238552 300544 238604
rect 490564 238552 490616 238604
rect 295064 238484 295116 238536
rect 485412 238484 485464 238536
rect 292120 238416 292172 238468
rect 484860 238416 484912 238468
rect 293592 238348 293644 238400
rect 491668 238348 491720 238400
rect 293500 238280 293552 238332
rect 492772 238280 492824 238332
rect 288072 238212 288124 238264
rect 496820 238212 496872 238264
rect 260012 238144 260064 238196
rect 287060 238144 287112 238196
rect 287980 238144 288032 238196
rect 499212 238144 499264 238196
rect 232596 238076 232648 238128
rect 465080 238076 465132 238128
rect 232688 238008 232740 238060
rect 468300 238008 468352 238060
rect 288348 237940 288400 237992
rect 475660 237940 475712 237992
rect 294604 237872 294656 237924
rect 471796 237872 471848 237924
rect 294788 237804 294840 237856
rect 467196 237804 467248 237856
rect 294880 237736 294932 237788
rect 470692 237736 470744 237788
rect 293316 237668 293368 237720
rect 463700 237668 463752 237720
rect 352564 237600 352616 237652
rect 481640 237600 481692 237652
rect 438216 237532 438268 237584
rect 500960 237532 501012 237584
rect 439688 237464 439740 237516
rect 492680 237464 492732 237516
rect 438124 237396 438176 237448
rect 481916 237396 481968 237448
rect 438584 237328 438636 237380
rect 471980 237328 472032 237380
rect 472072 237328 472124 237380
rect 523040 237328 523092 237380
rect 287888 237260 287940 237312
rect 495440 237260 495492 237312
rect 285496 237192 285548 237244
rect 493324 237192 493376 237244
rect 285404 237124 285456 237176
rect 487160 237124 487212 237176
rect 296352 237056 296404 237108
rect 496820 237056 496872 237108
rect 300216 236988 300268 237040
rect 499856 236988 499908 237040
rect 284760 236920 284812 236972
rect 483020 236920 483072 236972
rect 296444 236852 296496 236904
rect 488540 236852 488592 236904
rect 300308 236784 300360 236836
rect 491300 236784 491352 236836
rect 294972 236716 295024 236768
rect 484400 236716 484452 236768
rect 296536 236648 296588 236700
rect 485780 236648 485832 236700
rect 292304 236580 292356 236632
rect 480260 236580 480312 236632
rect 292396 236512 292448 236564
rect 480536 236512 480588 236564
rect 299204 236444 299256 236496
rect 477500 236444 477552 236496
rect 297548 236376 297600 236428
rect 473452 236376 473504 236428
rect 297640 236308 297692 236360
rect 472072 236308 472124 236360
rect 297732 236240 297784 236292
rect 471980 236240 472032 236292
rect 298928 236172 298980 236224
rect 460940 236172 460992 236224
rect 461584 236172 461636 236224
rect 485780 236172 485832 236224
rect 364340 236104 364392 236156
rect 477592 236104 477644 236156
rect 232504 236036 232556 236088
rect 462320 236036 462372 236088
rect 462412 235968 462464 236020
rect 297364 235900 297416 235952
rect 505100 235900 505152 235952
rect 296260 235832 296312 235884
rect 503720 235832 503772 235884
rect 296168 235764 296220 235816
rect 502432 235764 502484 235816
rect 296628 235696 296680 235748
rect 469220 235696 469272 235748
rect 276388 235356 276440 235408
rect 440240 235356 440292 235408
rect 272800 235288 272852 235340
rect 445760 235288 445812 235340
rect 280528 235220 280580 235272
rect 505100 235220 505152 235272
rect 286968 233180 287020 233232
rect 579988 233180 580040 233232
rect 289728 219376 289780 219428
rect 579988 219376 580040 219428
rect 2964 202784 3016 202836
rect 6552 202784 6604 202836
rect 298744 193128 298796 193180
rect 579620 193128 579672 193180
rect 2780 188912 2832 188964
rect 5172 188912 5224 188964
rect 289636 179324 289688 179376
rect 579620 179324 579672 179376
rect 108948 177624 109000 177676
rect 243360 177624 243412 177676
rect 104808 177556 104860 177608
rect 243268 177556 243320 177608
rect 268568 177556 268620 177608
rect 402980 177556 403032 177608
rect 64788 177488 64840 177540
rect 240876 177488 240928 177540
rect 269672 177488 269724 177540
rect 416780 177488 416832 177540
rect 53656 177420 53708 177472
rect 239220 177420 239272 177472
rect 271052 177420 271104 177472
rect 434720 177420 434772 177472
rect 9588 177352 9640 177404
rect 234896 177352 234948 177404
rect 280712 177352 280764 177404
rect 540980 177352 541032 177404
rect 4068 177284 4120 177336
rect 234988 177284 235040 177336
rect 280620 177284 280672 177336
rect 549260 177284 549312 177336
rect 274088 162120 274140 162172
rect 444380 162120 444432 162172
rect 286876 153144 286928 153196
rect 580172 153144 580224 153196
rect 3148 150356 3200 150408
rect 6460 150356 6512 150408
rect 286784 139340 286836 139392
rect 580172 139340 580224 139392
rect 2780 137232 2832 137284
rect 5080 137232 5132 137284
rect 286692 126896 286744 126948
rect 579620 126896 579672 126948
rect 286600 100648 286652 100700
rect 580172 100648 580224 100700
rect 3240 97860 3292 97912
rect 6368 97860 6420 97912
rect 219256 89088 219308 89140
rect 253204 89088 253256 89140
rect 210976 89020 211028 89072
rect 253296 89020 253348 89072
rect 258816 89020 258868 89072
rect 284392 89020 284444 89072
rect 202696 88952 202748 89004
rect 251824 88952 251876 89004
rect 270776 88952 270828 89004
rect 420920 88952 420972 89004
rect 253388 88680 253440 88732
rect 256148 88680 256200 88732
rect 253204 88272 253256 88324
rect 254492 88272 254544 88324
rect 260288 87796 260340 87848
rect 302240 87796 302292 87848
rect 200028 87728 200080 87780
rect 251732 87728 251784 87780
rect 268660 87728 268712 87780
rect 389180 87728 389232 87780
rect 115848 87660 115900 87712
rect 244832 87660 244884 87712
rect 269948 87660 270000 87712
rect 407212 87660 407264 87712
rect 84108 87592 84160 87644
rect 242072 87592 242124 87644
rect 274272 87592 274324 87644
rect 456800 87592 456852 87644
rect 285128 86912 285180 86964
rect 579620 86912 579672 86964
rect 216588 86436 216640 86488
rect 253112 86436 253164 86488
rect 195888 86368 195940 86420
rect 251640 86368 251692 86420
rect 102048 86300 102100 86352
rect 243176 86300 243228 86352
rect 49608 86232 49660 86284
rect 239128 86232 239180 86284
rect 2780 85212 2832 85264
rect 4988 85212 5040 85264
rect 212448 85076 212500 85128
rect 253020 85076 253072 85128
rect 260932 85076 260984 85128
rect 307852 85076 307904 85128
rect 162768 85008 162820 85060
rect 249156 85008 249208 85060
rect 267004 85008 267056 85060
rect 332600 85008 332652 85060
rect 111708 84940 111760 84992
rect 244740 84940 244792 84992
rect 252468 84940 252520 84992
rect 256056 84940 256108 84992
rect 264152 84940 264204 84992
rect 349160 84940 349212 84992
rect 79968 84872 80020 84924
rect 241980 84872 242032 84924
rect 265348 84872 265400 84924
rect 369860 84872 369912 84924
rect 77208 84804 77260 84856
rect 240784 84804 240836 84856
rect 272064 84804 272116 84856
rect 452660 84804 452712 84856
rect 276480 83580 276532 83632
rect 488540 83580 488592 83632
rect 160008 83512 160060 83564
rect 247500 83512 247552 83564
rect 278044 83512 278096 83564
rect 506480 83512 506532 83564
rect 135168 83444 135220 83496
rect 246396 83444 246448 83496
rect 279608 83444 279660 83496
rect 531320 83444 531372 83496
rect 184848 82084 184900 82136
rect 250444 82084 250496 82136
rect 272984 82084 273036 82136
rect 448612 82084 448664 82136
rect 234528 80860 234580 80912
rect 254400 80860 254452 80912
rect 261760 80860 261812 80912
rect 320180 80860 320232 80912
rect 155868 80792 155920 80844
rect 247408 80792 247460 80844
rect 264060 80792 264112 80844
rect 345020 80792 345072 80844
rect 131028 80724 131080 80776
rect 246304 80724 246356 80776
rect 264980 80724 265032 80776
rect 365720 80724 365772 80776
rect 73068 80656 73120 80708
rect 240692 80656 240744 80708
rect 267096 80656 267148 80708
rect 385040 80656 385092 80708
rect 275652 79296 275704 79348
rect 470600 79296 470652 79348
rect 286508 73108 286560 73160
rect 580172 73108 580224 73160
rect 2964 59168 3016 59220
rect 6276 59168 6328 59220
rect 2780 45500 2832 45552
rect 4896 45500 4948 45552
rect 286324 33056 286376 33108
rect 580172 33056 580224 33108
rect 311164 20612 311216 20664
rect 579988 20612 580040 20664
rect 2964 19456 3016 19508
rect 6184 19456 6236 19508
rect 340972 16532 341024 16584
rect 342168 16532 342220 16584
rect 448612 13268 448664 13320
rect 449808 13268 449860 13320
rect 193220 11704 193272 11756
rect 194416 11704 194468 11756
rect 209780 11704 209832 11756
rect 210976 11704 211028 11756
rect 235816 11704 235868 11756
rect 250536 11704 250588 11756
rect 271236 11704 271288 11756
rect 271512 11704 271564 11756
rect 284300 11704 284352 11756
rect 285404 11704 285456 11756
rect 316132 11704 316184 11756
rect 317328 11704 317380 11756
rect 423772 11704 423824 11756
rect 424968 11704 425020 11756
rect 262680 11636 262732 11688
rect 274824 11636 274876 11688
rect 262956 10752 263008 10804
rect 324320 10752 324372 10804
rect 262772 10684 262824 10736
rect 328736 10684 328788 10736
rect 263048 10616 263100 10668
rect 332692 10616 332744 10668
rect 262864 10548 262916 10600
rect 336280 10548 336332 10600
rect 267372 10480 267424 10532
rect 371240 10480 371292 10532
rect 267188 10412 267240 10464
rect 374000 10412 374052 10464
rect 267280 10344 267332 10396
rect 378416 10344 378468 10396
rect 267464 10276 267516 10328
rect 382372 10276 382424 10328
rect 283564 9596 283616 9648
rect 480536 9596 480588 9648
rect 283748 9528 283800 9580
rect 487620 9528 487672 9580
rect 285220 9460 285272 9512
rect 523040 9460 523092 9512
rect 285036 9392 285088 9444
rect 530124 9392 530176 9444
rect 281080 9324 281132 9376
rect 543188 9324 543240 9376
rect 280988 9256 281040 9308
rect 546684 9256 546736 9308
rect 282368 9188 282420 9240
rect 553768 9188 553820 9240
rect 253480 9120 253532 9172
rect 255964 9120 256016 9172
rect 282092 9120 282144 9172
rect 557356 9120 557408 9172
rect 282460 9052 282512 9104
rect 560852 9052 560904 9104
rect 282000 8984 282052 9036
rect 564440 8984 564492 9036
rect 283840 8916 283892 8968
rect 573916 8916 573968 8968
rect 252468 8848 252520 8900
rect 255872 8848 255924 8900
rect 272616 8848 272668 8900
rect 452108 8848 452160 8900
rect 272524 8780 272576 8832
rect 450912 8780 450964 8832
rect 273904 8712 273956 8764
rect 440332 8712 440384 8764
rect 270040 8644 270092 8696
rect 420184 8644 420236 8696
rect 270132 8576 270184 8628
rect 415492 8576 415544 8628
rect 268752 8508 268804 8560
rect 402520 8508 402572 8560
rect 269856 8440 269908 8492
rect 387156 8440 387208 8492
rect 268384 8372 268436 8424
rect 379980 8372 380032 8424
rect 271604 8304 271656 8356
rect 365812 8304 365864 8356
rect 109316 8236 109368 8288
rect 242256 8236 242308 8288
rect 276572 8236 276624 8288
rect 493508 8236 493560 8288
rect 98644 8168 98696 8220
rect 234344 8168 234396 8220
rect 276020 8168 276072 8220
rect 497096 8168 497148 8220
rect 102232 8100 102284 8152
rect 242164 8100 242216 8152
rect 277032 8100 277084 8152
rect 500592 8100 500644 8152
rect 77392 8032 77444 8084
rect 240508 8032 240560 8084
rect 278412 8032 278464 8084
rect 504180 8032 504232 8084
rect 73804 7964 73856 8016
rect 240416 7964 240468 8016
rect 278320 7964 278372 8016
rect 507676 7964 507728 8016
rect 70216 7896 70268 7948
rect 240600 7896 240652 7948
rect 278228 7896 278280 7948
rect 511264 7896 511316 7948
rect 66720 7828 66772 7880
rect 241244 7828 241296 7880
rect 278136 7828 278188 7880
rect 514760 7828 514812 7880
rect 63224 7760 63276 7812
rect 240324 7760 240376 7812
rect 277584 7760 277636 7812
rect 518348 7760 518400 7812
rect 59636 7692 59688 7744
rect 239036 7692 239088 7744
rect 279700 7692 279752 7744
rect 521844 7692 521896 7744
rect 21824 7624 21876 7676
rect 235356 7624 235408 7676
rect 279792 7624 279844 7676
rect 525432 7624 525484 7676
rect 13544 7556 13596 7608
rect 235264 7556 235316 7608
rect 278780 7556 278832 7608
rect 529020 7556 529072 7608
rect 105728 7488 105780 7540
rect 234160 7488 234212 7540
rect 276756 7488 276808 7540
rect 489920 7488 489972 7540
rect 116400 7420 116452 7472
rect 244648 7420 244700 7472
rect 276940 7420 276992 7472
rect 486424 7420 486476 7472
rect 112812 7352 112864 7404
rect 234252 7352 234304 7404
rect 275100 7352 275152 7404
rect 482836 7352 482888 7404
rect 119896 7284 119948 7336
rect 234068 7284 234120 7336
rect 275192 7284 275244 7336
rect 478144 7284 478196 7336
rect 275744 7216 275796 7268
rect 474556 7216 474608 7268
rect 274364 7148 274416 7200
rect 467472 7148 467524 7200
rect 273628 7080 273680 7132
rect 463976 7080 464028 7132
rect 273720 7012 273772 7064
rect 460388 7012 460440 7064
rect 270500 6944 270552 6996
rect 432052 6944 432104 6996
rect 160100 6808 160152 6860
rect 249064 6808 249116 6860
rect 260380 6808 260432 6860
rect 294880 6808 294932 6860
rect 295984 6808 296036 6860
rect 580172 6808 580224 6860
rect 156604 6740 156656 6792
rect 247316 6740 247368 6792
rect 264612 6740 264664 6792
rect 354036 6740 354088 6792
rect 153016 6672 153068 6724
rect 247224 6672 247276 6724
rect 265532 6672 265584 6724
rect 357532 6672 357584 6724
rect 149520 6604 149572 6656
rect 247776 6604 247828 6656
rect 265716 6604 265768 6656
rect 361120 6604 361172 6656
rect 145932 6536 145984 6588
rect 247592 6536 247644 6588
rect 265992 6536 266044 6588
rect 364616 6536 364668 6588
rect 2780 6468 2832 6520
rect 4804 6468 4856 6520
rect 142436 6468 142488 6520
rect 246028 6468 246080 6520
rect 266084 6468 266136 6520
rect 368204 6468 368256 6520
rect 138848 6400 138900 6452
rect 246212 6400 246264 6452
rect 266728 6400 266780 6452
rect 374092 6400 374144 6452
rect 135260 6332 135312 6384
rect 246120 6332 246172 6384
rect 266636 6332 266688 6384
rect 377680 6332 377732 6384
rect 122288 6264 122340 6316
rect 244464 6264 244516 6316
rect 267740 6264 267792 6316
rect 393044 6264 393096 6316
rect 118792 6196 118844 6248
rect 244556 6196 244608 6248
rect 267924 6196 267976 6248
rect 396540 6196 396592 6248
rect 44272 6128 44324 6180
rect 238116 6128 238168 6180
rect 268844 6128 268896 6180
rect 400128 6128 400180 6180
rect 188528 6060 188580 6112
rect 250260 6060 250312 6112
rect 264428 6060 264480 6112
rect 350448 6060 350500 6112
rect 192024 5992 192076 6044
rect 250352 5992 250404 6044
rect 264704 5992 264756 6044
rect 346952 5992 347004 6044
rect 206192 5924 206244 5976
rect 251548 5924 251600 5976
rect 264520 5924 264572 5976
rect 343364 5924 343416 5976
rect 213368 5856 213420 5908
rect 252928 5856 252980 5908
rect 263416 5856 263468 5908
rect 338672 5856 338724 5908
rect 216864 5788 216916 5840
rect 252836 5788 252888 5840
rect 263324 5788 263376 5840
rect 335084 5788 335136 5840
rect 220452 5720 220504 5772
rect 252744 5720 252796 5772
rect 262588 5720 262640 5772
rect 331588 5720 331640 5772
rect 223948 5652 224000 5704
rect 253664 5652 253716 5704
rect 263140 5652 263192 5704
rect 328000 5652 328052 5704
rect 227536 5584 227588 5636
rect 254308 5584 254360 5636
rect 262312 5584 262364 5636
rect 324412 5584 324464 5636
rect 231032 5516 231084 5568
rect 254216 5516 254268 5568
rect 260840 5516 260892 5568
rect 322112 5516 322164 5568
rect 177948 5448 178000 5500
rect 249984 5448 250036 5500
rect 259828 5448 259880 5500
rect 290188 5448 290240 5500
rect 174268 5380 174320 5432
rect 248696 5380 248748 5432
rect 260472 5380 260524 5432
rect 293132 5448 293184 5500
rect 293224 5448 293276 5500
rect 290556 5380 290608 5432
rect 465172 5448 465224 5500
rect 475752 5380 475804 5432
rect 173164 5312 173216 5364
rect 249616 5312 249668 5364
rect 257344 5312 257396 5364
rect 264152 5312 264204 5364
rect 277216 5312 277268 5364
rect 492312 5312 492364 5364
rect 170772 5244 170824 5296
rect 248788 5244 248840 5296
rect 257620 5244 257672 5296
rect 267740 5244 267792 5296
rect 276112 5244 276164 5296
rect 495900 5244 495952 5296
rect 169668 5176 169720 5228
rect 248972 5176 249024 5228
rect 257528 5176 257580 5228
rect 268844 5176 268896 5228
rect 277124 5176 277176 5228
rect 499396 5176 499448 5228
rect 167184 5108 167236 5160
rect 248880 5108 248932 5160
rect 257436 5108 257488 5160
rect 271236 5108 271288 5160
rect 277768 5108 277820 5160
rect 510068 5108 510120 5160
rect 166080 5040 166132 5092
rect 248604 5040 248656 5092
rect 257712 5040 257764 5092
rect 272432 5040 272484 5092
rect 278964 5040 279016 5092
rect 163688 4972 163740 5024
rect 249432 4972 249484 5024
rect 259092 4972 259144 5024
rect 276020 4972 276072 5024
rect 277400 4972 277452 5024
rect 141240 4904 141292 4956
rect 245936 4904 245988 4956
rect 246396 4904 246448 4956
rect 255688 4904 255740 4956
rect 258908 4904 258960 4956
rect 278320 4904 278372 4956
rect 278504 4972 278556 5024
rect 12348 4836 12400 4888
rect 235632 4836 235684 4888
rect 242900 4836 242952 4888
rect 255780 4836 255832 4888
rect 259184 4836 259236 4888
rect 279516 4836 279568 4888
rect 280252 4904 280304 4956
rect 513564 5040 513616 5092
rect 517152 4972 517204 5024
rect 281816 4836 281868 4888
rect 534908 4904 534960 4956
rect 7656 4768 7708 4820
rect 234436 4768 234488 4820
rect 234620 4768 234672 4820
rect 254124 4768 254176 4820
rect 258356 4768 258408 4820
rect 281908 4768 281960 4820
rect 545488 4836 545540 4888
rect 556160 4768 556212 4820
rect 181444 4700 181496 4752
rect 250628 4700 250680 4752
rect 259000 4700 259052 4752
rect 283104 4700 283156 4752
rect 291936 4700 291988 4752
rect 293132 4700 293184 4752
rect 293684 4700 293736 4752
rect 458088 4700 458140 4752
rect 184940 4632 184992 4684
rect 250720 4632 250772 4684
rect 264796 4632 264848 4684
rect 352840 4632 352892 4684
rect 187332 4564 187384 4616
rect 250168 4564 250220 4616
rect 263784 4564 263836 4616
rect 339868 4564 339920 4616
rect 190828 4496 190880 4548
rect 250076 4496 250128 4548
rect 261944 4496 261996 4548
rect 318524 4496 318576 4548
rect 194416 4428 194468 4480
rect 251456 4428 251508 4480
rect 261116 4428 261168 4480
rect 315028 4428 315080 4480
rect 197912 4360 197964 4412
rect 252284 4360 252336 4412
rect 261576 4360 261628 4412
rect 311440 4360 311492 4412
rect 201500 4292 201552 4344
rect 251364 4292 251416 4344
rect 259644 4292 259696 4344
rect 304356 4292 304408 4344
rect 205088 4224 205140 4276
rect 252192 4224 252244 4276
rect 259460 4224 259512 4276
rect 300768 4224 300820 4276
rect 218060 4156 218112 4208
rect 219348 4156 219400 4208
rect 222752 4156 222804 4208
rect 226248 4156 226300 4208
rect 226340 4156 226392 4208
rect 227628 4156 227680 4208
rect 227720 4156 227772 4208
rect 253388 4156 253440 4208
rect 260564 4156 260616 4208
rect 297272 4156 297324 4208
rect 440240 4156 440292 4208
rect 441528 4156 441580 4208
rect 57244 4088 57296 4140
rect 60832 4020 60884 4072
rect 61936 4020 61988 4072
rect 69112 4088 69164 4140
rect 70308 4088 70360 4140
rect 71504 4088 71556 4140
rect 234068 4088 234120 4140
rect 238392 4088 238444 4140
rect 284852 4088 284904 4140
rect 299664 4088 299716 4140
rect 300124 4088 300176 4140
rect 433248 4088 433300 4140
rect 434168 4088 434220 4140
rect 508872 4088 508924 4140
rect 239312 4020 239364 4072
rect 290464 4020 290516 4072
rect 422576 4020 422628 4072
rect 422944 4020 422996 4072
rect 50160 3952 50212 4004
rect 238024 3952 238076 4004
rect 289452 3952 289504 4004
rect 296168 3952 296220 4004
rect 429660 3952 429712 4004
rect 433984 4020 434036 4072
rect 512460 4020 512512 4072
rect 439136 3952 439188 4004
rect 439504 3952 439556 4004
rect 519544 3952 519596 4004
rect 46664 3884 46716 3936
rect 238852 3884 238904 3936
rect 291844 3884 291896 3936
rect 426164 3884 426216 3936
rect 434076 3884 434128 3936
rect 515956 3884 516008 3936
rect 45468 3816 45520 3868
rect 238208 3816 238260 3868
rect 269580 3816 269632 3868
rect 408408 3816 408460 3868
rect 408500 3816 408552 3868
rect 533712 3816 533764 3868
rect 39580 3748 39632 3800
rect 237472 3748 237524 3800
rect 247592 3748 247644 3800
rect 255504 3748 255556 3800
rect 289544 3748 289596 3800
rect 447416 3748 447468 3800
rect 38384 3680 38436 3732
rect 237656 3680 237708 3732
rect 242716 3680 242768 3732
rect 244096 3680 244148 3732
rect 251916 3680 251968 3732
rect 280804 3680 280856 3732
rect 443828 3680 443880 3732
rect 32404 3612 32456 3664
rect 237564 3612 237616 3664
rect 241704 3612 241756 3664
rect 252008 3612 252060 3664
rect 254676 3612 254728 3664
rect 258540 3612 258592 3664
rect 27712 3544 27764 3596
rect 28816 3544 28868 3596
rect 31300 3544 31352 3596
rect 232044 3544 232096 3596
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 19432 3476 19484 3528
rect 20628 3476 20680 3528
rect 24216 3476 24268 3528
rect 236460 3544 236512 3596
rect 232228 3476 232280 3528
rect 233148 3476 233200 3528
rect 233424 3476 233476 3528
rect 234528 3476 234580 3528
rect 238116 3476 238168 3528
rect 14740 3408 14792 3460
rect 237104 3408 237156 3460
rect 240508 3544 240560 3596
rect 257896 3544 257948 3596
rect 260656 3544 260708 3596
rect 290648 3612 290700 3664
rect 280712 3544 280764 3596
rect 287704 3544 287756 3596
rect 288992 3544 289044 3596
rect 289360 3544 289412 3596
rect 296076 3544 296128 3596
rect 454500 3612 454552 3664
rect 461584 3544 461636 3596
rect 244372 3476 244424 3528
rect 245200 3476 245252 3528
rect 254676 3476 254728 3528
rect 255412 3476 255464 3528
rect 257804 3476 257856 3528
rect 259460 3476 259512 3528
rect 260104 3476 260156 3528
rect 261760 3476 261812 3528
rect 276664 3476 276716 3528
rect 468668 3476 468720 3528
rect 254860 3408 254912 3460
rect 257160 3408 257212 3460
rect 265348 3408 265400 3460
rect 271144 3408 271196 3460
rect 316224 3408 316276 3460
rect 319444 3408 319496 3460
rect 583392 3408 583444 3460
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 35992 3340 36044 3392
rect 37188 3340 37240 3392
rect 41880 3340 41932 3392
rect 42708 3340 42760 3392
rect 43076 3340 43128 3392
rect 44088 3340 44140 3392
rect 48964 3340 49016 3392
rect 49608 3340 49660 3392
rect 51356 3340 51408 3392
rect 52368 3340 52420 3392
rect 52552 3340 52604 3392
rect 53656 3340 53708 3392
rect 58440 3340 58492 3392
rect 59268 3340 59320 3392
rect 64328 3340 64380 3392
rect 64788 3340 64840 3392
rect 65524 3340 65576 3392
rect 66168 3340 66220 3392
rect 67916 3340 67968 3392
rect 68928 3340 68980 3392
rect 72608 3340 72660 3392
rect 73068 3340 73120 3392
rect 75000 3340 75052 3392
rect 75828 3340 75880 3392
rect 76196 3340 76248 3392
rect 77208 3340 77260 3392
rect 80888 3340 80940 3392
rect 81348 3340 81400 3392
rect 82084 3340 82136 3392
rect 82728 3340 82780 3392
rect 83280 3340 83332 3392
rect 84108 3340 84160 3392
rect 84476 3340 84528 3392
rect 85488 3340 85540 3392
rect 85672 3340 85724 3392
rect 86684 3340 86736 3392
rect 91560 3340 91612 3392
rect 92388 3340 92440 3392
rect 6460 3272 6512 3324
rect 7564 3272 7616 3324
rect 78588 3272 78640 3324
rect 92756 3272 92808 3324
rect 93768 3272 93820 3324
rect 97448 3272 97500 3324
rect 97908 3272 97960 3324
rect 99840 3272 99892 3324
rect 100668 3272 100720 3324
rect 101036 3272 101088 3324
rect 102048 3272 102100 3324
rect 242624 3340 242676 3392
rect 251180 3340 251232 3392
rect 256424 3340 256476 3392
rect 268200 3340 268252 3392
rect 401324 3340 401376 3392
rect 403624 3340 403676 3392
rect 526628 3340 526680 3392
rect 89168 3204 89220 3256
rect 239312 3272 239364 3324
rect 244924 3272 244976 3324
rect 264244 3272 264296 3324
rect 270040 3272 270092 3324
rect 271512 3272 271564 3324
rect 305552 3272 305604 3324
rect 307760 3272 307812 3324
rect 309048 3272 309100 3324
rect 309140 3272 309192 3324
rect 436744 3272 436796 3324
rect 439596 3272 439648 3324
rect 448612 3272 448664 3324
rect 96252 3136 96304 3188
rect 243912 3204 243964 3256
rect 280896 3204 280948 3256
rect 394240 3204 394292 3256
rect 396724 3204 396776 3256
rect 498200 3204 498252 3256
rect 103336 3136 103388 3188
rect 243452 3136 243504 3188
rect 271420 3136 271472 3188
rect 273628 3136 273680 3188
rect 289268 3136 289320 3188
rect 390652 3136 390704 3188
rect 393964 3136 394016 3188
rect 494704 3136 494756 3188
rect 106924 3068 106976 3120
rect 107568 3068 107620 3120
rect 108120 3068 108172 3120
rect 108948 3068 109000 3120
rect 110512 3068 110564 3120
rect 243084 3068 243136 3120
rect 269764 3068 269816 3120
rect 340972 3068 341024 3120
rect 357440 3068 357492 3120
rect 358728 3068 358780 3120
rect 365720 3068 365772 3120
rect 367008 3068 367060 3120
rect 374000 3068 374052 3120
rect 375288 3068 375340 3120
rect 382280 3068 382332 3120
rect 383568 3068 383620 3120
rect 400864 3068 400916 3120
rect 501788 3068 501840 3120
rect 114008 3000 114060 3052
rect 114468 3000 114520 3052
rect 115204 3000 115256 3052
rect 115848 3000 115900 3052
rect 123484 3000 123536 3052
rect 124128 3000 124180 3052
rect 124680 3000 124732 3052
rect 125508 3000 125560 3052
rect 125876 3000 125928 3052
rect 126888 3000 126940 3052
rect 126980 3000 127032 3052
rect 128268 3000 128320 3052
rect 245292 3000 245344 3052
rect 249984 3000 250036 3052
rect 252468 3000 252520 3052
rect 271328 3000 271380 3052
rect 277124 3000 277176 3052
rect 289084 3000 289136 3052
rect 351644 3000 351696 3052
rect 391204 3000 391256 3052
rect 491116 3000 491168 3052
rect 121092 2932 121144 2984
rect 245384 2932 245436 2984
rect 117596 2864 117648 2916
rect 130568 2864 130620 2916
rect 131028 2864 131080 2916
rect 132960 2864 133012 2916
rect 133788 2864 133840 2916
rect 134156 2864 134208 2916
rect 135168 2864 135220 2916
rect 140044 2864 140096 2916
rect 140688 2864 140740 2916
rect 143540 2864 143592 2916
rect 144828 2864 144880 2916
rect 147128 2864 147180 2916
rect 147588 2864 147640 2916
rect 148324 2864 148376 2916
rect 148968 2864 149020 2916
rect 150624 2864 150676 2916
rect 151728 2864 151780 2916
rect 151820 2864 151872 2916
rect 153108 2864 153160 2916
rect 155408 2864 155460 2916
rect 155868 2864 155920 2916
rect 157800 2864 157852 2916
rect 158628 2864 158680 2916
rect 158904 2864 158956 2916
rect 160008 2864 160060 2916
rect 164884 2864 164936 2916
rect 165528 2864 165580 2916
rect 168380 2864 168432 2916
rect 169576 2864 169628 2916
rect 171968 2864 172020 2916
rect 175464 2796 175516 2848
rect 176660 2864 176712 2916
rect 177856 2864 177908 2916
rect 233976 2864 234028 2916
rect 237012 2864 237064 2916
rect 253204 2932 253256 2984
rect 289176 2932 289228 2984
rect 344560 2932 344612 2984
rect 415400 2932 415452 2984
rect 416688 2932 416740 2984
rect 417516 2932 417568 2984
rect 469864 2932 469916 2984
rect 248788 2864 248840 2916
rect 253296 2864 253348 2916
rect 286416 2864 286468 2916
rect 337476 2864 337528 2916
rect 409236 2864 409288 2916
rect 455696 2864 455748 2916
rect 233792 2796 233844 2848
rect 241060 2796 241112 2848
rect 282184 2796 282236 2848
rect 323308 2796 323360 2848
rect 324320 2796 324372 2848
rect 325608 2796 325660 2848
rect 332600 2796 332652 2848
rect 333888 2796 333940 2848
rect 414664 2796 414716 2848
rect 459192 2796 459244 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 8128 700466 8156 703520
rect 24320 700534 24348 703520
rect 40512 700602 40540 703520
rect 72988 700806 73016 703520
rect 89180 700874 89208 703520
rect 105464 701010 105492 703520
rect 105452 701004 105504 701010
rect 105452 700946 105504 700952
rect 89168 700868 89220 700874
rect 89168 700810 89220 700816
rect 72976 700800 73028 700806
rect 72976 700742 73028 700748
rect 40500 700596 40552 700602
rect 40500 700538 40552 700544
rect 24308 700528 24360 700534
rect 24308 700470 24360 700476
rect 8116 700460 8168 700466
rect 8116 700402 8168 700408
rect 137848 700126 137876 703520
rect 137836 700120 137888 700126
rect 137836 700062 137888 700068
rect 154132 700058 154160 703520
rect 154120 700052 154172 700058
rect 154120 699994 154172 700000
rect 170324 699990 170352 703520
rect 170312 699984 170364 699990
rect 170312 699926 170364 699932
rect 202800 699786 202828 703520
rect 202788 699780 202840 699786
rect 202788 699722 202840 699728
rect 218992 699718 219020 703520
rect 235184 699854 235212 703520
rect 262220 701004 262272 701010
rect 262220 700946 262272 700952
rect 256516 700936 256568 700942
rect 256516 700878 256568 700884
rect 256424 700732 256476 700738
rect 256424 700674 256476 700680
rect 255136 700392 255188 700398
rect 255136 700334 255188 700340
rect 255044 700324 255096 700330
rect 255044 700266 255096 700272
rect 235172 699848 235224 699854
rect 235172 699790 235224 699796
rect 235908 699848 235960 699854
rect 235908 699790 235960 699796
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 670818 3464 671191
rect 3424 670812 3476 670818
rect 3424 670754 3476 670760
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 235920 391542 235948 699790
rect 253572 696992 253624 696998
rect 253572 696934 253624 696940
rect 252468 643136 252520 643142
rect 252468 643078 252520 643084
rect 252376 630692 252428 630698
rect 252376 630634 252428 630640
rect 252284 616888 252336 616894
rect 252284 616830 252336 616836
rect 251088 590708 251140 590714
rect 251088 590650 251140 590656
rect 250996 576904 251048 576910
rect 250996 576846 251048 576852
rect 250904 563100 250956 563106
rect 250904 563042 250956 563048
rect 249708 536852 249760 536858
rect 249708 536794 249760 536800
rect 249616 524476 249668 524482
rect 249616 524418 249668 524424
rect 249524 510672 249576 510678
rect 249524 510614 249576 510620
rect 248328 484424 248380 484430
rect 248328 484366 248380 484372
rect 248236 456816 248288 456822
rect 248236 456758 248288 456764
rect 246948 430636 247000 430642
rect 246948 430578 247000 430584
rect 246856 404388 246908 404394
rect 246856 404330 246908 404336
rect 246868 393314 246896 404330
rect 246684 393286 246896 393314
rect 235908 391536 235960 391542
rect 235908 391478 235960 391484
rect 242072 390516 242124 390522
rect 242072 390458 242124 390464
rect 240048 390312 240100 390318
rect 240048 390254 240100 390260
rect 238668 390108 238720 390114
rect 238668 390050 238720 390056
rect 4712 389972 4764 389978
rect 4712 389914 4764 389920
rect 3332 389088 3384 389094
rect 3332 389030 3384 389036
rect 3344 371385 3372 389030
rect 4068 389020 4120 389026
rect 4068 388962 4120 388968
rect 3976 388748 4028 388754
rect 3976 388690 4028 388696
rect 3884 388612 3936 388618
rect 3884 388554 3936 388560
rect 3792 388544 3844 388550
rect 3792 388486 3844 388492
rect 3700 388476 3752 388482
rect 3700 388418 3752 388424
rect 3608 388408 3660 388414
rect 3608 388350 3660 388356
rect 3516 388340 3568 388346
rect 3516 388282 3568 388288
rect 3422 387968 3478 387977
rect 3422 387903 3478 387912
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 2780 358488 2832 358494
rect 2778 358456 2780 358465
rect 2832 358456 2834 358465
rect 2778 358391 2834 358400
rect 2780 345908 2832 345914
rect 2780 345850 2832 345856
rect 2792 345409 2820 345850
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 2686 333432 2742 333441
rect 2686 333367 2742 333376
rect 18 333296 74 333305
rect 18 333231 74 333240
rect 32 16574 60 333231
rect 32 16546 152 16574
rect 124 490 152 16546
rect 2700 3534 2728 333367
rect 3332 306264 3384 306270
rect 3330 306232 3332 306241
rect 3384 306232 3386 306241
rect 3330 306167 3386 306176
rect 2780 254652 2832 254658
rect 2780 254594 2832 254600
rect 2792 254153 2820 254594
rect 2778 254144 2834 254153
rect 2778 254079 2834 254088
rect 2780 241392 2832 241398
rect 2780 241334 2832 241340
rect 2792 241097 2820 241334
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 2964 202836 3016 202842
rect 2964 202778 3016 202784
rect 2976 201929 3004 202778
rect 2962 201920 3018 201929
rect 2962 201855 3018 201864
rect 2780 188964 2832 188970
rect 2780 188906 2832 188912
rect 2792 188873 2820 188906
rect 2778 188864 2834 188873
rect 2778 188799 2834 188808
rect 3148 150408 3200 150414
rect 3148 150350 3200 150356
rect 3160 149841 3188 150350
rect 3146 149832 3202 149841
rect 3146 149767 3202 149776
rect 2780 137284 2832 137290
rect 2780 137226 2832 137232
rect 2792 136785 2820 137226
rect 2778 136776 2834 136785
rect 2778 136711 2834 136720
rect 3240 97912 3292 97918
rect 3240 97854 3292 97860
rect 3252 97617 3280 97854
rect 3238 97608 3294 97617
rect 3238 97543 3294 97552
rect 2780 85264 2832 85270
rect 2780 85206 2832 85212
rect 2792 84697 2820 85206
rect 2778 84688 2834 84697
rect 2778 84623 2834 84632
rect 2964 59220 3016 59226
rect 2964 59162 3016 59168
rect 2976 58585 3004 59162
rect 2962 58576 3018 58585
rect 2962 58511 3018 58520
rect 2780 45552 2832 45558
rect 2778 45520 2780 45529
rect 2832 45520 2834 45529
rect 2778 45455 2834 45464
rect 3436 32473 3464 387903
rect 3528 71641 3556 388282
rect 3620 110673 3648 388350
rect 3712 162897 3740 388418
rect 3804 214985 3832 388486
rect 3896 267209 3924 388554
rect 3988 293185 4016 388690
rect 4080 319297 4108 388962
rect 4724 358494 4752 389914
rect 5356 389904 5408 389910
rect 5356 389846 5408 389852
rect 5172 389768 5224 389774
rect 5172 389710 5224 389716
rect 5080 389632 5132 389638
rect 5080 389574 5132 389580
rect 4988 389496 5040 389502
rect 4988 389438 5040 389444
rect 4896 389360 4948 389366
rect 4802 389328 4858 389337
rect 4896 389302 4948 389308
rect 4802 389263 4858 389272
rect 4712 358488 4764 358494
rect 4712 358430 4764 358436
rect 4066 319288 4122 319297
rect 4066 319223 4122 319232
rect 3974 293176 4030 293185
rect 3974 293111 4030 293120
rect 3882 267200 3938 267209
rect 3882 267135 3938 267144
rect 3790 214976 3846 214985
rect 3790 214911 3846 214920
rect 4068 177336 4120 177342
rect 4068 177278 4120 177284
rect 3698 162888 3754 162897
rect 3698 162823 3754 162832
rect 3606 110664 3662 110673
rect 3606 110599 3662 110608
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 2976 19417 3004 19450
rect 2962 19408 3018 19417
rect 2962 19343 3018 19352
rect 2780 6520 2832 6526
rect 2778 6488 2780 6497
rect 2832 6488 2834 6497
rect 2778 6423 2834 6432
rect 2870 4856 2926 4865
rect 2870 4791 2926 4800
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 400 598 612 626
rect 400 490 428 598
rect 124 462 428 490
rect 584 480 612 598
rect 1688 480 1716 3470
rect 2884 480 2912 4791
rect 4080 480 4108 177278
rect 4816 6526 4844 389263
rect 4908 45558 4936 389302
rect 5000 85270 5028 389438
rect 5092 137290 5120 389574
rect 5184 188970 5212 389710
rect 5264 388680 5316 388686
rect 5264 388622 5316 388628
rect 5276 241398 5304 388622
rect 5368 254658 5396 389846
rect 6552 389836 6604 389842
rect 6552 389778 6604 389784
rect 6460 389700 6512 389706
rect 6460 389642 6512 389648
rect 6368 389564 6420 389570
rect 6368 389506 6420 389512
rect 6182 389464 6238 389473
rect 6182 389399 6238 389408
rect 6276 389428 6328 389434
rect 5448 389156 5500 389162
rect 5448 389098 5500 389104
rect 5460 345914 5488 389098
rect 5448 345908 5500 345914
rect 5448 345850 5500 345856
rect 5448 336048 5500 336054
rect 5448 335990 5500 335996
rect 5356 254652 5408 254658
rect 5356 254594 5408 254600
rect 5264 241392 5316 241398
rect 5264 241334 5316 241340
rect 5172 188964 5224 188970
rect 5172 188906 5224 188912
rect 5080 137284 5132 137290
rect 5080 137226 5132 137232
rect 4988 85264 5040 85270
rect 4988 85206 5040 85212
rect 4896 45552 4948 45558
rect 4896 45494 4948 45500
rect 5460 6914 5488 335990
rect 6196 19514 6224 389399
rect 6276 389370 6328 389376
rect 6288 59226 6316 389370
rect 6380 97918 6408 389506
rect 6472 150414 6500 389642
rect 6564 202842 6592 389778
rect 236274 389600 236330 389609
rect 236274 389535 236330 389544
rect 6644 389224 6696 389230
rect 6644 389166 6696 389172
rect 6656 306270 6684 389166
rect 235584 388104 235640 388113
rect 235584 388039 235640 388048
rect 235598 387940 235626 388039
rect 236288 387954 236316 389535
rect 237194 389192 237250 389201
rect 237194 389127 237250 389136
rect 236872 388240 236928 388249
rect 236872 388175 236928 388184
rect 236072 387926 236316 387954
rect 236886 387940 236914 388175
rect 236736 387864 236788 387870
rect 234908 387790 235244 387818
rect 236440 387812 236736 387818
rect 236440 387806 236788 387812
rect 237208 387818 237236 389127
rect 237930 388376 237986 388385
rect 237930 388311 237986 388320
rect 237944 387954 237972 388311
rect 237728 387926 237972 387954
rect 238392 387864 238444 387870
rect 236440 387790 236776 387806
rect 237208 387790 237268 387818
rect 238096 387812 238392 387818
rect 238680 387818 238708 390050
rect 239588 388884 239640 388890
rect 239588 388826 239640 388832
rect 239220 388816 239272 388822
rect 239220 388758 239272 388764
rect 239232 387954 239260 388758
rect 239600 387954 239628 388826
rect 240060 387954 240088 390254
rect 241152 390040 241204 390046
rect 241152 389982 241204 389988
rect 240416 388000 240468 388006
rect 238924 387926 239260 387954
rect 239384 387926 239628 387954
rect 239752 387926 240088 387954
rect 240212 387948 240416 387954
rect 241164 387954 241192 389982
rect 240212 387942 240468 387948
rect 240212 387926 240456 387942
rect 240580 387938 240916 387954
rect 240580 387932 240928 387938
rect 240580 387926 240876 387932
rect 241040 387926 241192 387954
rect 241244 388000 241296 388006
rect 242084 387954 242112 390458
rect 246304 390448 246356 390454
rect 246304 390390 246356 390396
rect 245016 390380 245068 390386
rect 245016 390322 245068 390328
rect 243820 390244 243872 390250
rect 243820 390186 243872 390192
rect 242532 390176 242584 390182
rect 242532 390118 242584 390124
rect 242544 387954 242572 390118
rect 243360 389292 243412 389298
rect 243360 389234 243412 389240
rect 242808 388068 242860 388074
rect 242808 388010 242860 388016
rect 242820 387954 242848 388010
rect 243372 387954 243400 389234
rect 243832 387954 243860 390186
rect 244326 388204 244378 388210
rect 244326 388146 244378 388152
rect 243958 388136 244010 388142
rect 243958 388078 244010 388084
rect 241296 387948 241408 387954
rect 241244 387942 241408 387948
rect 241256 387926 241408 387942
rect 241868 387926 242112 387954
rect 242236 387926 242572 387954
rect 242696 387926 242848 387954
rect 243064 387926 243400 387954
rect 243524 387926 243860 387954
rect 243970 387940 243998 388078
rect 244338 387940 244366 388146
rect 245028 387954 245056 390322
rect 245476 388952 245528 388958
rect 245476 388894 245528 388900
rect 245488 387954 245516 388894
rect 245568 388272 245620 388278
rect 245568 388214 245620 388220
rect 244812 387926 245056 387954
rect 245180 387926 245516 387954
rect 245580 387954 245608 388214
rect 246316 387954 246344 390390
rect 246684 387954 246712 393286
rect 246960 387954 246988 430578
rect 248144 418192 248196 418198
rect 248144 418134 248196 418140
rect 248156 390318 248184 418134
rect 247500 390312 247552 390318
rect 247500 390254 247552 390260
rect 248144 390312 248196 390318
rect 248144 390254 248196 390260
rect 247512 387954 247540 390254
rect 248248 389174 248276 456758
rect 247972 389146 248276 389174
rect 247972 387954 248000 389146
rect 248340 387954 248368 484366
rect 249432 470620 249484 470626
rect 249432 470562 249484 470568
rect 249340 390584 249392 390590
rect 249340 390526 249392 390532
rect 248972 390312 249024 390318
rect 248972 390254 249024 390260
rect 248984 389174 249012 390254
rect 248800 389146 249012 389174
rect 248800 387954 248828 389146
rect 249352 388226 249380 390526
rect 249444 390318 249472 470562
rect 249432 390312 249484 390318
rect 249432 390254 249484 390260
rect 249156 388204 249208 388210
rect 249156 388146 249208 388152
rect 249306 388198 249380 388226
rect 249536 388210 249564 510614
rect 249524 388204 249576 388210
rect 249168 387954 249196 388146
rect 245580 387926 245640 387954
rect 246008 387926 246344 387954
rect 246468 387926 246712 387954
rect 246836 387926 246988 387954
rect 247296 387926 247540 387954
rect 247664 387926 248000 387954
rect 248124 387926 248368 387954
rect 248492 387926 248828 387954
rect 248952 387926 249196 387954
rect 249306 387940 249334 388198
rect 249524 388146 249576 388152
rect 249628 387954 249656 524418
rect 249720 390590 249748 536794
rect 249708 390584 249760 390590
rect 249708 390526 249760 390532
rect 250812 390584 250864 390590
rect 250812 390526 250864 390532
rect 250444 390312 250496 390318
rect 250444 390254 250496 390260
rect 250456 387954 250484 390254
rect 250824 387954 250852 390526
rect 250916 390318 250944 563042
rect 250904 390312 250956 390318
rect 250904 390254 250956 390260
rect 251008 388226 251036 576846
rect 251100 390590 251128 590650
rect 252296 393314 252324 616830
rect 251744 393286 252324 393314
rect 251088 390584 251140 390590
rect 251088 390526 251140 390532
rect 249628 387926 249780 387954
rect 250148 387926 250484 387954
rect 250608 387926 250852 387954
rect 250962 388198 251036 388226
rect 250962 387940 250990 388198
rect 251744 387954 251772 393286
rect 252100 390312 252152 390318
rect 252100 390254 252152 390260
rect 252112 387954 252140 390254
rect 252388 387954 252416 630634
rect 252480 390318 252508 643078
rect 253584 393314 253612 696934
rect 253756 683188 253808 683194
rect 253756 683130 253808 683136
rect 253664 670744 253716 670750
rect 253664 670686 253716 670692
rect 253400 393286 253612 393314
rect 252468 390312 252520 390318
rect 252468 390254 252520 390260
rect 252928 390312 252980 390318
rect 252928 390254 252980 390260
rect 252940 387954 252968 390254
rect 253400 387954 253428 393286
rect 253676 390318 253704 670686
rect 253664 390312 253716 390318
rect 253664 390254 253716 390260
rect 253768 387954 253796 683130
rect 253848 391264 253900 391270
rect 253848 391206 253900 391212
rect 251436 387926 251772 387954
rect 251896 387926 252140 387954
rect 252264 387926 252416 387954
rect 252724 387926 252968 387954
rect 253092 387926 253428 387954
rect 253552 387926 253796 387954
rect 253860 387954 253888 391206
rect 254584 390312 254636 390318
rect 254584 390254 254636 390260
rect 254596 387954 254624 390254
rect 255056 387954 255084 700266
rect 255148 390318 255176 700334
rect 256436 393314 256464 700674
rect 255884 393286 256464 393314
rect 255228 391332 255280 391338
rect 255228 391274 255280 391280
rect 255136 390312 255188 390318
rect 255136 390254 255188 390260
rect 255240 388226 255268 391274
rect 253860 387926 253920 387954
rect 254380 387926 254624 387954
rect 254748 387926 255084 387954
rect 255194 388198 255268 388226
rect 255194 387940 255222 388198
rect 255884 387954 255912 393286
rect 256240 390312 256292 390318
rect 256240 390254 256292 390260
rect 256252 387954 256280 390254
rect 256528 387954 256556 700878
rect 256608 700664 256660 700670
rect 256608 700606 256660 700612
rect 256620 390318 256648 700606
rect 257712 700256 257764 700262
rect 257712 700198 257764 700204
rect 257724 393314 257752 700198
rect 257804 700188 257856 700194
rect 257804 700130 257856 700136
rect 257540 393286 257752 393314
rect 256608 390312 256660 390318
rect 256608 390254 256660 390260
rect 257068 390312 257120 390318
rect 257068 390254 257120 390260
rect 257080 387954 257108 390254
rect 257540 387954 257568 393286
rect 257816 390318 257844 700130
rect 260932 700120 260984 700126
rect 260932 700062 260984 700068
rect 260840 699984 260892 699990
rect 260840 699926 260892 699932
rect 259184 699916 259236 699922
rect 259184 699858 259236 699864
rect 257896 699848 257948 699854
rect 257896 699790 257948 699796
rect 257908 402974 257936 699790
rect 257908 402946 258028 402974
rect 257896 391400 257948 391406
rect 257896 391342 257948 391348
rect 257804 390312 257856 390318
rect 257804 390254 257856 390260
rect 257908 387954 257936 391342
rect 255576 387926 255912 387954
rect 256036 387926 256280 387954
rect 256404 387926 256556 387954
rect 256864 387926 257108 387954
rect 257232 387926 257568 387954
rect 257692 387926 257936 387954
rect 258000 387954 258028 402946
rect 259196 393314 259224 699858
rect 259644 699780 259696 699786
rect 259644 699722 259696 699728
rect 259276 434716 259328 434722
rect 259276 434658 259328 434664
rect 258736 393286 259224 393314
rect 258736 387954 258764 393286
rect 259184 391468 259236 391474
rect 259184 391410 259236 391416
rect 259196 387954 259224 391410
rect 258000 387926 258060 387954
rect 258520 387926 258764 387954
rect 258888 387926 259224 387954
rect 259288 387954 259316 434658
rect 259656 402974 259684 699722
rect 259656 402946 260328 402974
rect 259828 391604 259880 391610
rect 259828 391546 259880 391552
rect 259644 391536 259696 391542
rect 259644 391478 259696 391484
rect 259656 387954 259684 391478
rect 259840 387954 259868 391546
rect 260300 387954 260328 402946
rect 260852 391678 260880 699926
rect 260840 391672 260892 391678
rect 260840 391614 260892 391620
rect 260944 390590 260972 700062
rect 261024 699712 261076 699718
rect 261024 699654 261076 699660
rect 261484 699712 261536 699718
rect 261484 699654 261536 699660
rect 260932 390584 260984 390590
rect 260932 390526 260984 390532
rect 261036 388634 261064 699654
rect 261496 434722 261524 699654
rect 261484 434716 261536 434722
rect 261484 434658 261536 434664
rect 261116 391672 261168 391678
rect 261116 391614 261168 391620
rect 260944 388606 261064 388634
rect 260944 387954 260972 388606
rect 261128 387954 261156 391614
rect 262232 390590 262260 700946
rect 262312 700868 262364 700874
rect 262312 700810 262364 700816
rect 262324 390658 262352 700810
rect 262496 700800 262548 700806
rect 262496 700742 262548 700748
rect 262404 700052 262456 700058
rect 262404 699994 262456 700000
rect 262312 390652 262364 390658
rect 262312 390594 262364 390600
rect 261576 390584 261628 390590
rect 261576 390526 261628 390532
rect 262220 390584 262272 390590
rect 262220 390526 262272 390532
rect 261588 387954 261616 390526
rect 262416 387954 262444 699994
rect 262508 402974 262536 700742
rect 263692 700596 263744 700602
rect 263692 700538 263744 700544
rect 263600 700528 263652 700534
rect 263600 700470 263652 700476
rect 262508 402946 262812 402974
rect 262496 390584 262548 390590
rect 262496 390526 262548 390532
rect 259288 387926 259348 387954
rect 259656 387926 259716 387954
rect 259840 387926 260176 387954
rect 260300 387926 260636 387954
rect 260944 387926 261004 387954
rect 261128 387926 261464 387954
rect 261588 387926 261832 387954
rect 262292 387926 262444 387954
rect 262508 387954 262536 390526
rect 262784 387954 262812 402946
rect 263232 390652 263284 390658
rect 263232 390594 263284 390600
rect 263244 387954 263272 390594
rect 263612 390590 263640 700470
rect 263600 390584 263652 390590
rect 263600 390526 263652 390532
rect 263704 387954 263732 700538
rect 263784 700460 263836 700466
rect 263784 700402 263836 700408
rect 263796 402974 263824 700402
rect 267660 699718 267688 703520
rect 283656 700528 283708 700534
rect 283656 700470 283708 700476
rect 269764 700460 269816 700466
rect 269764 700402 269816 700408
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 264980 683256 265032 683262
rect 264980 683198 265032 683204
rect 263796 402946 264100 402974
rect 264072 387954 264100 402946
rect 264428 390584 264480 390590
rect 264428 390526 264480 390532
rect 264440 387954 264468 390526
rect 264992 387954 265020 683198
rect 265072 670812 265124 670818
rect 265072 670754 265124 670760
rect 265084 390590 265112 670754
rect 265164 656940 265216 656946
rect 265164 656882 265216 656888
rect 265176 402974 265204 656882
rect 266360 632120 266412 632126
rect 266360 632062 266412 632068
rect 265176 402946 265296 402974
rect 265072 390584 265124 390590
rect 265072 390526 265124 390532
rect 265268 387954 265296 402946
rect 265716 390584 265768 390590
rect 265716 390526 265768 390532
rect 265728 387954 265756 390526
rect 266372 387954 266400 632062
rect 266452 618316 266504 618322
rect 266452 618258 266504 618264
rect 266464 390590 266492 618258
rect 266544 605872 266596 605878
rect 266544 605814 266596 605820
rect 266452 390584 266504 390590
rect 266452 390526 266504 390532
rect 266556 387954 266584 605814
rect 266636 579692 266688 579698
rect 266636 579634 266688 579640
rect 266648 402974 266676 579634
rect 267740 565888 267792 565894
rect 267740 565830 267792 565836
rect 266648 402946 267412 402974
rect 266912 390584 266964 390590
rect 266912 390526 266964 390532
rect 266924 387954 266952 390526
rect 267384 387954 267412 402946
rect 267752 390590 267780 565830
rect 267832 553444 267884 553450
rect 267832 553386 267884 553392
rect 267740 390584 267792 390590
rect 267740 390526 267792 390532
rect 267844 387954 267872 553386
rect 267924 527196 267976 527202
rect 267924 527138 267976 527144
rect 267936 402974 267964 527138
rect 269120 514820 269172 514826
rect 269120 514762 269172 514768
rect 267936 402946 268700 402974
rect 268200 390584 268252 390590
rect 268200 390526 268252 390532
rect 268212 387954 268240 390526
rect 268672 387954 268700 402946
rect 269132 390590 269160 514762
rect 269212 501016 269264 501022
rect 269212 500958 269264 500964
rect 269120 390584 269172 390590
rect 269120 390526 269172 390532
rect 269224 387954 269252 500958
rect 269304 474768 269356 474774
rect 269304 474710 269356 474716
rect 269316 402974 269344 474710
rect 269316 402946 269712 402974
rect 269488 390584 269540 390590
rect 269488 390526 269540 390532
rect 269500 387954 269528 390526
rect 269684 388090 269712 402946
rect 269776 391542 269804 700402
rect 283564 699712 283616 699718
rect 283564 699654 283616 699660
rect 270776 462392 270828 462398
rect 270776 462334 270828 462340
rect 270592 448588 270644 448594
rect 270592 448530 270644 448536
rect 270500 397520 270552 397526
rect 270500 397462 270552 397468
rect 269764 391536 269816 391542
rect 269764 391478 269816 391484
rect 270512 389978 270540 397462
rect 270500 389972 270552 389978
rect 270500 389914 270552 389920
rect 270222 389872 270278 389881
rect 270222 389807 270224 389816
rect 270276 389807 270278 389816
rect 270224 389778 270276 389784
rect 270604 388226 270632 448530
rect 270684 422340 270736 422346
rect 270684 422282 270736 422288
rect 270696 390590 270724 422282
rect 270684 390584 270736 390590
rect 270684 390526 270736 390532
rect 270558 388198 270632 388226
rect 269684 388062 269896 388090
rect 269868 387954 269896 388062
rect 262508 387926 262660 387954
rect 262784 387926 263120 387954
rect 263244 387926 263488 387954
rect 263704 387926 263948 387954
rect 264072 387926 264316 387954
rect 264440 387926 264776 387954
rect 264992 387926 265144 387954
rect 265268 387926 265604 387954
rect 265728 387926 265972 387954
rect 266372 387926 266432 387954
rect 266556 387926 266800 387954
rect 266924 387926 267260 387954
rect 267384 387926 267628 387954
rect 267844 387926 268088 387954
rect 268212 387926 268548 387954
rect 268672 387926 268916 387954
rect 269224 387926 269376 387954
rect 269500 387926 269744 387954
rect 269868 387926 270204 387954
rect 270558 387940 270586 388198
rect 270788 387954 270816 462334
rect 271880 409896 271932 409902
rect 271880 409838 271932 409844
rect 271892 402974 271920 409838
rect 271892 402946 272012 402974
rect 271144 390584 271196 390590
rect 271144 390526 271196 390532
rect 271156 387954 271184 390526
rect 271512 389972 271564 389978
rect 271512 389914 271564 389920
rect 271604 389972 271656 389978
rect 271604 389914 271656 389920
rect 271524 387954 271552 389914
rect 271616 389881 271644 389914
rect 271602 389872 271658 389881
rect 271602 389807 271658 389816
rect 271984 387954 272012 402946
rect 283576 391406 283604 699654
rect 283668 391474 283696 700470
rect 283852 700466 283880 703520
rect 300136 700534 300164 703520
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 283840 700460 283892 700466
rect 283840 700402 283892 700408
rect 283932 700460 283984 700466
rect 283932 700402 283984 700408
rect 283944 699718 283972 700402
rect 332520 699854 332548 703520
rect 348804 699922 348832 703520
rect 364996 700466 365024 703520
rect 364984 700460 365036 700466
rect 364984 700402 365036 700408
rect 397472 700194 397500 703520
rect 413664 700262 413692 703520
rect 429856 700942 429884 703520
rect 429844 700936 429896 700942
rect 429844 700878 429896 700884
rect 462332 700738 462360 703520
rect 462320 700732 462372 700738
rect 462320 700674 462372 700680
rect 478524 700670 478552 703520
rect 478512 700664 478564 700670
rect 478512 700606 478564 700612
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 348792 699916 348844 699922
rect 348792 699858 348844 699864
rect 332508 699848 332560 699854
rect 332508 699790 332560 699796
rect 283932 699712 283984 699718
rect 283932 699654 283984 699660
rect 283656 391468 283708 391474
rect 283656 391410 283708 391416
rect 283564 391400 283616 391406
rect 283564 391342 283616 391348
rect 494072 391338 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700398 527220 703520
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 494060 391332 494112 391338
rect 494060 391274 494112 391280
rect 558932 391270 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 558920 391264 558972 391270
rect 558920 391206 558972 391212
rect 289084 390516 289136 390522
rect 289084 390458 289136 390464
rect 288992 390448 289044 390454
rect 288992 390390 289044 390396
rect 286968 390312 287020 390318
rect 286968 390254 287020 390260
rect 286784 390244 286836 390250
rect 286784 390186 286836 390192
rect 286600 390108 286652 390114
rect 286600 390050 286652 390056
rect 276940 389972 276992 389978
rect 276940 389914 276992 389920
rect 273260 389904 273312 389910
rect 273260 389846 273312 389852
rect 272800 389156 272852 389162
rect 272800 389098 272852 389104
rect 272340 389088 272392 389094
rect 272340 389030 272392 389036
rect 272352 387954 272380 389030
rect 272812 387954 272840 389098
rect 273272 387954 273300 389846
rect 275652 389836 275704 389842
rect 275652 389778 275704 389784
rect 274640 389224 274692 389230
rect 274640 389166 274692 389172
rect 273628 389020 273680 389026
rect 273628 388962 273680 388968
rect 273640 387954 273668 388962
rect 273996 388748 274048 388754
rect 273996 388690 274048 388696
rect 274008 387954 274036 388690
rect 274652 387954 274680 389166
rect 275284 388680 275336 388686
rect 275284 388622 275336 388628
rect 274824 388612 274876 388618
rect 274824 388554 274876 388560
rect 274836 387954 274864 388554
rect 275296 387954 275324 388622
rect 275664 387954 275692 389778
rect 276480 389768 276532 389774
rect 276480 389710 276532 389716
rect 276112 388544 276164 388550
rect 276112 388486 276164 388492
rect 276124 387954 276152 388486
rect 276492 387954 276520 389710
rect 276952 387954 276980 389914
rect 278228 389700 278280 389706
rect 278228 389642 278280 389648
rect 277768 389632 277820 389638
rect 277768 389574 277820 389580
rect 277492 388476 277544 388482
rect 277492 388418 277544 388424
rect 277504 387954 277532 388418
rect 277780 387954 277808 389574
rect 278240 387954 278268 389642
rect 284208 389632 284260 389638
rect 284208 389574 284260 389580
rect 279424 389564 279476 389570
rect 279424 389506 279476 389512
rect 284116 389564 284168 389570
rect 284116 389506 284168 389512
rect 279056 389496 279108 389502
rect 279056 389438 279108 389444
rect 278780 388408 278832 388414
rect 278780 388350 278832 388356
rect 278792 387954 278820 388350
rect 279068 387954 279096 389438
rect 279436 387954 279464 389506
rect 283748 389496 283800 389502
rect 281906 389464 281962 389473
rect 280712 389428 280764 389434
rect 283748 389438 283800 389444
rect 281906 389399 281962 389408
rect 280712 389370 280764 389376
rect 280252 389360 280304 389366
rect 280252 389302 280304 389308
rect 279884 388340 279936 388346
rect 279884 388282 279936 388288
rect 279896 387954 279924 388282
rect 280264 387954 280292 389302
rect 280724 387954 280752 389370
rect 281538 389328 281594 389337
rect 281538 389263 281594 389272
rect 281078 387968 281134 387977
rect 270788 387926 271032 387954
rect 271156 387926 271400 387954
rect 271524 387926 271860 387954
rect 271984 387926 272228 387954
rect 272352 387926 272688 387954
rect 272812 387926 273056 387954
rect 273272 387926 273516 387954
rect 273640 387926 273884 387954
rect 274008 387926 274344 387954
rect 274652 387926 274712 387954
rect 274836 387926 275172 387954
rect 275296 387926 275540 387954
rect 275664 387926 276000 387954
rect 276124 387926 276368 387954
rect 276492 387926 276828 387954
rect 276952 387926 277288 387954
rect 277504 387926 277656 387954
rect 277780 387926 278116 387954
rect 278240 387926 278484 387954
rect 278792 387926 278944 387954
rect 279068 387926 279312 387954
rect 279436 387926 279772 387954
rect 279896 387926 280140 387954
rect 280264 387926 280600 387954
rect 280724 387926 280968 387954
rect 281552 387954 281580 389263
rect 281920 387954 281948 389399
rect 283288 389360 283340 389366
rect 283288 389302 283340 389308
rect 282828 389224 282880 389230
rect 282828 389166 282880 389172
rect 282840 387954 282868 389166
rect 283300 387954 283328 389302
rect 283760 387954 283788 389438
rect 284128 387954 284156 389506
rect 281134 387926 281428 387954
rect 281552 387926 281796 387954
rect 281920 387926 282256 387954
rect 282624 387926 282868 387954
rect 283084 387926 283328 387954
rect 283452 387926 283788 387954
rect 283912 387926 284156 387954
rect 284220 387954 284248 389574
rect 285036 389428 285088 389434
rect 285036 389370 285088 389376
rect 285048 387954 285076 389370
rect 286416 388952 286468 388958
rect 286416 388894 286468 388900
rect 285126 388376 285182 388385
rect 285126 388311 285182 388320
rect 284220 387926 284280 387954
rect 284740 387926 285076 387954
rect 281078 387903 281134 387912
rect 240876 387874 240928 387880
rect 238096 387806 238444 387812
rect 238096 387790 238432 387806
rect 238556 387790 238708 387818
rect 234908 386510 234936 387790
rect 234896 386504 234948 386510
rect 234896 386446 234948 386452
rect 233054 385248 233110 385257
rect 233054 385183 233110 385192
rect 232962 379672 233018 379681
rect 232962 379607 233018 379616
rect 232870 374096 232926 374105
rect 232870 374031 232926 374040
rect 232778 368520 232834 368529
rect 232778 368455 232834 368464
rect 232686 357368 232742 357377
rect 232686 357303 232742 357312
rect 232594 346216 232650 346225
rect 232594 346151 232650 346160
rect 232502 340776 232558 340785
rect 232502 340711 232558 340720
rect 86868 336728 86920 336734
rect 68926 336696 68982 336705
rect 86868 336670 86920 336676
rect 68926 336631 68982 336640
rect 62026 336560 62082 336569
rect 44088 336524 44140 336530
rect 62026 336495 62082 336504
rect 44088 336466 44140 336472
rect 42708 336388 42760 336394
rect 42708 336330 42760 336336
rect 28908 336320 28960 336326
rect 28908 336262 28960 336268
rect 37186 336288 37242 336297
rect 20628 336252 20680 336258
rect 20628 336194 20680 336200
rect 7564 336116 7616 336122
rect 7564 336058 7616 336064
rect 6644 306264 6696 306270
rect 6644 306206 6696 306212
rect 6552 202836 6604 202842
rect 6552 202778 6604 202784
rect 6460 150408 6512 150414
rect 6460 150350 6512 150356
rect 6368 97912 6420 97918
rect 6368 97854 6420 97860
rect 6276 59220 6328 59226
rect 6276 59162 6328 59168
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 5276 6886 5488 6914
rect 4804 6520 4856 6526
rect 4804 6462 4856 6468
rect 5276 480 5304 6886
rect 7576 3330 7604 336058
rect 19338 335608 19394 335617
rect 19338 335543 19394 335552
rect 11058 335472 11114 335481
rect 10968 335436 11020 335442
rect 11058 335407 11114 335416
rect 10968 335378 11020 335384
rect 9588 177404 9640 177410
rect 9588 177346 9640 177352
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 6460 3324 6512 3330
rect 6460 3266 6512 3272
rect 7564 3324 7616 3330
rect 7564 3266 7616 3272
rect 6472 480 6500 3266
rect 7668 480 7696 4762
rect 9600 3534 9628 177346
rect 10980 3534 11008 335378
rect 11072 16574 11100 335407
rect 16578 334656 16634 334665
rect 16578 334591 16634 334600
rect 16592 16574 16620 334591
rect 19248 331900 19300 331906
rect 19248 331842 19300 331848
rect 11072 16546 11192 16574
rect 16592 16546 17080 16574
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 11164 480 11192 16546
rect 13544 7608 13596 7614
rect 13544 7550 13596 7556
rect 12348 4888 12400 4894
rect 12348 4830 12400 4836
rect 12360 480 12388 4830
rect 13556 480 13584 7550
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14752 480 14780 3402
rect 15934 3360 15990 3369
rect 15934 3295 15990 3304
rect 15948 480 15976 3295
rect 17052 480 17080 16546
rect 19260 3534 19288 331842
rect 19352 16574 19380 335543
rect 19352 16546 20208 16574
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 18248 480 18276 3470
rect 19444 480 19472 3470
rect 20180 490 20208 16546
rect 20640 3534 20668 336194
rect 28814 336016 28870 336025
rect 28814 335951 28870 335960
rect 26238 334792 26294 334801
rect 26238 334727 26294 334736
rect 23388 330540 23440 330546
rect 23388 330482 23440 330488
rect 21824 7676 21876 7682
rect 21824 7618 21876 7624
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20456 598 20668 626
rect 20456 490 20484 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20180 462 20484 490
rect 20640 480 20668 598
rect 21836 480 21864 7618
rect 23400 6914 23428 330482
rect 26252 16574 26280 334727
rect 28828 16574 28856 335951
rect 26252 16546 26556 16574
rect 23032 6886 23428 6914
rect 23032 480 23060 6886
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 25318 3496 25374 3505
rect 24228 480 24256 3470
rect 25318 3431 25374 3440
rect 25332 480 25360 3431
rect 26528 480 26556 16546
rect 28736 16546 28856 16574
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 27724 480 27752 3538
rect 28736 3482 28764 16546
rect 28920 6914 28948 336262
rect 37186 336223 37242 336232
rect 35806 336152 35862 336161
rect 35806 336087 35862 336096
rect 33140 333328 33192 333334
rect 33140 333270 33192 333276
rect 29000 333260 29052 333266
rect 29000 333202 29052 333208
rect 29012 16574 29040 333202
rect 33152 16574 33180 333270
rect 29012 16546 30144 16574
rect 33152 16546 33640 16574
rect 28828 6886 28948 6914
rect 28828 3602 28856 6886
rect 28816 3596 28868 3602
rect 28816 3538 28868 3544
rect 28736 3454 28948 3482
rect 28920 480 28948 3454
rect 30116 480 30144 16546
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 31300 3596 31352 3602
rect 31300 3538 31352 3544
rect 31312 480 31340 3538
rect 32416 480 32444 3606
rect 33612 480 33640 16546
rect 35820 3398 35848 336087
rect 35900 333396 35952 333402
rect 35900 333338 35952 333344
rect 35912 16574 35940 333338
rect 35912 16546 36768 16574
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 34808 480 34836 3334
rect 36004 480 36032 3334
rect 36740 490 36768 16546
rect 37200 3398 37228 336223
rect 40040 331288 40092 331294
rect 40040 331230 40092 331236
rect 40052 16574 40080 331230
rect 40052 16546 40264 16574
rect 39580 3800 39632 3806
rect 39580 3742 39632 3748
rect 38384 3732 38436 3738
rect 38384 3674 38436 3680
rect 37188 3392 37240 3398
rect 37188 3334 37240 3340
rect 37016 598 37228 626
rect 37016 490 37044 598
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 36740 462 37044 490
rect 37200 480 37228 598
rect 38396 480 38424 3674
rect 39592 480 39620 3742
rect 40236 490 40264 16546
rect 42720 3398 42748 336330
rect 44100 3398 44128 336466
rect 53746 336424 53802 336433
rect 53746 336359 53802 336368
rect 52366 333704 52422 333713
rect 52366 333639 52422 333648
rect 48226 333568 48282 333577
rect 48226 333503 48282 333512
rect 48240 6914 48268 333503
rect 49608 86284 49660 86290
rect 49608 86226 49660 86232
rect 47872 6886 48268 6914
rect 44272 6180 44324 6186
rect 44272 6122 44324 6128
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 42708 3392 42760 3398
rect 42708 3334 42760 3340
rect 43076 3392 43128 3398
rect 43076 3334 43128 3340
rect 44088 3392 44140 3398
rect 44088 3334 44140 3340
rect 40512 598 40724 626
rect 40512 490 40540 598
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 462 40540 490
rect 40696 480 40724 598
rect 41892 480 41920 3334
rect 43088 480 43116 3334
rect 44284 480 44312 6122
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 45468 3868 45520 3874
rect 45468 3810 45520 3816
rect 45480 480 45508 3810
rect 46676 480 46704 3878
rect 47872 480 47900 6886
rect 49620 3398 49648 86226
rect 50160 4004 50212 4010
rect 50160 3946 50212 3952
rect 48964 3392 49016 3398
rect 48964 3334 49016 3340
rect 49608 3392 49660 3398
rect 49608 3334 49660 3340
rect 48976 480 49004 3334
rect 50172 480 50200 3946
rect 52380 3398 52408 333639
rect 53656 177472 53708 177478
rect 53656 177414 53708 177420
rect 53668 3398 53696 177414
rect 51356 3392 51408 3398
rect 51356 3334 51408 3340
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 52552 3392 52604 3398
rect 52552 3334 52604 3340
rect 53656 3392 53708 3398
rect 53656 3334 53708 3340
rect 51368 480 51396 3334
rect 52564 480 52592 3334
rect 53760 480 53788 336359
rect 55126 333840 55182 333849
rect 55126 333775 55182 333784
rect 55140 6914 55168 333775
rect 61936 333464 61988 333470
rect 61936 333406 61988 333412
rect 59268 331968 59320 331974
rect 59268 331910 59320 331916
rect 54956 6886 55168 6914
rect 54956 480 54984 6886
rect 56046 6216 56102 6225
rect 56046 6151 56102 6160
rect 56060 480 56088 6151
rect 57244 4140 57296 4146
rect 57244 4082 57296 4088
rect 57256 480 57284 4082
rect 59280 3398 59308 331910
rect 61948 16574 61976 333406
rect 61856 16546 61976 16574
rect 59636 7744 59688 7750
rect 59636 7686 59688 7692
rect 58440 3392 58492 3398
rect 58440 3334 58492 3340
rect 59268 3392 59320 3398
rect 59268 3334 59320 3340
rect 58452 480 58480 3334
rect 59648 480 59676 7686
rect 60832 4072 60884 4078
rect 60832 4014 60884 4020
rect 60844 480 60872 4014
rect 61856 3482 61884 16546
rect 62040 6914 62068 336495
rect 66168 333532 66220 333538
rect 66168 333474 66220 333480
rect 64788 177540 64840 177546
rect 64788 177482 64840 177488
rect 63224 7812 63276 7818
rect 63224 7754 63276 7760
rect 61948 6886 62068 6914
rect 61948 4078 61976 6886
rect 61936 4072 61988 4078
rect 61936 4014 61988 4020
rect 61856 3454 62068 3482
rect 62040 480 62068 3454
rect 63236 480 63264 7754
rect 64800 3398 64828 177482
rect 66180 3398 66208 333474
rect 66720 7880 66772 7886
rect 66720 7822 66772 7828
rect 64328 3392 64380 3398
rect 64328 3334 64380 3340
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 65524 3392 65576 3398
rect 65524 3334 65576 3340
rect 66168 3392 66220 3398
rect 66168 3334 66220 3340
rect 64340 480 64368 3334
rect 65536 480 65564 3334
rect 66732 480 66760 7822
rect 68940 3398 68968 336631
rect 82728 336592 82780 336598
rect 82728 336534 82780 336540
rect 75828 336456 75880 336462
rect 75828 336398 75880 336404
rect 70308 333600 70360 333606
rect 70308 333542 70360 333548
rect 70216 7948 70268 7954
rect 70216 7890 70268 7896
rect 69112 4140 69164 4146
rect 69112 4082 69164 4088
rect 67916 3392 67968 3398
rect 67916 3334 67968 3340
rect 68928 3392 68980 3398
rect 68928 3334 68980 3340
rect 67928 480 67956 3334
rect 69124 480 69152 4082
rect 70228 3482 70256 7890
rect 70320 4146 70348 333542
rect 73068 80708 73120 80714
rect 73068 80650 73120 80656
rect 70308 4140 70360 4146
rect 70308 4082 70360 4088
rect 71504 4140 71556 4146
rect 71504 4082 71556 4088
rect 70228 3454 70348 3482
rect 70320 480 70348 3454
rect 71516 480 71544 4082
rect 73080 3398 73108 80650
rect 73804 8016 73856 8022
rect 73804 7958 73856 7964
rect 72608 3392 72660 3398
rect 72608 3334 72660 3340
rect 73068 3392 73120 3398
rect 73068 3334 73120 3340
rect 72620 480 72648 3334
rect 73816 480 73844 7958
rect 75840 3398 75868 336398
rect 81348 332036 81400 332042
rect 81348 331978 81400 331984
rect 79968 84924 80020 84930
rect 79968 84866 80020 84872
rect 77208 84856 77260 84862
rect 77208 84798 77260 84804
rect 77220 3398 77248 84798
rect 77392 8084 77444 8090
rect 77392 8026 77444 8032
rect 75000 3392 75052 3398
rect 75000 3334 75052 3340
rect 75828 3392 75880 3398
rect 75828 3334 75880 3340
rect 76196 3392 76248 3398
rect 76196 3334 76248 3340
rect 77208 3392 77260 3398
rect 77208 3334 77260 3340
rect 75012 480 75040 3334
rect 76208 480 76236 3334
rect 77404 480 77432 8026
rect 79980 6914 80008 84866
rect 79704 6886 80008 6914
rect 78588 3324 78640 3330
rect 78588 3266 78640 3272
rect 78600 480 78628 3266
rect 79704 480 79732 6886
rect 81360 3398 81388 331978
rect 82740 3398 82768 336534
rect 85488 332104 85540 332110
rect 85488 332046 85540 332052
rect 84108 87644 84160 87650
rect 84108 87586 84160 87592
rect 84120 3398 84148 87586
rect 85500 3398 85528 332046
rect 86880 6914 86908 336670
rect 100668 336660 100720 336666
rect 100668 336602 100720 336608
rect 93768 335980 93820 335986
rect 93768 335922 93820 335928
rect 92386 334928 92442 334937
rect 92386 334863 92442 334872
rect 88248 333668 88300 333674
rect 88248 333610 88300 333616
rect 88260 6914 88288 333610
rect 86696 6886 86908 6914
rect 87984 6886 88288 6914
rect 86696 3398 86724 6886
rect 86866 6352 86922 6361
rect 86866 6287 86922 6296
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 81348 3392 81400 3398
rect 81348 3334 81400 3340
rect 82084 3392 82136 3398
rect 82084 3334 82136 3340
rect 82728 3392 82780 3398
rect 82728 3334 82780 3340
rect 83280 3392 83332 3398
rect 83280 3334 83332 3340
rect 84108 3392 84160 3398
rect 84108 3334 84160 3340
rect 84476 3392 84528 3398
rect 84476 3334 84528 3340
rect 85488 3392 85540 3398
rect 85488 3334 85540 3340
rect 85672 3392 85724 3398
rect 85672 3334 85724 3340
rect 86684 3392 86736 3398
rect 86684 3334 86736 3340
rect 80900 480 80928 3334
rect 82096 480 82124 3334
rect 83292 480 83320 3334
rect 84488 480 84516 3334
rect 85684 480 85712 3334
rect 86880 480 86908 6287
rect 87984 480 88012 6886
rect 90362 6488 90418 6497
rect 90362 6423 90418 6432
rect 89168 3256 89220 3262
rect 89168 3198 89220 3204
rect 89180 480 89208 3198
rect 90376 480 90404 6423
rect 92400 3398 92428 334863
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 92388 3392 92440 3398
rect 92388 3334 92440 3340
rect 91572 480 91600 3334
rect 93780 3330 93808 335922
rect 95148 333736 95200 333742
rect 95148 333678 95200 333684
rect 93950 6624 94006 6633
rect 93950 6559 94006 6568
rect 92756 3324 92808 3330
rect 92756 3266 92808 3272
rect 93768 3324 93820 3330
rect 93768 3266 93820 3272
rect 92768 480 92796 3266
rect 93964 480 93992 6559
rect 95160 480 95188 333678
rect 97908 332172 97960 332178
rect 97908 332114 97960 332120
rect 97920 3330 97948 332114
rect 98644 8220 98696 8226
rect 98644 8162 98696 8168
rect 97448 3324 97500 3330
rect 97448 3266 97500 3272
rect 97908 3324 97960 3330
rect 97908 3266 97960 3272
rect 96252 3188 96304 3194
rect 96252 3130 96304 3136
rect 96264 480 96292 3130
rect 97460 480 97488 3266
rect 98656 480 98684 8162
rect 100680 3330 100708 336602
rect 107568 335912 107620 335918
rect 107568 335854 107620 335860
rect 104808 177608 104860 177614
rect 104808 177550 104860 177556
rect 102048 86352 102100 86358
rect 102048 86294 102100 86300
rect 102060 3330 102088 86294
rect 102232 8152 102284 8158
rect 102232 8094 102284 8100
rect 99840 3324 99892 3330
rect 99840 3266 99892 3272
rect 100668 3324 100720 3330
rect 100668 3266 100720 3272
rect 101036 3324 101088 3330
rect 101036 3266 101088 3272
rect 102048 3324 102100 3330
rect 102048 3266 102100 3272
rect 99852 480 99880 3266
rect 101048 480 101076 3266
rect 102244 480 102272 8094
rect 104820 6914 104848 177550
rect 105728 7540 105780 7546
rect 105728 7482 105780 7488
rect 104544 6886 104848 6914
rect 103336 3188 103388 3194
rect 103336 3130 103388 3136
rect 103348 480 103376 3130
rect 104544 480 104572 6886
rect 105740 480 105768 7482
rect 107580 3126 107608 335854
rect 114468 335844 114520 335850
rect 114468 335786 114520 335792
rect 108948 177676 109000 177682
rect 108948 177618 109000 177624
rect 108960 3126 108988 177618
rect 111708 84992 111760 84998
rect 111708 84934 111760 84940
rect 109316 8288 109368 8294
rect 109316 8230 109368 8236
rect 106924 3120 106976 3126
rect 106924 3062 106976 3068
rect 107568 3120 107620 3126
rect 107568 3062 107620 3068
rect 108120 3120 108172 3126
rect 108120 3062 108172 3068
rect 108948 3120 109000 3126
rect 108948 3062 109000 3068
rect 106936 480 106964 3062
rect 108132 480 108160 3062
rect 109328 480 109356 8230
rect 111720 6914 111748 84934
rect 112812 7404 112864 7410
rect 112812 7346 112864 7352
rect 111628 6886 111748 6914
rect 110512 3120 110564 3126
rect 110512 3062 110564 3068
rect 110524 480 110552 3062
rect 111628 480 111656 6886
rect 112824 480 112852 7346
rect 114480 3058 114508 335786
rect 125508 335776 125560 335782
rect 125508 335718 125560 335724
rect 124128 335708 124180 335714
rect 124128 335650 124180 335656
rect 115848 87712 115900 87718
rect 115848 87654 115900 87660
rect 115860 3058 115888 87654
rect 116400 7472 116452 7478
rect 116400 7414 116452 7420
rect 114008 3052 114060 3058
rect 114008 2994 114060 3000
rect 114468 3052 114520 3058
rect 114468 2994 114520 3000
rect 115204 3052 115256 3058
rect 115204 2994 115256 3000
rect 115848 3052 115900 3058
rect 115848 2994 115900 3000
rect 114020 480 114048 2994
rect 115216 480 115244 2994
rect 116412 480 116440 7414
rect 119896 7336 119948 7342
rect 119896 7278 119948 7284
rect 118792 6248 118844 6254
rect 118792 6190 118844 6196
rect 117596 2916 117648 2922
rect 117596 2858 117648 2864
rect 117608 480 117636 2858
rect 118804 480 118832 6190
rect 119908 480 119936 7278
rect 122288 6316 122340 6322
rect 122288 6258 122340 6264
rect 121092 2984 121144 2990
rect 121092 2926 121144 2932
rect 121104 480 121132 2926
rect 122300 480 122328 6258
rect 124140 3058 124168 335650
rect 125520 3058 125548 335718
rect 136546 335336 136602 335345
rect 136546 335271 136602 335280
rect 219348 335300 219400 335306
rect 133786 335200 133842 335209
rect 133786 335135 133842 335144
rect 129646 335064 129702 335073
rect 129646 334999 129702 335008
rect 128268 333804 128320 333810
rect 128268 333746 128320 333752
rect 126888 332240 126940 332246
rect 126888 332182 126940 332188
rect 126900 3058 126928 332182
rect 128174 4992 128230 5001
rect 128174 4927 128230 4936
rect 123484 3052 123536 3058
rect 123484 2994 123536 3000
rect 124128 3052 124180 3058
rect 124128 2994 124180 3000
rect 124680 3052 124732 3058
rect 124680 2994 124732 3000
rect 125508 3052 125560 3058
rect 125508 2994 125560 3000
rect 125876 3052 125928 3058
rect 125876 2994 125928 3000
rect 126888 3052 126940 3058
rect 126888 2994 126940 3000
rect 126980 3052 127032 3058
rect 126980 2994 127032 3000
rect 123496 480 123524 2994
rect 124692 480 124720 2994
rect 125888 480 125916 2994
rect 126992 480 127020 2994
rect 128188 480 128216 4927
rect 128280 3058 128308 333746
rect 129660 6914 129688 334999
rect 131028 80776 131080 80782
rect 131028 80718 131080 80724
rect 129384 6886 129688 6914
rect 128268 3052 128320 3058
rect 128268 2994 128320 3000
rect 129384 480 129412 6886
rect 131040 2922 131068 80718
rect 131762 5128 131818 5137
rect 131762 5063 131818 5072
rect 130568 2916 130620 2922
rect 130568 2858 130620 2864
rect 131028 2916 131080 2922
rect 131028 2858 131080 2864
rect 130580 480 130608 2858
rect 131776 480 131804 5063
rect 133800 2922 133828 335135
rect 135168 83496 135220 83502
rect 135168 83438 135220 83444
rect 135180 2922 135208 83438
rect 136560 6914 136588 335271
rect 219348 335242 219400 335248
rect 201408 335232 201460 335238
rect 201408 335174 201460 335180
rect 194416 335164 194468 335170
rect 194416 335106 194468 335112
rect 190368 335028 190420 335034
rect 190368 334970 190420 334976
rect 186136 334960 186188 334966
rect 186136 334902 186188 334908
rect 183468 334892 183520 334898
rect 183468 334834 183520 334840
rect 179328 334824 179380 334830
rect 179328 334766 179380 334772
rect 169576 334756 169628 334762
rect 169576 334698 169628 334704
rect 165528 334688 165580 334694
rect 165528 334630 165580 334636
rect 158628 334620 158680 334626
rect 158628 334562 158680 334568
rect 144826 334520 144882 334529
rect 144826 334455 144882 334464
rect 144736 333872 144788 333878
rect 144736 333814 144788 333820
rect 140688 332308 140740 332314
rect 140688 332250 140740 332256
rect 136468 6886 136588 6914
rect 135260 6384 135312 6390
rect 135260 6326 135312 6332
rect 132960 2916 133012 2922
rect 132960 2858 133012 2864
rect 133788 2916 133840 2922
rect 133788 2858 133840 2864
rect 134156 2916 134208 2922
rect 134156 2858 134208 2864
rect 135168 2916 135220 2922
rect 135168 2858 135220 2864
rect 132972 480 133000 2858
rect 134168 480 134196 2858
rect 135272 480 135300 6326
rect 136468 480 136496 6886
rect 138848 6452 138900 6458
rect 138848 6394 138900 6400
rect 137650 5264 137706 5273
rect 137650 5199 137706 5208
rect 137664 480 137692 5199
rect 138860 480 138888 6394
rect 140700 2922 140728 332250
rect 142436 6520 142488 6526
rect 142436 6462 142488 6468
rect 141240 4956 141292 4962
rect 141240 4898 141292 4904
rect 140044 2916 140096 2922
rect 140044 2858 140096 2864
rect 140688 2916 140740 2922
rect 140688 2858 140740 2864
rect 140056 480 140084 2858
rect 141252 480 141280 4898
rect 142448 480 142476 6462
rect 143540 2916 143592 2922
rect 143540 2858 143592 2864
rect 143552 480 143580 2858
rect 144748 480 144776 333814
rect 144840 2922 144868 334455
rect 147588 333940 147640 333946
rect 147588 333882 147640 333888
rect 145932 6588 145984 6594
rect 145932 6530 145984 6536
rect 144828 2916 144880 2922
rect 144828 2858 144880 2864
rect 145944 480 145972 6530
rect 147600 2922 147628 333882
rect 148968 333192 149020 333198
rect 148968 333134 149020 333140
rect 148980 2922 149008 333134
rect 153108 333124 153160 333130
rect 153108 333066 153160 333072
rect 151728 333056 151780 333062
rect 151728 332998 151780 333004
rect 149520 6656 149572 6662
rect 149520 6598 149572 6604
rect 147128 2916 147180 2922
rect 147128 2858 147180 2864
rect 147588 2916 147640 2922
rect 147588 2858 147640 2864
rect 148324 2916 148376 2922
rect 148324 2858 148376 2864
rect 148968 2916 149020 2922
rect 148968 2858 149020 2864
rect 147140 480 147168 2858
rect 148336 480 148364 2858
rect 149532 480 149560 6598
rect 151740 2922 151768 332998
rect 153016 6724 153068 6730
rect 153016 6666 153068 6672
rect 150624 2916 150676 2922
rect 150624 2858 150676 2864
rect 151728 2916 151780 2922
rect 151728 2858 151780 2864
rect 151820 2916 151872 2922
rect 151820 2858 151872 2864
rect 150636 480 150664 2858
rect 151832 480 151860 2858
rect 153028 480 153056 6666
rect 153120 2922 153148 333066
rect 154488 332988 154540 332994
rect 154488 332930 154540 332936
rect 154500 6914 154528 332930
rect 155868 80844 155920 80850
rect 155868 80786 155920 80792
rect 154224 6886 154528 6914
rect 153108 2916 153160 2922
rect 153108 2858 153160 2864
rect 154224 480 154252 6886
rect 155880 2922 155908 80786
rect 156604 6792 156656 6798
rect 156604 6734 156656 6740
rect 155408 2916 155460 2922
rect 155408 2858 155460 2864
rect 155868 2916 155920 2922
rect 155868 2858 155920 2864
rect 155420 480 155448 2858
rect 156616 480 156644 6734
rect 158640 2922 158668 334562
rect 161388 332376 161440 332382
rect 161388 332318 161440 332324
rect 160008 83564 160060 83570
rect 160008 83506 160060 83512
rect 160020 2922 160048 83506
rect 161400 6914 161428 332318
rect 162768 85060 162820 85066
rect 162768 85002 162820 85008
rect 162780 6914 162808 85002
rect 161308 6886 161428 6914
rect 162504 6886 162808 6914
rect 160100 6860 160152 6866
rect 160100 6802 160152 6808
rect 157800 2916 157852 2922
rect 157800 2858 157852 2864
rect 158628 2916 158680 2922
rect 158628 2858 158680 2864
rect 158904 2916 158956 2922
rect 158904 2858 158956 2864
rect 160008 2916 160060 2922
rect 160008 2858 160060 2864
rect 157812 480 157840 2858
rect 158916 480 158944 2858
rect 160112 480 160140 6802
rect 161308 480 161336 6886
rect 162504 480 162532 6886
rect 163688 5024 163740 5030
rect 163688 4966 163740 4972
rect 163700 480 163728 4966
rect 165540 2922 165568 334630
rect 167184 5160 167236 5166
rect 167184 5102 167236 5108
rect 166080 5092 166132 5098
rect 166080 5034 166132 5040
rect 164884 2916 164936 2922
rect 164884 2858 164936 2864
rect 165528 2916 165580 2922
rect 165528 2858 165580 2864
rect 164896 480 164924 2858
rect 166092 480 166120 5034
rect 167196 480 167224 5102
rect 169588 2922 169616 334698
rect 177856 332444 177908 332450
rect 177856 332386 177908 332392
rect 174268 5432 174320 5438
rect 174268 5374 174320 5380
rect 173164 5364 173216 5370
rect 173164 5306 173216 5312
rect 170772 5296 170824 5302
rect 170772 5238 170824 5244
rect 169668 5228 169720 5234
rect 169668 5170 169720 5176
rect 168380 2916 168432 2922
rect 168380 2858 168432 2864
rect 169576 2916 169628 2922
rect 169576 2858 169628 2864
rect 168392 480 168420 2858
rect 169680 2666 169708 5170
rect 169588 2638 169708 2666
rect 169588 480 169616 2638
rect 170784 480 170812 5238
rect 171968 2916 172020 2922
rect 171968 2858 172020 2864
rect 171980 480 172008 2858
rect 173176 480 173204 5306
rect 174280 480 174308 5374
rect 177868 2922 177896 332386
rect 179340 6914 179368 334766
rect 180708 332920 180760 332926
rect 180708 332862 180760 332868
rect 179064 6886 179368 6914
rect 177948 5500 178000 5506
rect 177948 5442 178000 5448
rect 176660 2916 176712 2922
rect 176660 2858 176712 2864
rect 177856 2916 177908 2922
rect 177856 2858 177908 2864
rect 175464 2848 175516 2854
rect 175464 2790 175516 2796
rect 175476 480 175504 2790
rect 176672 480 176700 2858
rect 177960 2802 177988 5442
rect 177868 2774 177988 2802
rect 177868 480 177896 2774
rect 179064 480 179092 6886
rect 180260 598 180472 626
rect 180260 480 180288 598
rect 180444 490 180472 598
rect 180720 490 180748 332862
rect 183480 6914 183508 334834
rect 184848 82136 184900 82142
rect 184848 82078 184900 82084
rect 184860 6914 184888 82078
rect 182560 6886 183508 6914
rect 184216 6886 184888 6914
rect 181444 4752 181496 4758
rect 181444 4694 181496 4700
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180444 462 180748 490
rect 181456 480 181484 4694
rect 182560 480 182588 6886
rect 183756 598 183968 626
rect 183756 480 183784 598
rect 183940 490 183968 598
rect 184216 490 184244 6886
rect 184940 4684 184992 4690
rect 184940 4626 184992 4632
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 183940 462 184244 490
rect 184952 480 184980 4626
rect 186148 480 186176 334902
rect 190380 6914 190408 334970
rect 194428 11762 194456 335106
rect 197268 335096 197320 335102
rect 197268 335038 197320 335044
rect 195888 86420 195940 86426
rect 195888 86362 195940 86368
rect 193220 11756 193272 11762
rect 193220 11698 193272 11704
rect 194416 11756 194468 11762
rect 194416 11698 194468 11704
rect 189736 6886 190408 6914
rect 188528 6112 188580 6118
rect 188528 6054 188580 6060
rect 187332 4616 187384 4622
rect 187332 4558 187384 4564
rect 187344 480 187372 4558
rect 188540 480 188568 6054
rect 189736 480 189764 6886
rect 192024 6044 192076 6050
rect 192024 5986 192076 5992
rect 190828 4548 190880 4554
rect 190828 4490 190880 4496
rect 190840 480 190868 4490
rect 192036 480 192064 5986
rect 193232 480 193260 11698
rect 195900 6914 195928 86362
rect 195624 6886 195928 6914
rect 194416 4480 194468 4486
rect 194416 4422 194468 4428
rect 194428 480 194456 4422
rect 195624 480 195652 6886
rect 196820 598 197032 626
rect 196820 480 196848 598
rect 197004 490 197032 598
rect 197280 490 197308 335038
rect 200028 87780 200080 87786
rect 200028 87722 200080 87728
rect 200040 6914 200068 87722
rect 201420 6914 201448 335174
rect 204168 334552 204220 334558
rect 204168 334494 204220 334500
rect 202696 89004 202748 89010
rect 202696 88946 202748 88952
rect 199120 6886 200068 6914
rect 200776 6886 201448 6914
rect 197912 4412 197964 4418
rect 197912 4354 197964 4360
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197004 462 197308 490
rect 197924 480 197952 4354
rect 199120 480 199148 6886
rect 200316 598 200528 626
rect 200316 480 200344 598
rect 200500 490 200528 598
rect 200776 490 200804 6886
rect 201500 4344 201552 4350
rect 201500 4286 201552 4292
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 200500 462 200804 490
rect 201512 480 201540 4286
rect 202708 480 202736 88946
rect 204180 6914 204208 334494
rect 211068 334484 211120 334490
rect 211068 334426 211120 334432
rect 208308 334416 208360 334422
rect 208308 334358 208360 334364
rect 208320 6914 208348 334358
rect 209688 332852 209740 332858
rect 209688 332794 209740 332800
rect 209700 6914 209728 332794
rect 210976 89072 211028 89078
rect 210976 89014 211028 89020
rect 210988 11762 211016 89014
rect 209780 11756 209832 11762
rect 209780 11698 209832 11704
rect 210976 11756 211028 11762
rect 210976 11698 211028 11704
rect 203904 6886 204208 6914
rect 207400 6886 208348 6914
rect 209056 6886 209728 6914
rect 203904 480 203932 6886
rect 206192 5976 206244 5982
rect 206192 5918 206244 5924
rect 205088 4276 205140 4282
rect 205088 4218 205140 4224
rect 205100 480 205128 4218
rect 206204 480 206232 5918
rect 207400 480 207428 6886
rect 208596 598 208808 626
rect 208596 480 208624 598
rect 208780 490 208808 598
rect 209056 490 209084 6886
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 208780 462 209084 490
rect 209792 480 209820 11698
rect 211080 6914 211108 334426
rect 215208 334280 215260 334286
rect 215208 334222 215260 334228
rect 212448 85128 212500 85134
rect 212448 85070 212500 85076
rect 212460 6914 212488 85070
rect 215220 6914 215248 334222
rect 219256 89140 219308 89146
rect 219256 89082 219308 89088
rect 216588 86488 216640 86494
rect 216588 86430 216640 86436
rect 216600 6914 216628 86430
rect 210988 6886 211108 6914
rect 212184 6886 212488 6914
rect 214944 6886 215248 6914
rect 215680 6886 216628 6914
rect 210988 480 211016 6886
rect 212184 480 212212 6886
rect 213368 5908 213420 5914
rect 213368 5850 213420 5856
rect 213380 480 213408 5850
rect 214484 598 214696 626
rect 214484 480 214512 598
rect 214668 490 214696 598
rect 214944 490 214972 6886
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 214668 462 214972 490
rect 215680 480 215708 6886
rect 216864 5840 216916 5846
rect 216864 5782 216916 5788
rect 216876 480 216904 5782
rect 218060 4208 218112 4214
rect 218060 4150 218112 4156
rect 218072 480 218100 4150
rect 219268 480 219296 89082
rect 219360 4214 219388 335242
rect 222108 334348 222160 334354
rect 222108 334290 222160 334296
rect 222120 6914 222148 334290
rect 229008 334212 229060 334218
rect 229008 334154 229060 334160
rect 226248 334144 226300 334150
rect 226248 334086 226300 334092
rect 226260 6914 226288 334086
rect 227628 332784 227680 332790
rect 227628 332726 227680 332732
rect 221568 6886 222148 6914
rect 225616 6886 226288 6914
rect 220452 5772 220504 5778
rect 220452 5714 220504 5720
rect 219348 4208 219400 4214
rect 219348 4150 219400 4156
rect 220464 480 220492 5714
rect 221568 480 221596 6886
rect 223948 5704 224000 5710
rect 223948 5646 224000 5652
rect 222752 4208 222804 4214
rect 222752 4150 222804 4156
rect 222764 480 222792 4150
rect 223960 480 223988 5646
rect 225156 598 225368 626
rect 225156 480 225184 598
rect 225340 490 225368 598
rect 225616 490 225644 6886
rect 227536 5636 227588 5642
rect 227536 5578 227588 5584
rect 226248 4208 226300 4214
rect 226246 4176 226248 4185
rect 226340 4208 226392 4214
rect 226300 4176 226302 4185
rect 226340 4150 226392 4156
rect 226246 4111 226302 4120
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 225340 462 225644 490
rect 226352 480 226380 4150
rect 227548 480 227576 5578
rect 227640 4214 227668 332726
rect 229020 6914 229048 334154
rect 230388 332716 230440 332722
rect 230388 332658 230440 332664
rect 230400 6914 230428 332658
rect 232516 236094 232544 340711
rect 232608 238134 232636 346151
rect 232596 238128 232648 238134
rect 232596 238070 232648 238076
rect 232700 238066 232728 357303
rect 232792 240786 232820 368455
rect 232780 240780 232832 240786
rect 232780 240722 232832 240728
rect 232688 238060 232740 238066
rect 232688 238002 232740 238008
rect 232884 237969 232912 374031
rect 232976 238513 233004 379607
rect 233068 238649 233096 385183
rect 234526 362944 234582 362953
rect 234526 362879 234582 362888
rect 234434 351792 234490 351801
rect 234434 351727 234490 351736
rect 234252 335640 234304 335646
rect 234252 335582 234304 335588
rect 234068 335572 234120 335578
rect 234068 335514 234120 335520
rect 233976 334076 234028 334082
rect 233976 334018 234028 334024
rect 233884 334008 233936 334014
rect 233884 333950 233936 333956
rect 233148 332648 233200 332654
rect 233148 332590 233200 332596
rect 233054 238640 233110 238649
rect 233054 238575 233110 238584
rect 232962 238504 233018 238513
rect 232962 238439 233018 238448
rect 232870 237960 232926 237969
rect 232870 237895 232926 237904
rect 232504 236088 232556 236094
rect 232504 236030 232556 236036
rect 228744 6886 229048 6914
rect 229848 6886 230428 6914
rect 227628 4208 227680 4214
rect 227720 4208 227772 4214
rect 227628 4150 227680 4156
rect 227718 4176 227720 4185
rect 227772 4176 227774 4185
rect 227718 4111 227774 4120
rect 228744 480 228772 6886
rect 229848 480 229876 6886
rect 231032 5568 231084 5574
rect 231032 5510 231084 5516
rect 231044 480 231072 5510
rect 232042 4040 232098 4049
rect 232042 3975 232098 3984
rect 232056 3602 232084 3975
rect 232044 3596 232096 3602
rect 232044 3538 232096 3544
rect 233160 3534 233188 332590
rect 233896 6914 233924 333950
rect 233804 6886 233924 6914
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233424 3528 233476 3534
rect 233424 3470 233476 3476
rect 232240 480 232268 3470
rect 233436 480 233464 3470
rect 233804 2854 233832 6886
rect 233988 2922 234016 334018
rect 234080 7342 234108 335514
rect 234160 335504 234212 335510
rect 234160 335446 234212 335452
rect 234172 7546 234200 335446
rect 234160 7540 234212 7546
rect 234160 7482 234212 7488
rect 234264 7410 234292 335582
rect 234344 335368 234396 335374
rect 234344 335310 234396 335316
rect 234356 8226 234384 335310
rect 234448 237153 234476 351727
rect 234434 237144 234490 237153
rect 234434 237079 234490 237088
rect 234540 236337 234568 362879
rect 269730 338162 269758 338164
rect 269718 338156 269770 338162
rect 269718 338098 269770 338104
rect 234724 338014 235060 338042
rect 234724 333305 234752 338014
rect 234804 337952 234856 337958
rect 235138 337906 235166 338028
rect 235230 337958 235258 338028
rect 234804 337894 234856 337900
rect 234710 333296 234766 333305
rect 234710 333231 234766 333240
rect 234526 236328 234582 236337
rect 234526 236263 234582 236272
rect 234528 80912 234580 80918
rect 234528 80854 234580 80860
rect 234344 8220 234396 8226
rect 234344 8162 234396 8168
rect 234252 7404 234304 7410
rect 234252 7346 234304 7352
rect 234068 7336 234120 7342
rect 234068 7278 234120 7284
rect 234436 4820 234488 4826
rect 234436 4762 234488 4768
rect 234448 4729 234476 4762
rect 234434 4720 234490 4729
rect 234434 4655 234490 4664
rect 234068 4140 234120 4146
rect 234068 4082 234120 4088
rect 234080 4049 234108 4082
rect 234066 4040 234122 4049
rect 234066 3975 234122 3984
rect 234540 3534 234568 80854
rect 234816 4865 234844 337894
rect 234988 337884 235040 337890
rect 234988 337826 235040 337832
rect 235092 337878 235166 337906
rect 235218 337952 235270 337958
rect 235218 337894 235270 337900
rect 235000 321554 235028 337826
rect 235092 333441 235120 337878
rect 235322 337770 235350 338028
rect 235184 337742 235350 337770
rect 235078 333432 235134 333441
rect 235078 333367 235134 333376
rect 234908 321526 235028 321554
rect 234908 177410 234936 321526
rect 235184 316034 235212 337742
rect 235414 337668 235442 338028
rect 235506 337770 235534 338028
rect 235598 337929 235626 338028
rect 235690 337958 235718 338028
rect 235678 337952 235730 337958
rect 235584 337920 235640 337929
rect 235678 337894 235730 337900
rect 235584 337855 235640 337864
rect 235630 337784 235686 337793
rect 235506 337742 235580 337770
rect 235414 337640 235488 337668
rect 235264 336796 235316 336802
rect 235264 336738 235316 336744
rect 235000 316006 235212 316034
rect 234896 177404 234948 177410
rect 234896 177346 234948 177352
rect 235000 177342 235028 316006
rect 234988 177336 235040 177342
rect 234988 177278 235040 177284
rect 235276 7614 235304 336738
rect 235356 336660 235408 336666
rect 235356 336602 235408 336608
rect 235368 331214 235396 336602
rect 235460 336054 235488 337640
rect 235552 336122 235580 337742
rect 235782 337770 235810 338028
rect 235630 337719 235686 337728
rect 235736 337742 235810 337770
rect 235874 337770 235902 338028
rect 235966 337958 235994 338028
rect 235954 337952 236006 337958
rect 235954 337894 236006 337900
rect 236058 337770 236086 338028
rect 235874 337742 235948 337770
rect 235540 336116 235592 336122
rect 235540 336058 235592 336064
rect 235448 336048 235500 336054
rect 235448 335990 235500 335996
rect 235538 335472 235594 335481
rect 235538 335407 235594 335416
rect 235368 331186 235488 331214
rect 235460 321554 235488 331186
rect 235368 321526 235488 321554
rect 235368 7682 235396 321526
rect 235552 316034 235580 335407
rect 235644 326466 235672 337719
rect 235736 335442 235764 337742
rect 235816 337680 235868 337686
rect 235816 337622 235868 337628
rect 235724 335436 235776 335442
rect 235724 335378 235776 335384
rect 235632 326460 235684 326466
rect 235632 326402 235684 326408
rect 235828 326346 235856 337622
rect 235920 335481 235948 337742
rect 236012 337742 236086 337770
rect 236196 338014 236256 338042
rect 236012 336802 236040 337742
rect 236196 336802 236224 338014
rect 236334 337770 236362 338028
rect 236288 337742 236362 337770
rect 236426 337770 236454 338028
rect 236518 337958 236546 338028
rect 236506 337952 236558 337958
rect 236506 337894 236558 337900
rect 236610 337770 236638 338028
rect 236426 337742 236500 337770
rect 236000 336796 236052 336802
rect 236000 336738 236052 336744
rect 236184 336796 236236 336802
rect 236184 336738 236236 336744
rect 236288 335753 236316 337742
rect 236472 337634 236500 337742
rect 236380 337606 236500 337634
rect 236564 337742 236638 337770
rect 236702 337770 236730 338028
rect 236794 337890 236822 338028
rect 236782 337884 236834 337890
rect 236782 337826 236834 337832
rect 236886 337770 236914 338028
rect 236978 337890 237006 338028
rect 236966 337884 237018 337890
rect 236966 337826 237018 337832
rect 236702 337742 236776 337770
rect 236274 335744 236330 335753
rect 236274 335679 236330 335688
rect 235906 335472 235962 335481
rect 235906 335407 235962 335416
rect 236000 335436 236052 335442
rect 236000 335378 236052 335384
rect 236012 335322 236040 335378
rect 235920 335294 236040 335322
rect 236184 335368 236236 335374
rect 236184 335310 236236 335316
rect 235920 334665 235948 335294
rect 235906 334656 235962 334665
rect 235906 334591 235962 334600
rect 235460 316006 235580 316034
rect 235644 326318 235856 326346
rect 235460 238921 235488 316006
rect 235446 238912 235502 238921
rect 235446 238847 235502 238856
rect 235356 7676 235408 7682
rect 235356 7618 235408 7624
rect 235264 7608 235316 7614
rect 235264 7550 235316 7556
rect 235644 4894 235672 326318
rect 235724 326256 235776 326262
rect 235724 326198 235776 326204
rect 235632 4888 235684 4894
rect 234802 4856 234858 4865
rect 234620 4820 234672 4826
rect 235632 4830 235684 4836
rect 234802 4791 234858 4800
rect 234620 4762 234672 4768
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 233976 2916 234028 2922
rect 233976 2858 234028 2864
rect 233792 2848 233844 2854
rect 233792 2790 233844 2796
rect 234632 480 234660 4762
rect 235736 4729 235764 326198
rect 236196 316034 236224 335310
rect 236288 331214 236316 335679
rect 236380 335442 236408 337606
rect 236460 337544 236512 337550
rect 236460 337486 236512 337492
rect 236368 335436 236420 335442
rect 236368 335378 236420 335384
rect 236472 331906 236500 337486
rect 236564 336258 236592 337742
rect 236644 337068 236696 337074
rect 236644 337010 236696 337016
rect 236552 336252 236604 336258
rect 236552 336194 236604 336200
rect 236656 334801 236684 337010
rect 236748 335617 236776 337742
rect 236840 337742 236914 337770
rect 237070 337770 237098 338028
rect 237162 337872 237190 338028
rect 237254 337940 237282 338028
rect 237392 338014 237452 338042
rect 237254 337912 237328 337940
rect 237162 337844 237236 337872
rect 237070 337742 237144 337770
rect 236734 335608 236790 335617
rect 236734 335543 236790 335552
rect 236642 334792 236698 334801
rect 236642 334727 236698 334736
rect 236460 331900 236512 331906
rect 236460 331842 236512 331848
rect 236288 331186 236684 331214
rect 236460 326392 236512 326398
rect 236460 326334 236512 326340
rect 236104 316006 236224 316034
rect 236104 240145 236132 316006
rect 236090 240136 236146 240145
rect 236090 240071 236146 240080
rect 235816 11756 235868 11762
rect 235816 11698 235868 11704
rect 235722 4720 235778 4729
rect 235722 4655 235778 4664
rect 235828 480 235856 11698
rect 236472 3602 236500 326334
rect 236460 3596 236512 3602
rect 236460 3538 236512 3544
rect 236656 3369 236684 331186
rect 236748 321554 236776 335543
rect 236840 330546 236868 337742
rect 236920 337680 236972 337686
rect 236920 337622 236972 337628
rect 237010 337648 237066 337657
rect 236828 330540 236880 330546
rect 236828 330482 236880 330488
rect 236932 326398 236960 337622
rect 237010 337583 237066 337592
rect 237024 336705 237052 337583
rect 237116 336954 237144 337742
rect 237208 337074 237236 337844
rect 237196 337068 237248 337074
rect 237196 337010 237248 337016
rect 237116 336926 237236 336954
rect 237104 336796 237156 336802
rect 237104 336738 237156 336744
rect 237010 336696 237066 336705
rect 237010 336631 237066 336640
rect 237012 336252 237064 336258
rect 237012 336194 237064 336200
rect 237024 333742 237052 336194
rect 237012 333736 237064 333742
rect 237012 333678 237064 333684
rect 236920 326392 236972 326398
rect 236920 326334 236972 326340
rect 236748 321526 237052 321554
rect 236826 240136 236882 240145
rect 236826 240071 236882 240080
rect 236840 238785 236868 240071
rect 237024 239057 237052 321526
rect 237010 239048 237066 239057
rect 237010 238983 237066 238992
rect 236826 238776 236882 238785
rect 236826 238711 236882 238720
rect 236840 3505 236868 238711
rect 236826 3496 236882 3505
rect 237116 3466 237144 336738
rect 237208 335374 237236 336926
rect 237300 336326 237328 337912
rect 237288 336320 237340 336326
rect 237288 336262 237340 336268
rect 237392 336025 237420 338014
rect 237530 337958 237558 338028
rect 237622 337958 237650 338028
rect 237518 337952 237570 337958
rect 237518 337894 237570 337900
rect 237610 337952 237662 337958
rect 237610 337894 237662 337900
rect 237470 337784 237526 337793
rect 237714 337770 237742 338028
rect 237470 337719 237526 337728
rect 237576 337742 237742 337770
rect 237806 337770 237834 338028
rect 237898 337890 237926 338028
rect 237886 337884 237938 337890
rect 237886 337826 237938 337832
rect 237990 337822 238018 338028
rect 237978 337816 238030 337822
rect 237806 337742 237880 337770
rect 237978 337758 238030 337764
rect 237378 336016 237434 336025
rect 237378 335951 237434 335960
rect 237286 335880 237342 335889
rect 237286 335815 237342 335824
rect 237196 335368 237248 335374
rect 237196 335310 237248 335316
rect 237300 333266 237328 335815
rect 237288 333260 237340 333266
rect 237288 333202 237340 333208
rect 237484 3806 237512 337719
rect 237472 3800 237524 3806
rect 237472 3742 237524 3748
rect 237576 3670 237604 337742
rect 237656 337680 237708 337686
rect 237852 337668 237880 337742
rect 238082 337668 238110 338028
rect 238174 337770 238202 338028
rect 238266 337929 238294 338028
rect 238252 337920 238308 337929
rect 238252 337855 238308 337864
rect 238358 337770 238386 338028
rect 238174 337742 238248 337770
rect 237656 337622 237708 337628
rect 237760 337640 237880 337668
rect 238036 337640 238110 337668
rect 237668 335889 237696 337622
rect 237760 336802 237788 337640
rect 237932 337612 237984 337618
rect 237932 337554 237984 337560
rect 237840 337000 237892 337006
rect 237840 336942 237892 336948
rect 237748 336796 237800 336802
rect 237748 336738 237800 336744
rect 237654 335880 237710 335889
rect 237654 335815 237710 335824
rect 237760 333334 237788 336738
rect 237852 336161 237880 336942
rect 237944 336297 237972 337554
rect 237930 336288 237986 336297
rect 237930 336223 237986 336232
rect 237838 336152 237894 336161
rect 238036 336138 238064 337640
rect 237838 336087 237894 336096
rect 237944 336110 238064 336138
rect 237944 334121 237972 336110
rect 238022 335608 238078 335617
rect 238220 335594 238248 337742
rect 238022 335543 238078 335552
rect 238128 335566 238248 335594
rect 238312 337742 238386 337770
rect 238496 338014 238556 338042
rect 237930 334112 237986 334121
rect 237930 334047 237986 334056
rect 237944 333402 237972 334047
rect 237932 333396 237984 333402
rect 237932 333338 237984 333344
rect 237748 333328 237800 333334
rect 237748 333270 237800 333276
rect 237656 326392 237708 326398
rect 237656 326334 237708 326340
rect 237668 3738 237696 326334
rect 237748 321836 237800 321842
rect 237748 321778 237800 321784
rect 237760 278798 237788 321778
rect 237748 278792 237800 278798
rect 237748 278734 237800 278740
rect 238036 4010 238064 335543
rect 238128 326398 238156 335566
rect 238208 333260 238260 333266
rect 238208 333202 238260 333208
rect 238116 326392 238168 326398
rect 238116 326334 238168 326340
rect 238116 278792 238168 278798
rect 238116 278734 238168 278740
rect 238128 6186 238156 278734
rect 238116 6180 238168 6186
rect 238116 6122 238168 6128
rect 238024 4004 238076 4010
rect 238024 3946 238076 3952
rect 238220 3874 238248 333202
rect 238312 331294 238340 337742
rect 238392 337680 238444 337686
rect 238392 337622 238444 337628
rect 238300 331288 238352 331294
rect 238300 331230 238352 331236
rect 238312 327758 238340 331230
rect 238300 327752 238352 327758
rect 238300 327694 238352 327700
rect 238404 4146 238432 337622
rect 238496 336190 238524 338014
rect 238634 337958 238662 338028
rect 238622 337952 238674 337958
rect 238622 337894 238674 337900
rect 238726 337770 238754 338028
rect 238818 337958 238846 338028
rect 238910 337958 238938 338028
rect 238806 337952 238858 337958
rect 238806 337894 238858 337900
rect 238898 337952 238950 337958
rect 238898 337894 238950 337900
rect 238680 337742 238754 337770
rect 238852 337816 238904 337822
rect 239002 337770 239030 338028
rect 238852 337758 238904 337764
rect 238484 336184 238536 336190
rect 238484 336126 238536 336132
rect 238576 336048 238628 336054
rect 238576 335990 238628 335996
rect 238588 334937 238616 335990
rect 238574 334928 238630 334937
rect 238574 334863 238630 334872
rect 238680 321842 238708 337742
rect 238668 321836 238720 321842
rect 238668 321778 238720 321784
rect 238392 4140 238444 4146
rect 238392 4082 238444 4088
rect 238864 3942 238892 337758
rect 238956 337742 239030 337770
rect 239094 337770 239122 338028
rect 239186 337890 239214 338028
rect 239174 337884 239226 337890
rect 239174 337826 239226 337832
rect 239278 337770 239306 338028
rect 239094 337742 239168 337770
rect 238956 333577 238984 337742
rect 239036 337680 239088 337686
rect 239036 337622 239088 337628
rect 239048 335617 239076 337622
rect 239034 335608 239090 335617
rect 239034 335543 239090 335552
rect 238942 333568 238998 333577
rect 238942 333503 238998 333512
rect 239036 333260 239088 333266
rect 239036 333202 239088 333208
rect 238944 323876 238996 323882
rect 238944 323818 238996 323824
rect 238956 6225 238984 323818
rect 239048 7750 239076 333202
rect 239140 86290 239168 337742
rect 239232 337742 239306 337770
rect 239232 333713 239260 337742
rect 239370 337668 239398 338028
rect 239462 337958 239490 338028
rect 239450 337952 239502 337958
rect 239554 337940 239582 338028
rect 239692 338014 239752 338042
rect 239554 337912 239628 337940
rect 239450 337894 239502 337900
rect 239496 337816 239548 337822
rect 239496 337758 239548 337764
rect 239324 337640 239398 337668
rect 239218 333704 239274 333713
rect 239218 333639 239274 333648
rect 239324 331214 239352 337640
rect 239508 336433 239536 337758
rect 239494 336424 239550 336433
rect 239494 336359 239550 336368
rect 239600 333849 239628 337912
rect 239586 333840 239642 333849
rect 239586 333775 239642 333784
rect 239232 331186 239352 331214
rect 239232 177478 239260 331186
rect 239692 323882 239720 338014
rect 239830 337940 239858 338028
rect 239784 337912 239858 337940
rect 239680 323876 239732 323882
rect 239680 323818 239732 323824
rect 239784 316034 239812 337912
rect 239922 337872 239950 338028
rect 239876 337844 239950 337872
rect 239876 331974 239904 337844
rect 240014 337770 240042 338028
rect 239968 337742 240042 337770
rect 239968 333266 239996 337742
rect 240106 337668 240134 338028
rect 240060 337640 240134 337668
rect 240198 337668 240226 338028
rect 240290 337770 240318 338028
rect 240382 337929 240410 338028
rect 240474 337958 240502 338028
rect 240462 337952 240514 337958
rect 240368 337920 240424 337929
rect 240462 337894 240514 337900
rect 240368 337855 240424 337864
rect 240566 337822 240594 338028
rect 240554 337816 240606 337822
rect 240414 337784 240470 337793
rect 240290 337742 240364 337770
rect 240198 337640 240272 337668
rect 240060 336569 240088 337640
rect 240046 336560 240102 336569
rect 240046 336495 240102 336504
rect 240244 333470 240272 337640
rect 240232 333464 240284 333470
rect 240232 333406 240284 333412
rect 239956 333260 240008 333266
rect 239956 333202 240008 333208
rect 239864 331968 239916 331974
rect 239864 331910 239916 331916
rect 239324 316006 239812 316034
rect 239220 177472 239272 177478
rect 239220 177414 239272 177420
rect 239128 86284 239180 86290
rect 239128 86226 239180 86232
rect 239036 7744 239088 7750
rect 239036 7686 239088 7692
rect 238942 6216 238998 6225
rect 238942 6151 238998 6160
rect 239324 4078 239352 316006
rect 240336 7818 240364 337742
rect 240554 337758 240606 337764
rect 240658 337770 240686 338028
rect 240750 337906 240778 338028
rect 240888 338014 240948 338042
rect 240750 337878 240824 337906
rect 240658 337742 240732 337770
rect 240414 337719 240470 337728
rect 240428 326398 240456 337719
rect 240508 337680 240560 337686
rect 240704 337657 240732 337742
rect 240508 337622 240560 337628
rect 240690 337648 240746 337657
rect 240416 326392 240468 326398
rect 240416 326334 240468 326340
rect 240416 326256 240468 326262
rect 240416 326198 240468 326204
rect 240428 8022 240456 326198
rect 240520 8090 240548 337622
rect 240796 337634 240824 337878
rect 240888 337754 240916 338014
rect 241026 337770 241054 338028
rect 241118 337890 241146 338028
rect 241106 337884 241158 337890
rect 241106 337826 241158 337832
rect 241210 337770 241238 338028
rect 240876 337748 240928 337754
rect 241026 337742 241100 337770
rect 240876 337690 240928 337696
rect 240796 337606 240916 337634
rect 240690 337583 240746 337592
rect 240692 337544 240744 337550
rect 240692 337486 240744 337492
rect 240704 326466 240732 337486
rect 240784 335844 240836 335850
rect 240784 335786 240836 335792
rect 240796 332110 240824 335786
rect 240888 333606 240916 337606
rect 240876 333600 240928 333606
rect 240876 333542 240928 333548
rect 240784 332104 240836 332110
rect 240784 332046 240836 332052
rect 240784 331968 240836 331974
rect 240784 331910 240836 331916
rect 240692 326460 240744 326466
rect 240692 326402 240744 326408
rect 240796 322674 240824 331910
rect 240876 326392 240928 326398
rect 240876 326334 240928 326340
rect 240612 322646 240824 322674
rect 240508 8084 240560 8090
rect 240508 8026 240560 8032
rect 240416 8016 240468 8022
rect 240416 7958 240468 7964
rect 240612 7954 240640 322646
rect 240784 322108 240836 322114
rect 240784 322050 240836 322056
rect 240692 321088 240744 321094
rect 240692 321030 240744 321036
rect 240704 80714 240732 321030
rect 240796 84862 240824 322050
rect 240888 177546 240916 326334
rect 240876 177540 240928 177546
rect 240876 177482 240928 177488
rect 240784 84856 240836 84862
rect 240784 84798 240836 84804
rect 240692 80708 240744 80714
rect 240692 80650 240744 80656
rect 240600 7948 240652 7954
rect 240600 7890 240652 7896
rect 240324 7812 240376 7818
rect 240324 7754 240376 7760
rect 239312 4072 239364 4078
rect 239312 4014 239364 4020
rect 238852 3936 238904 3942
rect 238852 3878 238904 3884
rect 238208 3868 238260 3874
rect 238208 3810 238260 3816
rect 237656 3732 237708 3738
rect 237656 3674 237708 3680
rect 237564 3664 237616 3670
rect 237564 3606 237616 3612
rect 240508 3596 240560 3602
rect 240508 3538 240560 3544
rect 238116 3528 238168 3534
rect 238116 3470 238168 3476
rect 236826 3431 236882 3440
rect 237104 3460 237156 3466
rect 237104 3402 237156 3408
rect 236642 3360 236698 3369
rect 236642 3295 236698 3304
rect 237012 2916 237064 2922
rect 237012 2858 237064 2864
rect 237024 480 237052 2858
rect 238128 480 238156 3470
rect 239312 3324 239364 3330
rect 239312 3266 239364 3272
rect 239324 480 239352 3266
rect 240520 480 240548 3538
rect 241072 2854 241100 337742
rect 241164 337742 241238 337770
rect 241164 326262 241192 337742
rect 241302 337668 241330 338028
rect 241394 337770 241422 338028
rect 241486 337890 241514 338028
rect 241474 337884 241526 337890
rect 241474 337826 241526 337832
rect 241394 337742 241468 337770
rect 241256 337640 241330 337668
rect 241256 336462 241284 337640
rect 241244 336456 241296 336462
rect 241244 336398 241296 336404
rect 241244 333260 241296 333266
rect 241244 333202 241296 333208
rect 241152 326256 241204 326262
rect 241152 326198 241204 326204
rect 241256 7886 241284 333202
rect 241440 322114 241468 337742
rect 241578 337668 241606 338028
rect 241670 337770 241698 338028
rect 241762 337958 241790 338028
rect 241854 338008 241882 338028
rect 241854 337980 241928 338008
rect 241750 337952 241802 337958
rect 241750 337894 241802 337900
rect 241670 337742 241836 337770
rect 241704 337680 241756 337686
rect 241578 337640 241652 337668
rect 241520 337544 241572 337550
rect 241520 337486 241572 337492
rect 241532 335850 241560 337486
rect 241520 335844 241572 335850
rect 241520 335786 241572 335792
rect 241624 326534 241652 337640
rect 241704 337622 241756 337628
rect 241716 336326 241744 337622
rect 241704 336320 241756 336326
rect 241704 336262 241756 336268
rect 241704 336116 241756 336122
rect 241704 336058 241756 336064
rect 241716 334286 241744 336058
rect 241704 334280 241756 334286
rect 241704 334222 241756 334228
rect 241808 331214 241836 337742
rect 241900 336598 241928 337980
rect 242038 337770 242066 338028
rect 242130 337958 242158 338028
rect 242118 337952 242170 337958
rect 242118 337894 242170 337900
rect 242222 337770 242250 338028
rect 242314 337822 242342 338028
rect 242038 337742 242112 337770
rect 241978 337648 242034 337657
rect 241978 337583 242034 337592
rect 241888 336592 241940 336598
rect 241888 336534 241940 336540
rect 241888 336320 241940 336326
rect 241888 336262 241940 336268
rect 241900 332042 241928 336262
rect 241992 335986 242020 337583
rect 241980 335980 242032 335986
rect 241980 335922 242032 335928
rect 241888 332036 241940 332042
rect 241888 331978 241940 331984
rect 241808 331186 242020 331214
rect 241612 326528 241664 326534
rect 241612 326470 241664 326476
rect 241796 326460 241848 326466
rect 241796 326402 241848 326408
rect 241704 326324 241756 326330
rect 241704 326266 241756 326272
rect 241428 322108 241480 322114
rect 241428 322050 241480 322056
rect 241244 7880 241296 7886
rect 241244 7822 241296 7828
rect 241716 6633 241744 326266
rect 241702 6624 241758 6633
rect 241702 6559 241758 6568
rect 241808 6497 241836 326402
rect 241888 326392 241940 326398
rect 241888 326334 241940 326340
rect 241794 6488 241850 6497
rect 241794 6423 241850 6432
rect 241900 6361 241928 326334
rect 241992 84930 242020 331186
rect 242084 87650 242112 337742
rect 242176 337742 242250 337770
rect 242302 337816 242354 337822
rect 242302 337758 242354 337764
rect 242176 336734 242204 337742
rect 242406 337736 242434 338028
rect 242498 337890 242526 338028
rect 242486 337884 242538 337890
rect 242486 337826 242538 337832
rect 242590 337770 242618 338028
rect 242682 337958 242710 338028
rect 242670 337952 242722 337958
rect 242670 337894 242722 337900
rect 242774 337827 242802 338028
rect 242866 337958 242894 338028
rect 242854 337952 242906 337958
rect 242854 337894 242906 337900
rect 242760 337818 242816 337827
rect 242958 337822 242986 338028
rect 242590 337742 242664 337770
rect 242760 337753 242816 337762
rect 242946 337816 242998 337822
rect 243050 337804 243078 338028
rect 243188 338014 243248 338042
rect 243188 337890 243216 338014
rect 243326 337958 243354 338028
rect 243314 337952 243366 337958
rect 243314 337894 243366 337900
rect 243176 337884 243228 337890
rect 243176 337826 243228 337832
rect 243418 337822 243446 338028
rect 243510 337958 243538 338028
rect 243498 337952 243550 337958
rect 243498 337894 243550 337900
rect 243406 337816 243458 337822
rect 243050 337776 243124 337804
rect 242946 337758 242998 337764
rect 243096 337770 243124 337776
rect 243096 337742 243216 337770
rect 243602 337804 243630 338028
rect 243406 337758 243458 337764
rect 243556 337776 243630 337804
rect 242406 337708 242480 337736
rect 242256 337680 242308 337686
rect 242256 337622 242308 337628
rect 242164 336728 242216 336734
rect 242164 336670 242216 336676
rect 242164 333260 242216 333266
rect 242164 333202 242216 333208
rect 242072 87644 242124 87650
rect 242072 87586 242124 87592
rect 241980 84924 242032 84930
rect 241980 84866 242032 84872
rect 242176 8158 242204 333202
rect 242268 326398 242296 337622
rect 242348 335844 242400 335850
rect 242348 335786 242400 335792
rect 242256 326392 242308 326398
rect 242256 326334 242308 326340
rect 242360 316034 242388 335786
rect 242452 333674 242480 337708
rect 242532 337680 242584 337686
rect 242532 337622 242584 337628
rect 242440 333668 242492 333674
rect 242440 333610 242492 333616
rect 242544 321554 242572 337622
rect 242636 326466 242664 337742
rect 243188 337668 243216 337742
rect 243096 337640 243216 337668
rect 243452 337680 243504 337686
rect 242808 337612 242860 337618
rect 242808 337554 242860 337560
rect 242716 326528 242768 326534
rect 242716 326470 242768 326476
rect 242624 326460 242676 326466
rect 242624 326402 242676 326408
rect 242544 321526 242664 321554
rect 242268 316006 242388 316034
rect 242268 8294 242296 316006
rect 242256 8288 242308 8294
rect 242256 8230 242308 8236
rect 242164 8152 242216 8158
rect 242164 8094 242216 8100
rect 241886 6352 241942 6361
rect 241886 6287 241942 6296
rect 241704 3664 241756 3670
rect 241704 3606 241756 3612
rect 241060 2848 241112 2854
rect 241060 2790 241112 2796
rect 241716 480 241744 3606
rect 242636 3398 242664 321526
rect 242728 3738 242756 326470
rect 242820 326330 242848 337554
rect 242992 336456 243044 336462
rect 242992 336398 243044 336404
rect 243004 335442 243032 336398
rect 242992 335436 243044 335442
rect 242992 335378 243044 335384
rect 243096 326466 243124 337640
rect 243452 337622 243504 337628
rect 243360 336252 243412 336258
rect 243360 336194 243412 336200
rect 243372 335889 243400 336194
rect 243358 335880 243414 335889
rect 243358 335815 243414 335824
rect 243176 335436 243228 335442
rect 243176 335378 243228 335384
rect 243084 326460 243136 326466
rect 243084 326402 243136 326408
rect 242808 326324 242860 326330
rect 242808 326266 242860 326272
rect 243084 326324 243136 326330
rect 243084 326266 243136 326272
rect 242900 4888 242952 4894
rect 242900 4830 242952 4836
rect 242716 3732 242768 3738
rect 242716 3674 242768 3680
rect 242624 3392 242676 3398
rect 242624 3334 242676 3340
rect 242912 480 242940 4830
rect 243096 3126 243124 326266
rect 243188 86358 243216 335378
rect 243268 333328 243320 333334
rect 243268 333270 243320 333276
rect 243280 177614 243308 333270
rect 243464 332178 243492 337622
rect 243556 333266 243584 337776
rect 243694 337736 243722 338028
rect 243786 337958 243814 338028
rect 243774 337952 243826 337958
rect 243774 337894 243826 337900
rect 243878 337770 243906 338028
rect 243970 337890 243998 338028
rect 243958 337884 244010 337890
rect 243958 337826 244010 337832
rect 244062 337770 244090 338028
rect 243648 337708 243722 337736
rect 243832 337742 243906 337770
rect 244016 337742 244090 337770
rect 244154 337770 244182 338028
rect 244246 337890 244274 338028
rect 244234 337884 244286 337890
rect 244234 337826 244286 337832
rect 244430 337770 244458 338028
rect 244522 337958 244550 338028
rect 244510 337952 244562 337958
rect 244510 337894 244562 337900
rect 244614 337770 244642 338028
rect 244706 337890 244734 338028
rect 244694 337884 244746 337890
rect 244694 337826 244746 337832
rect 244798 337822 244826 338028
rect 244890 337890 244918 338028
rect 244982 337963 245010 338028
rect 244968 337954 245024 337963
rect 245074 337958 245102 338028
rect 245166 337958 245194 338028
rect 244878 337884 244930 337890
rect 244968 337889 245024 337898
rect 245062 337952 245114 337958
rect 245062 337894 245114 337900
rect 245154 337952 245206 337958
rect 245154 337894 245206 337900
rect 244878 337826 244930 337832
rect 244786 337816 244838 337822
rect 244154 337742 244228 337770
rect 244430 337742 244504 337770
rect 244614 337742 244688 337770
rect 244786 337758 244838 337764
rect 244968 337784 245024 337793
rect 243544 333260 243596 333266
rect 243544 333202 243596 333208
rect 243452 332172 243504 332178
rect 243452 332114 243504 332120
rect 243360 326392 243412 326398
rect 243360 326334 243412 326340
rect 243372 177682 243400 326334
rect 243648 316034 243676 337708
rect 243726 337648 243782 337657
rect 243726 337583 243782 337592
rect 243740 333810 243768 337583
rect 243832 335986 243860 337742
rect 243912 337680 243964 337686
rect 243912 337622 243964 337628
rect 243820 335980 243872 335986
rect 243820 335922 243872 335928
rect 243924 335918 243952 337622
rect 243912 335912 243964 335918
rect 243912 335854 243964 335860
rect 243728 333804 243780 333810
rect 243728 333746 243780 333752
rect 243912 326460 243964 326466
rect 243912 326402 243964 326408
rect 243464 316006 243676 316034
rect 243360 177676 243412 177682
rect 243360 177618 243412 177624
rect 243268 177608 243320 177614
rect 243268 177550 243320 177556
rect 243176 86352 243228 86358
rect 243176 86294 243228 86300
rect 243464 3194 243492 316006
rect 243924 3262 243952 326402
rect 244016 326398 244044 337742
rect 244096 337680 244148 337686
rect 244096 337622 244148 337628
rect 244108 331214 244136 337622
rect 244200 335850 244228 337742
rect 244280 336524 244332 336530
rect 244280 336466 244332 336472
rect 244188 335844 244240 335850
rect 244188 335786 244240 335792
rect 244292 334762 244320 336466
rect 244372 335980 244424 335986
rect 244372 335922 244424 335928
rect 244280 334756 244332 334762
rect 244280 334698 244332 334704
rect 244108 331186 244228 331214
rect 244004 326392 244056 326398
rect 244004 326334 244056 326340
rect 244200 326330 244228 331186
rect 244188 326324 244240 326330
rect 244188 326266 244240 326272
rect 244096 3732 244148 3738
rect 244096 3674 244148 3680
rect 243912 3256 243964 3262
rect 243912 3198 243964 3204
rect 243452 3188 243504 3194
rect 243452 3130 243504 3136
rect 243084 3120 243136 3126
rect 243084 3062 243136 3068
rect 244108 480 244136 3674
rect 244384 3534 244412 335922
rect 244476 326262 244504 337742
rect 244556 337680 244608 337686
rect 244556 337622 244608 337628
rect 244568 335646 244596 337622
rect 244660 335714 244688 337742
rect 245258 337770 245286 338028
rect 245350 337958 245378 338028
rect 245488 338014 245548 338042
rect 245338 337952 245390 337958
rect 245338 337894 245390 337900
rect 245488 337822 245516 338014
rect 245626 337822 245654 338028
rect 245718 337963 245746 338028
rect 245704 337954 245760 337963
rect 245704 337889 245760 337898
rect 245810 337822 245838 338028
rect 245902 337963 245930 338028
rect 245888 337954 245944 337963
rect 245888 337889 245944 337898
rect 245476 337816 245528 337822
rect 245258 337742 245332 337770
rect 245476 337758 245528 337764
rect 245614 337816 245666 337822
rect 245614 337758 245666 337764
rect 245798 337816 245850 337822
rect 245994 337770 246022 338028
rect 245798 337758 245850 337764
rect 245024 337728 245056 337736
rect 244968 337719 245056 337728
rect 244982 337708 245056 337719
rect 244740 337680 244792 337686
rect 244740 337622 244792 337628
rect 244832 337680 244884 337686
rect 244832 337622 244884 337628
rect 244648 335708 244700 335714
rect 244648 335650 244700 335656
rect 244556 335640 244608 335646
rect 244556 335582 244608 335588
rect 244648 326800 244700 326806
rect 244648 326742 244700 326748
rect 244556 326460 244608 326466
rect 244556 326402 244608 326408
rect 244464 326256 244516 326262
rect 244464 326198 244516 326204
rect 244464 326120 244516 326126
rect 244464 326062 244516 326068
rect 244476 6322 244504 326062
rect 244464 6316 244516 6322
rect 244464 6258 244516 6264
rect 244568 6254 244596 326402
rect 244660 7478 244688 326742
rect 244752 326738 244780 337622
rect 244844 326806 244872 337622
rect 244924 333804 244976 333810
rect 244924 333746 244976 333752
rect 244832 326800 244884 326806
rect 244832 326742 244884 326748
rect 244740 326732 244792 326738
rect 244740 326674 244792 326680
rect 244832 326528 244884 326534
rect 244832 326470 244884 326476
rect 244740 326256 244792 326262
rect 244740 326198 244792 326204
rect 244752 84998 244780 326198
rect 244844 87718 244872 326470
rect 244936 326346 244964 333746
rect 245028 326466 245056 337708
rect 245200 337612 245252 337618
rect 245200 337554 245252 337560
rect 245108 335708 245160 335714
rect 245108 335650 245160 335656
rect 245120 335170 245148 335650
rect 245108 335164 245160 335170
rect 245108 335106 245160 335112
rect 245108 334756 245160 334762
rect 245108 334698 245160 334704
rect 245120 326482 245148 334698
rect 245212 327026 245240 337554
rect 245304 328454 245332 337742
rect 245948 337742 246022 337770
rect 245842 337648 245898 337657
rect 245842 337583 245898 337592
rect 245568 336388 245620 336394
rect 245568 336330 245620 336336
rect 245384 335640 245436 335646
rect 245384 335582 245436 335588
rect 245396 332994 245424 335582
rect 245580 334150 245608 336330
rect 245856 334966 245884 337583
rect 245844 334960 245896 334966
rect 245844 334902 245896 334908
rect 245568 334144 245620 334150
rect 245568 334086 245620 334092
rect 245384 332988 245436 332994
rect 245384 332930 245436 332936
rect 245304 328426 245516 328454
rect 245212 326998 245424 327026
rect 245016 326460 245068 326466
rect 245120 326454 245332 326482
rect 245016 326402 245068 326408
rect 244936 326318 245056 326346
rect 244924 326052 244976 326058
rect 244924 325994 244976 326000
rect 244832 87712 244884 87718
rect 244832 87654 244884 87660
rect 244740 84992 244792 84998
rect 244740 84934 244792 84940
rect 244648 7472 244700 7478
rect 244648 7414 244700 7420
rect 244556 6248 244608 6254
rect 244556 6190 244608 6196
rect 244372 3528 244424 3534
rect 244372 3470 244424 3476
rect 244936 3330 244964 325994
rect 245028 321554 245056 326318
rect 245304 326058 245332 326454
rect 245292 326052 245344 326058
rect 245292 325994 245344 326000
rect 245028 321526 245332 321554
rect 245200 3528 245252 3534
rect 245200 3470 245252 3476
rect 244924 3324 244976 3330
rect 244924 3266 244976 3272
rect 245212 480 245240 3470
rect 245304 3058 245332 321526
rect 245292 3052 245344 3058
rect 245292 2994 245344 3000
rect 245396 2990 245424 326998
rect 245488 326126 245516 328426
rect 245844 326732 245896 326738
rect 245844 326674 245896 326680
rect 245476 326120 245528 326126
rect 245476 326062 245528 326068
rect 245856 5137 245884 326674
rect 245948 326618 245976 337742
rect 246086 337668 246114 338028
rect 246040 337640 246114 337668
rect 246178 337668 246206 338028
rect 246270 337770 246298 338028
rect 246362 337890 246390 338028
rect 246350 337884 246402 337890
rect 246350 337826 246402 337832
rect 246454 337770 246482 338028
rect 246546 337890 246574 338028
rect 246684 338014 246744 338042
rect 246534 337884 246586 337890
rect 246534 337826 246586 337832
rect 246270 337742 246344 337770
rect 246454 337742 246620 337770
rect 246178 337640 246252 337668
rect 246040 326738 246068 337640
rect 246224 335209 246252 337640
rect 246210 335200 246266 335209
rect 246210 335135 246266 335144
rect 246028 326732 246080 326738
rect 246028 326674 246080 326680
rect 245948 326590 246252 326618
rect 246120 326460 246172 326466
rect 246120 326402 246172 326408
rect 246028 326256 246080 326262
rect 246028 326198 246080 326204
rect 245936 326188 245988 326194
rect 245936 326130 245988 326136
rect 245842 5128 245898 5137
rect 245842 5063 245898 5072
rect 245948 4962 245976 326130
rect 246040 6526 246068 326198
rect 246028 6520 246080 6526
rect 246028 6462 246080 6468
rect 246132 6390 246160 326402
rect 246224 326210 246252 326590
rect 246316 326346 246344 337742
rect 246396 337680 246448 337686
rect 246396 337622 246448 337628
rect 246488 337680 246540 337686
rect 246488 337622 246540 337628
rect 246408 326466 246436 337622
rect 246396 326460 246448 326466
rect 246396 326402 246448 326408
rect 246316 326318 246436 326346
rect 246224 326182 246344 326210
rect 246212 326120 246264 326126
rect 246212 326062 246264 326068
rect 246224 6458 246252 326062
rect 246316 80782 246344 326182
rect 246408 83502 246436 326318
rect 246396 83496 246448 83502
rect 246396 83438 246448 83444
rect 246304 80776 246356 80782
rect 246304 80718 246356 80724
rect 246212 6452 246264 6458
rect 246212 6394 246264 6400
rect 246120 6384 246172 6390
rect 246120 6326 246172 6332
rect 246500 5273 246528 337622
rect 246592 335345 246620 337742
rect 246578 335336 246634 335345
rect 246578 335271 246634 335280
rect 246580 333260 246632 333266
rect 246580 333202 246632 333208
rect 246486 5264 246542 5273
rect 246486 5199 246542 5208
rect 246592 5001 246620 333202
rect 246684 326126 246712 338014
rect 246822 337940 246850 338028
rect 246776 337912 246850 337940
rect 246776 332314 246804 337912
rect 246914 337872 246942 338028
rect 246868 337844 246942 337872
rect 246764 332308 246816 332314
rect 246764 332250 246816 332256
rect 246868 326194 246896 337844
rect 247006 337770 247034 338028
rect 247098 337822 247126 338028
rect 246960 337742 247034 337770
rect 247086 337816 247138 337822
rect 247086 337758 247138 337764
rect 247190 337770 247218 338028
rect 247282 337890 247310 338028
rect 247374 337958 247402 338028
rect 247362 337952 247414 337958
rect 247362 337894 247414 337900
rect 247466 337890 247494 338028
rect 247270 337884 247322 337890
rect 247270 337826 247322 337832
rect 247454 337884 247506 337890
rect 247454 337826 247506 337832
rect 247406 337784 247462 337793
rect 247190 337742 247264 337770
rect 246960 326262 246988 337742
rect 247040 337680 247092 337686
rect 247040 337622 247092 337628
rect 247052 334529 247080 337622
rect 247038 334520 247094 334529
rect 247038 334455 247094 334464
rect 247236 333878 247264 337742
rect 247558 337770 247586 338028
rect 247650 337822 247678 338028
rect 247788 338014 247848 338042
rect 247788 337890 247816 338014
rect 247776 337884 247828 337890
rect 247776 337826 247828 337832
rect 247406 337719 247462 337728
rect 247512 337742 247586 337770
rect 247638 337816 247690 337822
rect 247638 337758 247690 337764
rect 247774 337784 247830 337793
rect 247316 337680 247368 337686
rect 247316 337622 247368 337628
rect 247224 333872 247276 333878
rect 247224 333814 247276 333820
rect 247328 333198 247356 337622
rect 247420 334694 247448 337719
rect 247512 334778 247540 337742
rect 247926 337770 247954 338028
rect 248018 337793 248046 338028
rect 248110 337890 248138 338028
rect 248202 337958 248230 338028
rect 248294 337963 248322 338028
rect 248190 337952 248242 337958
rect 248190 337894 248242 337900
rect 248280 337954 248336 337963
rect 248098 337884 248150 337890
rect 248280 337889 248336 337898
rect 248386 337890 248414 338028
rect 248098 337826 248150 337832
rect 248374 337884 248426 337890
rect 248374 337826 248426 337832
rect 247774 337719 247830 337728
rect 247880 337742 247954 337770
rect 248004 337784 248060 337793
rect 247788 335646 247816 337719
rect 247776 335640 247828 335646
rect 247776 335582 247828 335588
rect 247512 334750 247816 334778
rect 247408 334688 247460 334694
rect 247408 334630 247460 334636
rect 247592 334620 247644 334626
rect 247592 334562 247644 334568
rect 247316 333192 247368 333198
rect 247316 333134 247368 333140
rect 247408 333192 247460 333198
rect 247408 333134 247460 333140
rect 247316 326460 247368 326466
rect 247316 326402 247368 326408
rect 246948 326256 247000 326262
rect 246948 326198 247000 326204
rect 246856 326188 246908 326194
rect 246856 326130 246908 326136
rect 246672 326120 246724 326126
rect 246672 326062 246724 326068
rect 247224 324420 247276 324426
rect 247224 324362 247276 324368
rect 247236 6730 247264 324362
rect 247328 6798 247356 326402
rect 247420 80850 247448 333134
rect 247500 326392 247552 326398
rect 247500 326334 247552 326340
rect 247512 83570 247540 326334
rect 247500 83564 247552 83570
rect 247500 83506 247552 83512
rect 247408 80844 247460 80850
rect 247408 80786 247460 80792
rect 247316 6792 247368 6798
rect 247316 6734 247368 6740
rect 247224 6724 247276 6730
rect 247224 6666 247276 6672
rect 247604 6594 247632 334562
rect 247788 6662 247816 334750
rect 247880 324426 247908 337742
rect 248478 337770 248506 338028
rect 248570 337890 248598 338028
rect 248558 337884 248610 337890
rect 248558 337826 248610 337832
rect 248662 337770 248690 338028
rect 248754 337872 248782 338028
rect 248846 337940 248874 338028
rect 248984 338014 249044 338042
rect 248846 337912 248920 337940
rect 248754 337844 248828 337872
rect 248004 337719 248060 337728
rect 248328 337748 248380 337754
rect 248478 337742 248552 337770
rect 248662 337742 248736 337770
rect 248328 337690 248380 337696
rect 247960 337680 248012 337686
rect 247960 337622 248012 337628
rect 247972 333130 248000 337622
rect 248144 337612 248196 337618
rect 248144 337554 248196 337560
rect 247960 333124 248012 333130
rect 247960 333066 248012 333072
rect 248156 326466 248184 337554
rect 248144 326460 248196 326466
rect 248144 326402 248196 326408
rect 248340 326398 248368 337690
rect 248420 337680 248472 337686
rect 248420 337622 248472 337628
rect 248432 332382 248460 337622
rect 248420 332376 248472 332382
rect 248420 332318 248472 332324
rect 248328 326392 248380 326398
rect 248328 326334 248380 326340
rect 248524 326126 248552 337742
rect 248708 326602 248736 337742
rect 248800 334626 248828 337844
rect 248892 336326 248920 337912
rect 248880 336320 248932 336326
rect 248880 336262 248932 336268
rect 248788 334620 248840 334626
rect 248788 334562 248840 334568
rect 248984 331786 249012 338014
rect 249122 337940 249150 338028
rect 248800 331758 249012 331786
rect 249076 337912 249150 337940
rect 248696 326596 248748 326602
rect 248696 326538 248748 326544
rect 248800 326482 248828 331758
rect 248972 331696 249024 331702
rect 248972 331638 249024 331644
rect 248880 331628 248932 331634
rect 248880 331570 248932 331576
rect 248616 326454 248828 326482
rect 248512 326120 248564 326126
rect 248512 326062 248564 326068
rect 247868 324420 247920 324426
rect 247868 324362 247920 324368
rect 247776 6656 247828 6662
rect 247776 6598 247828 6604
rect 247592 6588 247644 6594
rect 247592 6530 247644 6536
rect 248616 5098 248644 326454
rect 248696 326392 248748 326398
rect 248892 326346 248920 331570
rect 248696 326334 248748 326340
rect 248708 5438 248736 326334
rect 248800 326318 248920 326346
rect 248696 5432 248748 5438
rect 248696 5374 248748 5380
rect 248800 5302 248828 326318
rect 248880 326256 248932 326262
rect 248880 326198 248932 326204
rect 248788 5296 248840 5302
rect 248788 5238 248840 5244
rect 248892 5166 248920 326198
rect 248984 5234 249012 331638
rect 249076 326262 249104 337912
rect 249214 337872 249242 338028
rect 249168 337844 249242 337872
rect 249168 336530 249196 337844
rect 249306 337770 249334 338028
rect 249260 337742 249334 337770
rect 249156 336524 249208 336530
rect 249156 336466 249208 336472
rect 249156 335776 249208 335782
rect 249156 335718 249208 335724
rect 249168 334218 249196 335718
rect 249156 334212 249208 334218
rect 249156 334154 249208 334160
rect 249154 334112 249210 334121
rect 249154 334047 249210 334056
rect 249168 331214 249196 334047
rect 249260 331702 249288 337742
rect 249398 337668 249426 338028
rect 249352 337640 249426 337668
rect 249248 331696 249300 331702
rect 249248 331638 249300 331644
rect 249352 331634 249380 337640
rect 249490 337498 249518 338028
rect 249582 337668 249610 338028
rect 249674 337770 249702 338028
rect 249766 337958 249794 338028
rect 249858 337958 249886 338028
rect 249754 337952 249806 337958
rect 249754 337894 249806 337900
rect 249846 337952 249898 337958
rect 249846 337894 249898 337900
rect 249950 337872 249978 338028
rect 250042 337940 250070 338028
rect 250042 337912 250116 337940
rect 249950 337844 250024 337872
rect 249674 337742 249748 337770
rect 249582 337640 249656 337668
rect 249490 337470 249564 337498
rect 249432 334620 249484 334626
rect 249432 334562 249484 334568
rect 249340 331628 249392 331634
rect 249340 331570 249392 331576
rect 249168 331186 249288 331214
rect 249156 326596 249208 326602
rect 249156 326538 249208 326544
rect 249064 326256 249116 326262
rect 249064 326198 249116 326204
rect 249064 326120 249116 326126
rect 249064 326062 249116 326068
rect 249076 6866 249104 326062
rect 249168 85066 249196 326538
rect 249260 271862 249288 331186
rect 249248 271856 249300 271862
rect 249248 271798 249300 271804
rect 249156 85060 249208 85066
rect 249156 85002 249208 85008
rect 249064 6860 249116 6866
rect 249064 6802 249116 6808
rect 248972 5228 249024 5234
rect 248972 5170 249024 5176
rect 248880 5160 248932 5166
rect 248880 5102 248932 5108
rect 248604 5092 248656 5098
rect 248604 5034 248656 5040
rect 249444 5030 249472 334562
rect 249536 334082 249564 337470
rect 249524 334076 249576 334082
rect 249524 334018 249576 334024
rect 249628 5370 249656 337640
rect 249720 326398 249748 337742
rect 249708 326392 249760 326398
rect 249708 326334 249760 326340
rect 249996 5506 250024 337844
rect 250088 337754 250116 337912
rect 250226 337822 250254 338028
rect 250214 337816 250266 337822
rect 250214 337758 250266 337764
rect 250318 337770 250346 338028
rect 250410 337890 250438 338028
rect 250502 337963 250530 338028
rect 250488 337954 250544 337963
rect 250398 337884 250450 337890
rect 250488 337889 250544 337898
rect 250398 337826 250450 337832
rect 250594 337804 250622 338028
rect 250686 337963 250714 338028
rect 250672 337954 250728 337963
rect 250778 337958 250806 338028
rect 250870 337958 250898 338028
rect 250672 337889 250728 337898
rect 250766 337952 250818 337958
rect 250766 337894 250818 337900
rect 250858 337952 250910 337958
rect 250858 337894 250910 337900
rect 250812 337816 250864 337822
rect 250442 337784 250498 337793
rect 250076 337748 250128 337754
rect 250318 337742 250392 337770
rect 250076 337690 250128 337696
rect 250260 337680 250312 337686
rect 250260 337622 250312 337628
rect 250076 337612 250128 337618
rect 250076 337554 250128 337560
rect 249984 5500 250036 5506
rect 249984 5442 250036 5448
rect 249616 5364 249668 5370
rect 249616 5306 249668 5312
rect 249432 5024 249484 5030
rect 246578 4992 246634 5001
rect 245936 4956 245988 4962
rect 245936 4898 245988 4904
rect 246396 4956 246448 4962
rect 249432 4966 249484 4972
rect 246578 4927 246634 4936
rect 246396 4898 246448 4904
rect 245384 2984 245436 2990
rect 245384 2926 245436 2932
rect 246408 480 246436 4898
rect 250088 4554 250116 337554
rect 250168 333192 250220 333198
rect 250168 333134 250220 333140
rect 250180 4622 250208 333134
rect 250272 332926 250300 337622
rect 250260 332920 250312 332926
rect 250260 332862 250312 332868
rect 250260 326460 250312 326466
rect 250260 326402 250312 326408
rect 250272 6118 250300 326402
rect 250364 326398 250392 337742
rect 250594 337776 250760 337804
rect 250442 337719 250498 337728
rect 250352 326392 250404 326398
rect 250352 326334 250404 326340
rect 250352 326256 250404 326262
rect 250352 326198 250404 326204
rect 250260 6112 250312 6118
rect 250260 6054 250312 6060
rect 250364 6050 250392 326198
rect 250456 82142 250484 337719
rect 250536 336184 250588 336190
rect 250536 336126 250588 336132
rect 250444 82136 250496 82142
rect 250444 82078 250496 82084
rect 250548 11762 250576 336126
rect 250628 326392 250680 326398
rect 250628 326334 250680 326340
rect 250536 11756 250588 11762
rect 250536 11698 250588 11704
rect 250352 6044 250404 6050
rect 250352 5986 250404 5992
rect 250640 4758 250668 326334
rect 250628 4752 250680 4758
rect 250628 4694 250680 4700
rect 250732 4690 250760 337776
rect 250962 337770 250990 338028
rect 251054 337890 251082 338028
rect 251042 337884 251094 337890
rect 251042 337826 251094 337832
rect 251146 337770 251174 338028
rect 250812 337758 250864 337764
rect 250824 326466 250852 337758
rect 250916 337742 250990 337770
rect 251100 337742 251174 337770
rect 251284 338014 251344 338042
rect 251284 337754 251312 338014
rect 251422 337770 251450 338028
rect 251514 337958 251542 338028
rect 251606 337963 251634 338028
rect 251502 337952 251554 337958
rect 251502 337894 251554 337900
rect 251592 337954 251648 337963
rect 251592 337889 251648 337898
rect 251698 337890 251726 338028
rect 251686 337884 251738 337890
rect 251686 337826 251738 337832
rect 251546 337784 251602 337793
rect 251272 337748 251324 337754
rect 250916 335034 250944 337742
rect 250904 335028 250956 335034
rect 250904 334970 250956 334976
rect 250812 326460 250864 326466
rect 250812 326402 250864 326408
rect 251100 326262 251128 337742
rect 251422 337742 251496 337770
rect 251272 337690 251324 337696
rect 251270 337648 251326 337657
rect 251270 337583 251326 337592
rect 251180 336524 251232 336530
rect 251180 336466 251232 336472
rect 251192 332654 251220 336466
rect 251180 332648 251232 332654
rect 251180 332590 251232 332596
rect 251284 328454 251312 337583
rect 251364 334824 251416 334830
rect 251364 334766 251416 334772
rect 251376 334422 251404 334766
rect 251364 334416 251416 334422
rect 251364 334358 251416 334364
rect 251284 328426 251404 328454
rect 251088 326256 251140 326262
rect 251088 326198 251140 326204
rect 250720 4684 250772 4690
rect 250720 4626 250772 4632
rect 250168 4616 250220 4622
rect 250168 4558 250220 4564
rect 250076 4548 250128 4554
rect 250076 4490 250128 4496
rect 251376 4350 251404 328426
rect 251468 4486 251496 337742
rect 251790 337736 251818 338028
rect 251882 337770 251910 338028
rect 251974 337963 252002 338028
rect 251960 337954 252016 337963
rect 251960 337889 252016 337898
rect 252066 337890 252094 338028
rect 252054 337884 252106 337890
rect 252054 337826 252106 337832
rect 252158 337770 252186 338028
rect 251882 337742 251956 337770
rect 251546 337719 251602 337728
rect 251560 335102 251588 337719
rect 251744 337708 251818 337736
rect 251640 337544 251692 337550
rect 251640 337486 251692 337492
rect 251548 335096 251600 335102
rect 251548 335038 251600 335044
rect 251548 326392 251600 326398
rect 251548 326334 251600 326340
rect 251560 5982 251588 326334
rect 251652 86426 251680 337486
rect 251744 87786 251772 337708
rect 251824 337612 251876 337618
rect 251824 337554 251876 337560
rect 251836 89010 251864 337554
rect 251928 335238 251956 337742
rect 252112 337742 252186 337770
rect 251916 335232 251968 335238
rect 251916 335174 251968 335180
rect 252112 334490 252140 337742
rect 252250 337668 252278 338028
rect 252342 337736 252370 338028
rect 252480 338014 252540 338042
rect 252342 337708 252416 337736
rect 252204 337640 252278 337668
rect 252100 334484 252152 334490
rect 252100 334426 252152 334432
rect 251916 334416 251968 334422
rect 251916 334358 251968 334364
rect 251824 89004 251876 89010
rect 251824 88946 251876 88952
rect 251732 87780 251784 87786
rect 251732 87722 251784 87728
rect 251640 86420 251692 86426
rect 251640 86362 251692 86368
rect 251548 5976 251600 5982
rect 251548 5918 251600 5924
rect 251456 4480 251508 4486
rect 251456 4422 251508 4428
rect 251364 4344 251416 4350
rect 251364 4286 251416 4292
rect 247592 3800 247644 3806
rect 247592 3742 247644 3748
rect 247604 480 247632 3742
rect 251928 3738 251956 334358
rect 252100 332648 252152 332654
rect 252100 332590 252152 332596
rect 252112 316034 252140 332590
rect 252020 316006 252140 316034
rect 251916 3732 251968 3738
rect 251916 3674 251968 3680
rect 252020 3670 252048 316006
rect 252204 4282 252232 337640
rect 252388 334642 252416 337708
rect 252480 334830 252508 338014
rect 252618 337958 252646 338028
rect 252606 337952 252658 337958
rect 252606 337894 252658 337900
rect 252710 337736 252738 338028
rect 252802 337890 252830 338028
rect 252790 337884 252842 337890
rect 252790 337826 252842 337832
rect 252894 337770 252922 338028
rect 252664 337708 252738 337736
rect 252848 337742 252922 337770
rect 252560 336048 252612 336054
rect 252560 335990 252612 335996
rect 252468 334824 252520 334830
rect 252468 334766 252520 334772
rect 252388 334614 252508 334642
rect 252376 333192 252428 333198
rect 252376 333134 252428 333140
rect 252388 16574 252416 333134
rect 252480 326398 252508 334614
rect 252572 331974 252600 335990
rect 252560 331968 252612 331974
rect 252560 331910 252612 331916
rect 252468 326392 252520 326398
rect 252468 326334 252520 326340
rect 252664 326262 252692 337708
rect 252744 326460 252796 326466
rect 252744 326402 252796 326408
rect 252652 326256 252704 326262
rect 252652 326198 252704 326204
rect 252756 326210 252784 326402
rect 252848 326398 252876 337742
rect 252986 337668 253014 338028
rect 253078 337890 253106 338028
rect 253066 337884 253118 337890
rect 253066 337826 253118 337832
rect 253170 337770 253198 338028
rect 252940 337640 253014 337668
rect 253124 337742 253198 337770
rect 253262 337770 253290 338028
rect 253354 337890 253382 338028
rect 253342 337884 253394 337890
rect 253342 337826 253394 337832
rect 253446 337770 253474 338028
rect 253262 337742 253336 337770
rect 252836 326392 252888 326398
rect 252836 326334 252888 326340
rect 252756 326182 252876 326210
rect 252744 326120 252796 326126
rect 252744 326062 252796 326068
rect 252468 84992 252520 84998
rect 252468 84934 252520 84940
rect 252296 16546 252416 16574
rect 252296 4418 252324 16546
rect 252480 11778 252508 84934
rect 252388 11750 252508 11778
rect 252284 4412 252336 4418
rect 252284 4354 252336 4360
rect 252192 4276 252244 4282
rect 252192 4218 252244 4224
rect 252008 3664 252060 3670
rect 252008 3606 252060 3612
rect 251180 3392 251232 3398
rect 251180 3334 251232 3340
rect 249984 3052 250036 3058
rect 249984 2994 250036 3000
rect 248788 2916 248840 2922
rect 248788 2858 248840 2864
rect 248800 480 248828 2858
rect 249996 480 250024 2994
rect 251192 480 251220 3334
rect 252388 480 252416 11750
rect 252468 8900 252520 8906
rect 252468 8842 252520 8848
rect 252480 3058 252508 8842
rect 252756 5778 252784 326062
rect 252848 5846 252876 326182
rect 252940 5914 252968 337640
rect 253020 326392 253072 326398
rect 253020 326334 253072 326340
rect 253032 85134 253060 326334
rect 253124 86494 253152 337742
rect 253204 337680 253256 337686
rect 253204 337622 253256 337628
rect 253216 335306 253244 337622
rect 253204 335300 253256 335306
rect 253204 335242 253256 335248
rect 253308 326466 253336 337742
rect 253400 337742 253474 337770
rect 253296 326460 253348 326466
rect 253296 326402 253348 326408
rect 253400 326346 253428 337742
rect 253538 337736 253566 338028
rect 253676 338014 253736 338042
rect 253538 337708 253612 337736
rect 253478 337512 253534 337521
rect 253478 337447 253534 337456
rect 253492 335986 253520 337447
rect 253480 335980 253532 335986
rect 253480 335922 253532 335928
rect 253584 334234 253612 337708
rect 253676 334354 253704 338014
rect 253814 337940 253842 338028
rect 253768 337912 253842 337940
rect 253664 334348 253716 334354
rect 253664 334290 253716 334296
rect 253584 334206 253704 334234
rect 253572 334144 253624 334150
rect 253572 334086 253624 334092
rect 253216 326318 253428 326346
rect 253216 89146 253244 326318
rect 253296 326256 253348 326262
rect 253296 326198 253348 326204
rect 253204 89140 253256 89146
rect 253204 89082 253256 89088
rect 253308 89078 253336 326198
rect 253584 316034 253612 334086
rect 253676 326126 253704 334206
rect 253768 334150 253796 337912
rect 253906 337872 253934 338028
rect 253860 337844 253934 337872
rect 253756 334144 253808 334150
rect 253756 334086 253808 334092
rect 253664 326120 253716 326126
rect 253664 326062 253716 326068
rect 253860 316034 253888 337844
rect 253998 337736 254026 338028
rect 254090 337822 254118 338028
rect 254182 337963 254210 338028
rect 254168 337954 254224 337963
rect 254274 337958 254302 338028
rect 254168 337889 254224 337898
rect 254262 337952 254314 337958
rect 254262 337894 254314 337900
rect 254078 337816 254130 337822
rect 254366 337770 254394 338028
rect 254458 337890 254486 338028
rect 254446 337884 254498 337890
rect 254446 337826 254498 337832
rect 254078 337758 254130 337764
rect 253952 337708 254026 337736
rect 254320 337742 254394 337770
rect 253952 336394 253980 337708
rect 254214 337648 254270 337657
rect 254214 337583 254270 337592
rect 253940 336388 253992 336394
rect 253940 336330 253992 336336
rect 254124 326392 254176 326398
rect 254228 326380 254256 337583
rect 254320 332722 254348 337742
rect 254550 337736 254578 338028
rect 254504 337708 254578 337736
rect 254400 337680 254452 337686
rect 254400 337622 254452 337628
rect 254308 332716 254360 332722
rect 254308 332658 254360 332664
rect 254412 326505 254440 337622
rect 254504 336530 254532 337708
rect 254642 337668 254670 338028
rect 254596 337640 254670 337668
rect 254780 338014 254840 338042
rect 254492 336524 254544 336530
rect 254492 336466 254544 336472
rect 254596 331214 254624 337640
rect 254504 331186 254624 331214
rect 254398 326496 254454 326505
rect 254398 326431 254454 326440
rect 254504 326380 254532 331186
rect 254780 326398 254808 338014
rect 254918 337958 254946 338028
rect 254906 337952 254958 337958
rect 254906 337894 254958 337900
rect 255010 337770 255038 338028
rect 255102 337958 255130 338028
rect 255090 337952 255142 337958
rect 255090 337894 255142 337900
rect 254872 337742 255038 337770
rect 254228 326352 254348 326380
rect 254124 326334 254176 326340
rect 253492 316006 253612 316034
rect 253676 316006 253888 316034
rect 253296 89072 253348 89078
rect 253296 89014 253348 89020
rect 253388 88732 253440 88738
rect 253388 88674 253440 88680
rect 253204 88324 253256 88330
rect 253204 88266 253256 88272
rect 253112 86488 253164 86494
rect 253112 86430 253164 86436
rect 253020 85128 253072 85134
rect 253020 85070 253072 85076
rect 252928 5908 252980 5914
rect 252928 5850 252980 5856
rect 252836 5840 252888 5846
rect 252836 5782 252888 5788
rect 252744 5772 252796 5778
rect 252744 5714 252796 5720
rect 252468 3052 252520 3058
rect 252468 2994 252520 3000
rect 253216 2990 253244 88266
rect 253400 16574 253428 88674
rect 253308 16546 253428 16574
rect 253204 2984 253256 2990
rect 253204 2926 253256 2932
rect 253308 2922 253336 16546
rect 253492 11778 253520 316006
rect 253400 11750 253520 11778
rect 253400 4214 253428 11750
rect 253480 9172 253532 9178
rect 253480 9114 253532 9120
rect 253388 4208 253440 4214
rect 253388 4150 253440 4156
rect 253296 2916 253348 2922
rect 253296 2858 253348 2864
rect 253492 480 253520 9114
rect 253676 5710 253704 316006
rect 253664 5704 253716 5710
rect 253664 5646 253716 5652
rect 254136 4826 254164 326334
rect 254214 326224 254270 326233
rect 254214 326159 254270 326168
rect 254228 5574 254256 326159
rect 254320 5642 254348 326352
rect 254412 326352 254532 326380
rect 254768 326392 254820 326398
rect 254412 80918 254440 326352
rect 254768 326334 254820 326340
rect 254872 326108 254900 337742
rect 255194 337736 255222 338028
rect 255148 337708 255222 337736
rect 254952 337680 255004 337686
rect 254952 337622 255004 337628
rect 255044 337680 255096 337686
rect 255044 337622 255096 337628
rect 254964 336190 254992 337622
rect 254952 336184 255004 336190
rect 254952 336126 255004 336132
rect 254952 335640 255004 335646
rect 254952 335582 255004 335588
rect 254964 334762 254992 335582
rect 254952 334756 255004 334762
rect 254952 334698 255004 334704
rect 254504 326080 254900 326108
rect 254504 88330 254532 326080
rect 254676 325984 254728 325990
rect 254676 325926 254728 325932
rect 254492 88324 254544 88330
rect 254492 88266 254544 88272
rect 254400 80912 254452 80918
rect 254400 80854 254452 80860
rect 254308 5636 254360 5642
rect 254308 5578 254360 5584
rect 254216 5568 254268 5574
rect 254216 5510 254268 5516
rect 254124 4820 254176 4826
rect 254124 4762 254176 4768
rect 254688 3670 254716 325926
rect 255056 316034 255084 337622
rect 255148 335646 255176 337708
rect 255286 337634 255314 338028
rect 255378 337890 255406 338028
rect 255470 337890 255498 338028
rect 255366 337884 255418 337890
rect 255366 337826 255418 337832
rect 255458 337884 255510 337890
rect 255458 337826 255510 337832
rect 255562 337634 255590 338028
rect 255654 337895 255682 338028
rect 255640 337886 255696 337895
rect 255640 337821 255696 337830
rect 255746 337736 255774 338028
rect 255838 337890 255866 338028
rect 255826 337884 255878 337890
rect 255826 337826 255878 337832
rect 255240 337606 255314 337634
rect 255424 337606 255590 337634
rect 255700 337708 255774 337736
rect 256022 337736 256050 338028
rect 256114 337890 256142 338028
rect 256206 337958 256234 338028
rect 256194 337952 256246 337958
rect 256194 337894 256246 337900
rect 256102 337884 256154 337890
rect 256102 337826 256154 337832
rect 256146 337784 256202 337793
rect 256022 337708 256096 337736
rect 256146 337719 256202 337728
rect 255136 335640 255188 335646
rect 255136 335582 255188 335588
rect 255136 335436 255188 335442
rect 255136 335378 255188 335384
rect 255148 332042 255176 335378
rect 255136 332036 255188 332042
rect 255136 331978 255188 331984
rect 255240 325990 255268 337606
rect 255318 335472 255374 335481
rect 255318 335407 255374 335416
rect 255332 326126 255360 335407
rect 255424 334422 255452 337606
rect 255596 337544 255648 337550
rect 255596 337486 255648 337492
rect 255504 337476 255556 337482
rect 255504 337418 255556 337424
rect 255412 334416 255464 334422
rect 255412 334358 255464 334364
rect 255412 326596 255464 326602
rect 255412 326538 255464 326544
rect 255320 326120 255372 326126
rect 255320 326062 255372 326068
rect 255228 325984 255280 325990
rect 255228 325926 255280 325932
rect 254872 316006 255084 316034
rect 254676 3664 254728 3670
rect 254676 3606 254728 3612
rect 254676 3528 254728 3534
rect 254676 3470 254728 3476
rect 254688 480 254716 3470
rect 254872 3466 254900 316006
rect 255424 3534 255452 326538
rect 255516 326534 255544 337418
rect 255504 326528 255556 326534
rect 255504 326470 255556 326476
rect 255608 326380 255636 337486
rect 255516 326352 255636 326380
rect 255516 3806 255544 326352
rect 255596 326188 255648 326194
rect 255596 326130 255648 326136
rect 255504 3800 255556 3806
rect 255504 3742 255556 3748
rect 255412 3528 255464 3534
rect 255412 3470 255464 3476
rect 255608 3482 255636 326130
rect 255700 4962 255728 337708
rect 255780 337612 255832 337618
rect 255780 337554 255832 337560
rect 255792 332654 255820 337554
rect 255872 337544 255924 337550
rect 255872 337486 255924 337492
rect 255780 332648 255832 332654
rect 255780 332590 255832 332596
rect 255780 326528 255832 326534
rect 255780 326470 255832 326476
rect 255688 4956 255740 4962
rect 255688 4898 255740 4904
rect 255792 4894 255820 326470
rect 255884 8906 255912 337486
rect 255964 326528 256016 326534
rect 255964 326470 256016 326476
rect 255976 9178 256004 326470
rect 256068 326380 256096 337708
rect 256160 326534 256188 337719
rect 256298 337668 256326 338028
rect 256390 337793 256418 338028
rect 256376 337784 256432 337793
rect 256376 337719 256432 337728
rect 256298 337640 256372 337668
rect 256240 337544 256292 337550
rect 256240 337486 256292 337492
rect 256148 326528 256200 326534
rect 256148 326470 256200 326476
rect 256252 326380 256280 337486
rect 256344 326482 256372 337640
rect 256482 337634 256510 338028
rect 256436 337606 256510 337634
rect 256436 326602 256464 337606
rect 256574 337498 256602 338028
rect 256528 337470 256602 337498
rect 256424 326596 256476 326602
rect 256424 326538 256476 326544
rect 256344 326454 256464 326482
rect 256068 326352 256188 326380
rect 256252 326352 256372 326380
rect 256056 326256 256108 326262
rect 256056 326198 256108 326204
rect 256068 84998 256096 326198
rect 256160 88738 256188 326352
rect 256240 326120 256292 326126
rect 256240 326062 256292 326068
rect 256252 239193 256280 326062
rect 256344 321554 256372 326352
rect 256436 326262 256464 326454
rect 256424 326256 256476 326262
rect 256424 326198 256476 326204
rect 256528 326194 256556 337470
rect 256666 337362 256694 338028
rect 256758 337668 256786 338028
rect 256850 337736 256878 338028
rect 256942 338008 256970 338028
rect 257080 338014 257140 338042
rect 256942 337980 257016 338008
rect 256850 337708 256924 337736
rect 256758 337640 256832 337668
rect 256620 337334 256694 337362
rect 256620 335374 256648 337334
rect 256804 335510 256832 337640
rect 256792 335504 256844 335510
rect 256792 335446 256844 335452
rect 256608 335368 256660 335374
rect 256608 335310 256660 335316
rect 256896 326262 256924 337708
rect 256988 333334 257016 337980
rect 257080 335646 257108 338014
rect 257218 337736 257246 338028
rect 257310 337929 257338 338028
rect 257402 337958 257430 338028
rect 257390 337952 257442 337958
rect 257296 337920 257352 337929
rect 257390 337894 257442 337900
rect 257296 337855 257352 337864
rect 257494 337822 257522 338028
rect 257586 337958 257614 338028
rect 257678 337963 257706 338028
rect 257574 337952 257626 337958
rect 257574 337894 257626 337900
rect 257664 337954 257720 337963
rect 257770 337958 257798 338028
rect 257862 337958 257890 338028
rect 257664 337889 257720 337898
rect 257758 337952 257810 337958
rect 257758 337894 257810 337900
rect 257850 337952 257902 337958
rect 257850 337894 257902 337900
rect 257482 337816 257534 337822
rect 257342 337784 257398 337793
rect 257218 337708 257292 337736
rect 257482 337758 257534 337764
rect 257342 337719 257398 337728
rect 257804 337748 257856 337754
rect 257160 337612 257212 337618
rect 257160 337554 257212 337560
rect 257068 335640 257120 335646
rect 257068 335582 257120 335588
rect 257068 335368 257120 335374
rect 257068 335310 257120 335316
rect 256976 333328 257028 333334
rect 256976 333270 257028 333276
rect 256884 326256 256936 326262
rect 256884 326198 256936 326204
rect 256516 326188 256568 326194
rect 256516 326130 256568 326136
rect 256344 321526 256464 321554
rect 256238 239184 256294 239193
rect 256238 239119 256294 239128
rect 256148 88732 256200 88738
rect 256148 88674 256200 88680
rect 256056 84992 256108 84998
rect 256056 84934 256108 84940
rect 255964 9172 256016 9178
rect 255964 9114 256016 9120
rect 255872 8900 255924 8906
rect 255872 8842 255924 8848
rect 255780 4888 255832 4894
rect 255780 4830 255832 4836
rect 254860 3460 254912 3466
rect 255608 3454 255912 3482
rect 254860 3402 254912 3408
rect 255884 480 255912 3454
rect 256436 3398 256464 321526
rect 256424 3392 256476 3398
rect 256424 3334 256476 3340
rect 257080 480 257108 335310
rect 257172 3466 257200 337554
rect 257264 336122 257292 337708
rect 257252 336116 257304 336122
rect 257252 336058 257304 336064
rect 257252 335912 257304 335918
rect 257252 335854 257304 335860
rect 257264 333266 257292 335854
rect 257252 333260 257304 333266
rect 257252 333202 257304 333208
rect 257356 5370 257384 337719
rect 257954 337736 257982 338028
rect 258046 337890 258074 338028
rect 258034 337884 258086 337890
rect 258034 337826 258086 337832
rect 258138 337770 258166 338028
rect 257804 337690 257856 337696
rect 257908 337708 257982 337736
rect 258092 337742 258166 337770
rect 258276 338014 258336 338042
rect 257620 337680 257672 337686
rect 257434 337648 257490 337657
rect 257620 337622 257672 337628
rect 257434 337583 257490 337592
rect 257448 328454 257476 337583
rect 257448 328426 257568 328454
rect 257436 326528 257488 326534
rect 257436 326470 257488 326476
rect 257344 5364 257396 5370
rect 257344 5306 257396 5312
rect 257448 5166 257476 326470
rect 257540 5234 257568 328426
rect 257632 5302 257660 337622
rect 257816 326534 257844 337690
rect 257804 326528 257856 326534
rect 257804 326470 257856 326476
rect 257908 326380 257936 337708
rect 258092 335782 258120 337742
rect 258080 335776 258132 335782
rect 258080 335718 258132 335724
rect 258172 335708 258224 335714
rect 258172 335650 258224 335656
rect 258080 335504 258132 335510
rect 258080 335446 258132 335452
rect 257988 333328 258040 333334
rect 257988 333270 258040 333276
rect 257724 326352 257936 326380
rect 257620 5296 257672 5302
rect 257620 5238 257672 5244
rect 257528 5228 257580 5234
rect 257528 5170 257580 5176
rect 257436 5160 257488 5166
rect 257436 5102 257488 5108
rect 257724 5098 257752 326352
rect 257804 326256 257856 326262
rect 257804 326198 257856 326204
rect 257712 5092 257764 5098
rect 257712 5034 257764 5040
rect 257816 3534 257844 326198
rect 258000 316034 258028 333270
rect 257908 316006 258028 316034
rect 257908 3602 257936 316006
rect 258092 16574 258120 335446
rect 258184 333402 258212 335650
rect 258276 335510 258304 338014
rect 258414 337736 258442 338028
rect 258368 337708 258442 337736
rect 258506 337736 258534 338028
rect 258598 337890 258626 338028
rect 258586 337884 258638 337890
rect 258586 337826 258638 337832
rect 258690 337736 258718 338028
rect 258506 337708 258580 337736
rect 258368 335714 258396 337708
rect 258356 335708 258408 335714
rect 258356 335650 258408 335656
rect 258264 335504 258316 335510
rect 258264 335446 258316 335452
rect 258448 335436 258500 335442
rect 258448 335378 258500 335384
rect 258356 335368 258408 335374
rect 258356 335310 258408 335316
rect 258172 333396 258224 333402
rect 258172 333338 258224 333344
rect 258092 16546 258304 16574
rect 257896 3596 257948 3602
rect 257896 3538 257948 3544
rect 257804 3528 257856 3534
rect 257804 3470 257856 3476
rect 257160 3460 257212 3466
rect 257160 3402 257212 3408
rect 258276 480 258304 16546
rect 258368 4826 258396 335310
rect 258460 239834 258488 335378
rect 258552 326398 258580 337708
rect 258644 337708 258718 337736
rect 258540 326392 258592 326398
rect 258540 326334 258592 326340
rect 258644 316034 258672 337708
rect 258782 337668 258810 338028
rect 258874 337958 258902 338028
rect 258862 337952 258914 337958
rect 258862 337894 258914 337900
rect 258966 337770 258994 338028
rect 258736 337640 258810 337668
rect 258920 337742 258994 337770
rect 259058 337770 259086 338028
rect 259150 337958 259178 338028
rect 259138 337952 259190 337958
rect 259138 337894 259190 337900
rect 259242 337906 259270 338028
rect 259334 338008 259362 338028
rect 259472 338014 259532 338042
rect 259334 337980 259408 338008
rect 259242 337878 259316 337906
rect 259058 337742 259132 337770
rect 258736 335374 258764 337640
rect 258816 336252 258868 336258
rect 258816 336194 258868 336200
rect 258724 335368 258776 335374
rect 258724 335310 258776 335316
rect 258828 332110 258856 336194
rect 258816 332104 258868 332110
rect 258816 332046 258868 332052
rect 258920 331214 258948 337742
rect 259000 337680 259052 337686
rect 259000 337622 259052 337628
rect 258552 316006 258672 316034
rect 258828 331186 258948 331214
rect 258448 239828 258500 239834
rect 258448 239770 258500 239776
rect 258356 4820 258408 4826
rect 258356 4762 258408 4768
rect 258552 3670 258580 316006
rect 258828 89078 258856 331186
rect 258908 326392 258960 326398
rect 258908 326334 258960 326340
rect 258816 89072 258868 89078
rect 258816 89014 258868 89020
rect 258920 4962 258948 326334
rect 258908 4956 258960 4962
rect 258908 4898 258960 4904
rect 259012 4758 259040 337622
rect 259104 335442 259132 337742
rect 259184 337612 259236 337618
rect 259184 337554 259236 337560
rect 259092 335436 259144 335442
rect 259092 335378 259144 335384
rect 259092 335300 259144 335306
rect 259092 335242 259144 335248
rect 259104 5030 259132 335242
rect 259092 5024 259144 5030
rect 259092 4966 259144 4972
rect 259196 4894 259224 337554
rect 259288 335442 259316 337878
rect 259276 335436 259328 335442
rect 259276 335378 259328 335384
rect 259276 335300 259328 335306
rect 259276 335242 259328 335248
rect 259288 331906 259316 335242
rect 259380 334082 259408 337980
rect 259472 335714 259500 338014
rect 259610 337736 259638 338028
rect 259564 337708 259638 337736
rect 259460 335708 259512 335714
rect 259460 335650 259512 335656
rect 259564 335594 259592 337708
rect 259702 337668 259730 338028
rect 259794 337736 259822 338028
rect 259886 337890 259914 338028
rect 259874 337884 259926 337890
rect 259874 337826 259926 337832
rect 259978 337736 260006 338028
rect 260070 337890 260098 338028
rect 260162 337958 260190 338028
rect 260254 337958 260282 338028
rect 260150 337952 260202 337958
rect 260150 337894 260202 337900
rect 260242 337952 260294 337958
rect 260242 337894 260294 337900
rect 260058 337884 260110 337890
rect 260058 337826 260110 337832
rect 260346 337770 260374 338028
rect 260438 337872 260466 338028
rect 260576 338014 260636 338042
rect 260438 337844 260512 337872
rect 260300 337742 260374 337770
rect 259794 337708 259868 337736
rect 259978 337708 260052 337736
rect 259702 337640 259776 337668
rect 259748 335850 259776 337640
rect 259736 335844 259788 335850
rect 259736 335786 259788 335792
rect 259736 335708 259788 335714
rect 259736 335650 259788 335656
rect 259460 335572 259512 335578
rect 259564 335566 259684 335594
rect 259460 335514 259512 335520
rect 259368 334076 259420 334082
rect 259368 334018 259420 334024
rect 259276 331900 259328 331906
rect 259276 331842 259328 331848
rect 259184 4888 259236 4894
rect 259184 4830 259236 4836
rect 259000 4752 259052 4758
rect 259000 4694 259052 4700
rect 259472 4282 259500 335514
rect 259552 335504 259604 335510
rect 259552 335446 259604 335452
rect 259564 332178 259592 335446
rect 259552 332172 259604 332178
rect 259552 332114 259604 332120
rect 259656 331702 259684 335566
rect 259644 331696 259696 331702
rect 259644 331638 259696 331644
rect 259644 326188 259696 326194
rect 259644 326130 259696 326136
rect 259656 4350 259684 326130
rect 259748 321554 259776 335650
rect 259840 335510 259868 337708
rect 259920 337612 259972 337618
rect 259920 337554 259972 337560
rect 259828 335504 259880 335510
rect 259828 335446 259880 335452
rect 259932 335374 259960 337554
rect 260024 335714 260052 337708
rect 260196 337544 260248 337550
rect 260196 337486 260248 337492
rect 260012 335708 260064 335714
rect 260012 335650 260064 335656
rect 260104 335640 260156 335646
rect 260104 335582 260156 335588
rect 260012 335436 260064 335442
rect 260012 335378 260064 335384
rect 259920 335368 259972 335374
rect 259920 335310 259972 335316
rect 259828 335300 259880 335306
rect 259828 335242 259880 335248
rect 259840 326194 259868 335242
rect 259828 326188 259880 326194
rect 259828 326130 259880 326136
rect 259748 321526 259868 321554
rect 259840 5506 259868 321526
rect 260024 238202 260052 335378
rect 260012 238196 260064 238202
rect 260012 238138 260064 238144
rect 259828 5500 259880 5506
rect 259828 5442 259880 5448
rect 259644 4344 259696 4350
rect 259644 4286 259696 4292
rect 259460 4276 259512 4282
rect 259460 4218 259512 4224
rect 258540 3664 258592 3670
rect 258540 3606 258592 3612
rect 260116 3534 260144 335582
rect 260208 326262 260236 337486
rect 260300 335578 260328 337742
rect 260484 335918 260512 337844
rect 260472 335912 260524 335918
rect 260472 335854 260524 335860
rect 260380 335708 260432 335714
rect 260380 335650 260432 335656
rect 260288 335572 260340 335578
rect 260288 335514 260340 335520
rect 260392 335458 260420 335650
rect 260300 335430 260420 335458
rect 260472 335504 260524 335510
rect 260472 335446 260524 335452
rect 260300 334150 260328 335430
rect 260380 335368 260432 335374
rect 260380 335310 260432 335316
rect 260288 334144 260340 334150
rect 260288 334086 260340 334092
rect 260288 326392 260340 326398
rect 260288 326334 260340 326340
rect 260196 326256 260248 326262
rect 260196 326198 260248 326204
rect 260300 87854 260328 326334
rect 260288 87848 260340 87854
rect 260288 87790 260340 87796
rect 260392 6866 260420 335310
rect 260380 6860 260432 6866
rect 260380 6802 260432 6808
rect 260484 5438 260512 335446
rect 260576 326398 260604 338014
rect 260714 337872 260742 338028
rect 260668 337844 260742 337872
rect 260668 335374 260696 337844
rect 260806 337736 260834 338028
rect 260898 337890 260926 338028
rect 260886 337884 260938 337890
rect 260886 337826 260938 337832
rect 260990 337736 261018 338028
rect 260760 337708 260834 337736
rect 260944 337708 261018 337736
rect 260760 336530 260788 337708
rect 260840 337612 260892 337618
rect 260840 337554 260892 337560
rect 260748 336524 260800 336530
rect 260748 336466 260800 336472
rect 260852 336462 260880 337554
rect 260840 336456 260892 336462
rect 260840 336398 260892 336404
rect 260840 335436 260892 335442
rect 260840 335378 260892 335384
rect 260656 335368 260708 335374
rect 260656 335310 260708 335316
rect 260564 326392 260616 326398
rect 260564 326334 260616 326340
rect 260564 326256 260616 326262
rect 260564 326198 260616 326204
rect 260472 5432 260524 5438
rect 260472 5374 260524 5380
rect 260576 4214 260604 326198
rect 260852 5574 260880 335378
rect 260944 85134 260972 337708
rect 261082 337668 261110 338028
rect 261036 337640 261110 337668
rect 261036 332586 261064 337640
rect 261174 337498 261202 338028
rect 261266 337634 261294 338028
rect 261358 337770 261386 338028
rect 261450 337890 261478 338028
rect 261438 337884 261490 337890
rect 261438 337826 261490 337832
rect 261542 337770 261570 338028
rect 261634 337906 261662 338028
rect 261818 337958 261846 338028
rect 261910 337963 261938 338028
rect 261806 337952 261858 337958
rect 261634 337878 261708 337906
rect 261806 337894 261858 337900
rect 261896 337954 261952 337963
rect 262002 337958 262030 338028
rect 261896 337889 261952 337898
rect 261990 337952 262042 337958
rect 261990 337894 262042 337900
rect 261358 337742 261432 337770
rect 261266 337606 261340 337634
rect 261174 337470 261248 337498
rect 261220 334286 261248 337470
rect 261312 335374 261340 337606
rect 261404 336054 261432 337742
rect 261496 337742 261570 337770
rect 261392 336048 261444 336054
rect 261392 335990 261444 335996
rect 261300 335368 261352 335374
rect 261300 335310 261352 335316
rect 261208 334280 261260 334286
rect 261208 334222 261260 334228
rect 261024 332580 261076 332586
rect 261024 332522 261076 332528
rect 261496 316034 261524 337742
rect 261576 337680 261628 337686
rect 261576 337622 261628 337628
rect 261588 335458 261616 337622
rect 261680 336870 261708 337878
rect 262094 337822 262122 338028
rect 262186 337890 262214 338028
rect 262174 337884 262226 337890
rect 262174 337826 262226 337832
rect 261760 337816 261812 337822
rect 262082 337816 262134 337822
rect 261760 337758 261812 337764
rect 261942 337784 261998 337793
rect 261668 336864 261720 336870
rect 261668 336806 261720 336812
rect 261588 335430 261708 335458
rect 261576 335368 261628 335374
rect 261576 335310 261628 335316
rect 261128 316006 261524 316034
rect 260932 85128 260984 85134
rect 260932 85070 260984 85076
rect 260840 5568 260892 5574
rect 260840 5510 260892 5516
rect 261128 4486 261156 316006
rect 261116 4480 261168 4486
rect 261116 4422 261168 4428
rect 261588 4418 261616 335310
rect 261680 332722 261708 335430
rect 261668 332716 261720 332722
rect 261668 332658 261720 332664
rect 261772 80918 261800 337758
rect 262082 337758 262134 337764
rect 262278 337736 262306 338028
rect 261942 337719 261998 337728
rect 261760 80912 261812 80918
rect 261760 80854 261812 80860
rect 261956 4554 261984 337719
rect 262232 337708 262306 337736
rect 262128 337680 262180 337686
rect 262128 337622 262180 337628
rect 262140 335442 262168 337622
rect 262128 335436 262180 335442
rect 262128 335378 262180 335384
rect 262232 334626 262260 337708
rect 262370 337668 262398 338028
rect 262324 337640 262398 337668
rect 262462 337668 262490 338028
rect 262554 337822 262582 338028
rect 262646 337890 262674 338028
rect 262634 337884 262686 337890
rect 262738 337872 262766 338028
rect 262830 337940 262858 338028
rect 262968 338014 263028 338042
rect 262830 337912 262904 337940
rect 262738 337844 262812 337872
rect 262634 337826 262686 337832
rect 262542 337816 262594 337822
rect 262542 337758 262594 337764
rect 262462 337640 262536 337668
rect 262220 334620 262272 334626
rect 262220 334562 262272 334568
rect 262220 334484 262272 334490
rect 262220 334426 262272 334432
rect 261944 4548 261996 4554
rect 261944 4490 261996 4496
rect 261576 4412 261628 4418
rect 261576 4354 261628 4360
rect 260564 4208 260616 4214
rect 260564 4150 260616 4156
rect 260656 3596 260708 3602
rect 260656 3538 260708 3544
rect 259460 3528 259512 3534
rect 259460 3470 259512 3476
rect 260104 3528 260156 3534
rect 260104 3470 260156 3476
rect 259472 480 259500 3470
rect 260668 480 260696 3538
rect 261760 3528 261812 3534
rect 261760 3470 261812 3476
rect 261772 480 261800 3470
rect 262232 490 262260 334426
rect 262324 5642 262352 337640
rect 262404 335912 262456 335918
rect 262404 335854 262456 335860
rect 262416 331838 262444 335854
rect 262508 335442 262536 337640
rect 262680 335708 262732 335714
rect 262680 335650 262732 335656
rect 262496 335436 262548 335442
rect 262496 335378 262548 335384
rect 262588 335368 262640 335374
rect 262588 335310 262640 335316
rect 262404 331832 262456 331838
rect 262404 331774 262456 331780
rect 262600 5778 262628 335310
rect 262692 11694 262720 335650
rect 262680 11688 262732 11694
rect 262680 11630 262732 11636
rect 262784 10742 262812 337844
rect 262876 335578 262904 337912
rect 262864 335572 262916 335578
rect 262864 335514 262916 335520
rect 262864 335436 262916 335442
rect 262864 335378 262916 335384
rect 262876 331214 262904 335378
rect 262968 335374 262996 338014
rect 263106 337736 263134 338028
rect 263060 337708 263134 337736
rect 262956 335368 263008 335374
rect 262956 335310 263008 335316
rect 262876 331186 262996 331214
rect 262864 323468 262916 323474
rect 262864 323410 262916 323416
rect 262772 10736 262824 10742
rect 262772 10678 262824 10684
rect 262876 10606 262904 323410
rect 262968 10810 262996 331186
rect 262956 10804 263008 10810
rect 262956 10746 263008 10752
rect 263060 10674 263088 337708
rect 263198 337668 263226 338028
rect 263290 337736 263318 338028
rect 263382 337929 263410 338028
rect 263368 337920 263424 337929
rect 263474 337890 263502 338028
rect 263368 337855 263424 337864
rect 263462 337884 263514 337890
rect 263462 337826 263514 337832
rect 263414 337784 263470 337793
rect 263290 337708 263364 337736
rect 263566 337736 263594 338028
rect 263658 337958 263686 338028
rect 263750 337963 263778 338028
rect 263646 337952 263698 337958
rect 263646 337894 263698 337900
rect 263736 337954 263792 337963
rect 263736 337889 263792 337898
rect 263842 337822 263870 338028
rect 263934 338008 263962 338028
rect 263934 337980 264008 338008
rect 263830 337816 263882 337822
rect 263830 337758 263882 337764
rect 263414 337719 263470 337728
rect 263152 337640 263226 337668
rect 263152 335578 263180 337640
rect 263232 335776 263284 335782
rect 263232 335718 263284 335724
rect 263140 335572 263192 335578
rect 263140 335514 263192 335520
rect 263140 335368 263192 335374
rect 263140 335310 263192 335316
rect 263152 323474 263180 335310
rect 263140 323468 263192 323474
rect 263140 323410 263192 323416
rect 263244 316034 263272 335718
rect 263152 316006 263272 316034
rect 263048 10668 263100 10674
rect 263048 10610 263100 10616
rect 262864 10600 262916 10606
rect 262864 10542 262916 10548
rect 262588 5772 262640 5778
rect 262588 5714 262640 5720
rect 263152 5710 263180 316006
rect 263336 5846 263364 337708
rect 263428 335374 263456 337719
rect 263520 337708 263594 337736
rect 263416 335368 263468 335374
rect 263416 335310 263468 335316
rect 263520 328454 263548 337708
rect 263784 337680 263836 337686
rect 263784 337622 263836 337628
rect 263600 336048 263652 336054
rect 263600 335990 263652 335996
rect 263612 332518 263640 335990
rect 263692 335368 263744 335374
rect 263692 335310 263744 335316
rect 263704 332654 263732 335310
rect 263692 332648 263744 332654
rect 263692 332590 263744 332596
rect 263600 332512 263652 332518
rect 263600 332454 263652 332460
rect 263428 328426 263548 328454
rect 263428 5914 263456 328426
rect 263416 5908 263468 5914
rect 263416 5850 263468 5856
rect 263324 5840 263376 5846
rect 263324 5782 263376 5788
rect 263140 5704 263192 5710
rect 263140 5646 263192 5652
rect 262312 5636 262364 5642
rect 262312 5578 262364 5584
rect 263796 4622 263824 337622
rect 263876 336184 263928 336190
rect 263876 336126 263928 336132
rect 263888 326398 263916 336126
rect 263980 333334 264008 337980
rect 264118 337736 264146 338028
rect 264210 337890 264238 338028
rect 264198 337884 264250 337890
rect 264198 337826 264250 337832
rect 264302 337736 264330 338028
rect 264118 337708 264192 337736
rect 264060 337612 264112 337618
rect 264060 337554 264112 337560
rect 263968 333328 264020 333334
rect 263968 333270 264020 333276
rect 263876 326392 263928 326398
rect 263876 326334 263928 326340
rect 264072 80850 264100 337554
rect 264164 335986 264192 337708
rect 264256 337708 264330 337736
rect 264394 337736 264422 338028
rect 264486 337929 264514 338028
rect 264472 337920 264528 337929
rect 264578 337890 264606 338028
rect 264472 337855 264528 337864
rect 264566 337884 264618 337890
rect 264566 337826 264618 337832
rect 264670 337736 264698 338028
rect 264394 337708 264560 337736
rect 264152 335980 264204 335986
rect 264152 335922 264204 335928
rect 264152 335640 264204 335646
rect 264152 335582 264204 335588
rect 264164 334218 264192 335582
rect 264256 335442 264284 337708
rect 264334 337648 264390 337657
rect 264334 337583 264390 337592
rect 264428 337612 264480 337618
rect 264244 335436 264296 335442
rect 264244 335378 264296 335384
rect 264152 334212 264204 334218
rect 264152 334154 264204 334160
rect 264348 331214 264376 337583
rect 264428 337554 264480 337560
rect 264164 331186 264376 331214
rect 264164 84998 264192 331186
rect 264244 326392 264296 326398
rect 264244 326334 264296 326340
rect 264152 84992 264204 84998
rect 264152 84934 264204 84940
rect 264060 80844 264112 80850
rect 264060 80786 264112 80792
rect 264152 5364 264204 5370
rect 264152 5306 264204 5312
rect 263784 4616 263836 4622
rect 263784 4558 263836 4564
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262232 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 5306
rect 264256 3330 264284 326334
rect 264440 6118 264468 337554
rect 264532 335578 264560 337708
rect 264624 337708 264698 337736
rect 264624 336734 264652 337708
rect 264762 337634 264790 338028
rect 264854 337770 264882 338028
rect 264946 337958 264974 338028
rect 264934 337952 264986 337958
rect 264934 337894 264986 337900
rect 265038 337906 265066 338028
rect 265130 338008 265158 338028
rect 265268 338014 265328 338042
rect 265130 337980 265204 338008
rect 265038 337878 265112 337906
rect 264854 337742 264928 337770
rect 264762 337606 264836 337634
rect 264612 336728 264664 336734
rect 264612 336670 264664 336676
rect 264704 335980 264756 335986
rect 264704 335922 264756 335928
rect 264716 335646 264744 335922
rect 264704 335640 264756 335646
rect 264704 335582 264756 335588
rect 264520 335572 264572 335578
rect 264520 335514 264572 335520
rect 264704 335436 264756 335442
rect 264704 335378 264756 335384
rect 264612 335368 264664 335374
rect 264612 335310 264664 335316
rect 264520 333328 264572 333334
rect 264520 333270 264572 333276
rect 264428 6112 264480 6118
rect 264428 6054 264480 6060
rect 264532 5982 264560 333270
rect 264624 6798 264652 335310
rect 264612 6792 264664 6798
rect 264612 6734 264664 6740
rect 264716 6050 264744 335378
rect 264704 6044 264756 6050
rect 264704 5986 264756 5992
rect 264520 5976 264572 5982
rect 264520 5918 264572 5924
rect 264808 4690 264836 337606
rect 264900 335374 264928 337742
rect 264888 335368 264940 335374
rect 264888 335310 264940 335316
rect 264980 335368 265032 335374
rect 264980 335310 265032 335316
rect 264992 80782 265020 335310
rect 265084 332858 265112 337878
rect 265072 332852 265124 332858
rect 265072 332794 265124 332800
rect 265176 327690 265204 337980
rect 265268 336598 265296 338014
rect 265406 337872 265434 338028
rect 265360 337844 265434 337872
rect 265256 336592 265308 336598
rect 265256 336534 265308 336540
rect 265256 333328 265308 333334
rect 265256 333270 265308 333276
rect 265164 327684 265216 327690
rect 265164 327626 265216 327632
rect 265268 321554 265296 333270
rect 265360 332926 265388 337844
rect 265498 337668 265526 338028
rect 265590 337770 265618 338028
rect 265682 337890 265710 338028
rect 265670 337884 265722 337890
rect 265670 337826 265722 337832
rect 265774 337770 265802 338028
rect 265866 337890 265894 338028
rect 265854 337884 265906 337890
rect 265854 337826 265906 337832
rect 265958 337770 265986 338028
rect 265590 337742 265664 337770
rect 265774 337742 265848 337770
rect 265498 337640 265572 337668
rect 265348 332920 265400 332926
rect 265348 332862 265400 332868
rect 265544 328454 265572 337640
rect 265636 335986 265664 337742
rect 265716 337680 265768 337686
rect 265716 337622 265768 337628
rect 265624 335980 265676 335986
rect 265624 335922 265676 335928
rect 265728 332994 265756 337622
rect 265716 332988 265768 332994
rect 265716 332930 265768 332936
rect 265820 331214 265848 337742
rect 265912 337742 265986 337770
rect 266050 337770 266078 338028
rect 266142 337872 266170 338028
rect 266234 338008 266262 338028
rect 266372 338014 266432 338042
rect 266234 337980 266308 338008
rect 266142 337844 266216 337872
rect 266050 337742 266124 337770
rect 265912 335374 265940 337742
rect 265992 337680 266044 337686
rect 265992 337622 266044 337628
rect 266004 336054 266032 337622
rect 265992 336048 266044 336054
rect 265992 335990 266044 335996
rect 265900 335368 265952 335374
rect 265900 335310 265952 335316
rect 265820 331186 266032 331214
rect 265544 328426 265756 328454
rect 265532 327684 265584 327690
rect 265532 327626 265584 327632
rect 265268 321526 265388 321554
rect 265360 84930 265388 321526
rect 265348 84924 265400 84930
rect 265348 84866 265400 84872
rect 264980 80776 265032 80782
rect 264980 80718 265032 80724
rect 265544 6730 265572 327626
rect 265532 6724 265584 6730
rect 265532 6666 265584 6672
rect 265728 6662 265756 328426
rect 265716 6656 265768 6662
rect 265716 6598 265768 6604
rect 266004 6594 266032 331186
rect 265992 6588 266044 6594
rect 265992 6530 266044 6536
rect 266096 6526 266124 337742
rect 266188 336734 266216 337844
rect 266176 336728 266228 336734
rect 266176 336670 266228 336676
rect 266280 333334 266308 337980
rect 266372 335442 266400 338014
rect 266510 337872 266538 338028
rect 266464 337844 266538 337872
rect 266464 336462 266492 337844
rect 266602 337736 266630 338028
rect 266556 337708 266630 337736
rect 266452 336456 266504 336462
rect 266452 336398 266504 336404
rect 266556 336326 266584 337708
rect 266694 337634 266722 338028
rect 266786 337770 266814 338028
rect 266878 337890 266906 338028
rect 266970 337890 266998 338028
rect 266866 337884 266918 337890
rect 266866 337826 266918 337832
rect 266958 337884 267010 337890
rect 266958 337826 267010 337832
rect 267062 337770 267090 338028
rect 267154 337890 267182 338028
rect 267246 337958 267274 338028
rect 267338 337958 267366 338028
rect 267234 337952 267286 337958
rect 267234 337894 267286 337900
rect 267326 337952 267378 337958
rect 267326 337894 267378 337900
rect 267430 337906 267458 338028
rect 267568 338014 267628 338042
rect 267430 337890 267504 337906
rect 267142 337884 267194 337890
rect 267430 337884 267516 337890
rect 267430 337878 267464 337884
rect 267142 337826 267194 337832
rect 267464 337826 267516 337832
rect 266786 337742 266952 337770
rect 267062 337742 267228 337770
rect 266648 337606 266722 337634
rect 266820 337680 266872 337686
rect 266820 337622 266872 337628
rect 266452 336320 266504 336326
rect 266452 336262 266504 336268
rect 266544 336320 266596 336326
rect 266544 336262 266596 336268
rect 266360 335436 266412 335442
rect 266360 335378 266412 335384
rect 266268 333328 266320 333334
rect 266268 333270 266320 333276
rect 266464 331770 266492 336262
rect 266544 335844 266596 335850
rect 266544 335786 266596 335792
rect 266452 331764 266504 331770
rect 266452 331706 266504 331712
rect 266084 6520 266136 6526
rect 266084 6462 266136 6468
rect 264796 4684 264848 4690
rect 264796 4626 264848 4632
rect 265348 3460 265400 3466
rect 265348 3402 265400 3408
rect 264244 3324 264296 3330
rect 264244 3266 264296 3272
rect 265360 480 265388 3402
rect 266556 480 266584 335786
rect 266648 335782 266676 337606
rect 266728 336320 266780 336326
rect 266728 336262 266780 336268
rect 266636 335776 266688 335782
rect 266636 335718 266688 335724
rect 266636 335368 266688 335374
rect 266636 335310 266688 335316
rect 266648 6390 266676 335310
rect 266740 6458 266768 336262
rect 266832 335374 266860 337622
rect 266924 336394 266952 337742
rect 267004 337680 267056 337686
rect 267004 337622 267056 337628
rect 266912 336388 266964 336394
rect 266912 336330 266964 336336
rect 266912 335504 266964 335510
rect 266912 335446 266964 335452
rect 266820 335368 266872 335374
rect 266820 335310 266872 335316
rect 266924 321554 266952 335446
rect 267016 329118 267044 337622
rect 267096 335776 267148 335782
rect 267096 335718 267148 335724
rect 267108 335458 267136 335718
rect 267200 335578 267228 337742
rect 267464 337748 267516 337754
rect 267464 337690 267516 337696
rect 267188 335572 267240 335578
rect 267188 335514 267240 335520
rect 267108 335430 267228 335458
rect 267096 335368 267148 335374
rect 267096 335310 267148 335316
rect 267004 329112 267056 329118
rect 267004 329054 267056 329060
rect 266924 321526 267044 321554
rect 267016 85066 267044 321526
rect 267004 85060 267056 85066
rect 267004 85002 267056 85008
rect 267108 80714 267136 335310
rect 267096 80708 267148 80714
rect 267096 80650 267148 80656
rect 267200 10470 267228 335430
rect 267372 335300 267424 335306
rect 267372 335242 267424 335248
rect 267280 329112 267332 329118
rect 267280 329054 267332 329060
rect 267188 10464 267240 10470
rect 267188 10406 267240 10412
rect 267292 10402 267320 329054
rect 267384 10538 267412 335242
rect 267372 10532 267424 10538
rect 267372 10474 267424 10480
rect 267280 10396 267332 10402
rect 267280 10338 267332 10344
rect 267476 10334 267504 337690
rect 267568 335374 267596 338014
rect 267706 337872 267734 338028
rect 267660 337844 267734 337872
rect 267660 335646 267688 337844
rect 267798 337736 267826 338028
rect 267890 337890 267918 338028
rect 267878 337884 267930 337890
rect 267878 337826 267930 337832
rect 267798 337708 267872 337736
rect 267648 335640 267700 335646
rect 267648 335582 267700 335588
rect 267556 335368 267608 335374
rect 267556 335310 267608 335316
rect 267844 334558 267872 337708
rect 267982 337600 268010 338028
rect 268074 337668 268102 338028
rect 268166 337770 268194 338028
rect 268258 337958 268286 338028
rect 268246 337952 268298 337958
rect 268246 337894 268298 337900
rect 268350 337895 268378 338028
rect 268336 337886 268392 337895
rect 268336 337821 268392 337830
rect 268166 337754 268332 337770
rect 268166 337748 268344 337754
rect 268166 337742 268292 337748
rect 268442 337736 268470 338028
rect 268534 337872 268562 338028
rect 268626 338008 268654 338028
rect 268626 337980 268700 338008
rect 268534 337844 268608 337872
rect 268292 337690 268344 337696
rect 268396 337708 268470 337736
rect 268074 337640 268148 337668
rect 267982 337572 268056 337600
rect 268028 335850 268056 337572
rect 268016 335844 268068 335850
rect 268016 335786 268068 335792
rect 267924 335368 267976 335374
rect 267924 335310 267976 335316
rect 267832 334552 267884 334558
rect 267832 334494 267884 334500
rect 267740 333328 267792 333334
rect 267740 333270 267792 333276
rect 267464 10328 267516 10334
rect 267464 10270 267516 10276
rect 266728 6452 266780 6458
rect 266728 6394 266780 6400
rect 266636 6384 266688 6390
rect 266636 6326 266688 6332
rect 267752 6322 267780 333270
rect 267740 6316 267792 6322
rect 267740 6258 267792 6264
rect 267936 6254 267964 335310
rect 268120 333130 268148 337640
rect 268292 337612 268344 337618
rect 268292 337554 268344 337560
rect 268200 337408 268252 337414
rect 268200 337350 268252 337356
rect 268212 334694 268240 337350
rect 268200 334688 268252 334694
rect 268200 334630 268252 334636
rect 268108 333124 268160 333130
rect 268108 333066 268160 333072
rect 268304 321554 268332 337554
rect 268396 335374 268424 337708
rect 268474 337648 268530 337657
rect 268474 337583 268530 337592
rect 268488 335730 268516 337583
rect 268580 336598 268608 337844
rect 268568 336592 268620 336598
rect 268568 336534 268620 336540
rect 268488 335702 268608 335730
rect 268580 335578 268608 335702
rect 268476 335572 268528 335578
rect 268476 335514 268528 335520
rect 268568 335572 268620 335578
rect 268568 335514 268620 335520
rect 268384 335368 268436 335374
rect 268384 335310 268436 335316
rect 268382 333296 268438 333305
rect 268382 333231 268438 333240
rect 268396 321706 268424 333231
rect 268384 321700 268436 321706
rect 268384 321642 268436 321648
rect 268212 321526 268332 321554
rect 267924 6248 267976 6254
rect 267924 6190 267976 6196
rect 267740 5296 267792 5302
rect 267740 5238 267792 5244
rect 267752 480 267780 5238
rect 268212 3398 268240 321526
rect 268488 316034 268516 335514
rect 268568 335436 268620 335442
rect 268568 335378 268620 335384
rect 268396 316006 268516 316034
rect 268396 8430 268424 316006
rect 268580 177614 268608 335378
rect 268672 333810 268700 337980
rect 268810 337736 268838 338028
rect 268902 337890 268930 338028
rect 268890 337884 268942 337890
rect 268890 337826 268942 337832
rect 268994 337736 269022 338028
rect 268810 337708 268884 337736
rect 268752 335368 268804 335374
rect 268752 335310 268804 335316
rect 268660 333804 268712 333810
rect 268660 333746 268712 333752
rect 268660 333328 268712 333334
rect 268660 333270 268712 333276
rect 268568 177608 268620 177614
rect 268568 177550 268620 177556
rect 268672 87786 268700 333270
rect 268660 87780 268712 87786
rect 268660 87722 268712 87728
rect 268764 8566 268792 335310
rect 268752 8560 268804 8566
rect 268752 8502 268804 8508
rect 268384 8424 268436 8430
rect 268384 8366 268436 8372
rect 268856 6186 268884 337708
rect 268948 337708 269022 337736
rect 268948 335374 268976 337708
rect 269086 337634 269114 338028
rect 269040 337606 269114 337634
rect 269178 337634 269206 338028
rect 269270 337890 269298 338028
rect 269258 337884 269310 337890
rect 269258 337826 269310 337832
rect 269362 337770 269390 338028
rect 269454 337890 269482 338028
rect 269442 337884 269494 337890
rect 269442 337826 269494 337832
rect 269546 337770 269574 338028
rect 269638 337872 269666 338028
rect 269868 338014 269928 338042
rect 269764 337884 269816 337890
rect 269638 337844 269712 337872
rect 269316 337742 269390 337770
rect 269500 337742 269574 337770
rect 269178 337606 269252 337634
rect 269040 335442 269068 337606
rect 269224 336666 269252 337606
rect 269212 336660 269264 336666
rect 269212 336602 269264 336608
rect 269120 335776 269172 335782
rect 269118 335744 269120 335753
rect 269172 335744 269174 335753
rect 269118 335679 269174 335688
rect 269120 335572 269172 335578
rect 269120 335514 269172 335520
rect 269028 335436 269080 335442
rect 269028 335378 269080 335384
rect 268936 335368 268988 335374
rect 268936 335310 268988 335316
rect 268936 335164 268988 335170
rect 268936 335106 268988 335112
rect 268948 333878 268976 335106
rect 268936 333872 268988 333878
rect 268936 333814 268988 333820
rect 269132 333742 269160 335514
rect 269212 335504 269264 335510
rect 269212 335446 269264 335452
rect 269120 333736 269172 333742
rect 269120 333678 269172 333684
rect 269224 333674 269252 335446
rect 269316 335442 269344 337742
rect 269396 337680 269448 337686
rect 269396 337622 269448 337628
rect 269408 335458 269436 337622
rect 269500 335578 269528 337742
rect 269580 337612 269632 337618
rect 269580 337554 269632 337560
rect 269488 335572 269540 335578
rect 269488 335514 269540 335520
rect 269304 335436 269356 335442
rect 269408 335430 269528 335458
rect 269304 335378 269356 335384
rect 269396 335368 269448 335374
rect 269396 335310 269448 335316
rect 269212 333668 269264 333674
rect 269212 333610 269264 333616
rect 269118 333568 269174 333577
rect 269118 333503 269174 333512
rect 269132 326126 269160 333503
rect 269120 326120 269172 326126
rect 269120 326062 269172 326068
rect 269408 6497 269436 335310
rect 269500 335102 269528 335430
rect 269488 335096 269540 335102
rect 269488 335038 269540 335044
rect 269394 6488 269450 6497
rect 269394 6423 269450 6432
rect 268844 6180 268896 6186
rect 268844 6122 268896 6128
rect 268844 5228 268896 5234
rect 268844 5170 268896 5176
rect 268200 3392 268252 3398
rect 268200 3334 268252 3340
rect 268856 480 268884 5170
rect 269592 3874 269620 337554
rect 269684 335374 269712 337844
rect 269764 337826 269816 337832
rect 269672 335368 269724 335374
rect 269672 335310 269724 335316
rect 269776 328454 269804 337826
rect 269868 335578 269896 338014
rect 270006 337958 270034 338028
rect 269994 337952 270046 337958
rect 269994 337894 270046 337900
rect 270098 337736 270126 338028
rect 270190 337958 270218 338028
rect 270178 337952 270230 337958
rect 270178 337894 270230 337900
rect 270282 337890 270310 338028
rect 270270 337884 270322 337890
rect 270270 337826 270322 337832
rect 270374 337736 270402 338028
rect 270098 337708 270172 337736
rect 269856 335572 269908 335578
rect 269856 335514 269908 335520
rect 269856 335436 269908 335442
rect 269856 335378 269908 335384
rect 270040 335436 270092 335442
rect 270040 335378 270092 335384
rect 269684 328426 269804 328454
rect 269684 177546 269712 328426
rect 269764 326460 269816 326466
rect 269764 326402 269816 326408
rect 269776 326210 269804 326402
rect 269868 326346 269896 335378
rect 269948 335232 270000 335238
rect 269948 335174 270000 335180
rect 269960 326466 269988 335174
rect 269948 326460 270000 326466
rect 269948 326402 270000 326408
rect 269868 326318 269988 326346
rect 269776 326182 269896 326210
rect 269764 326120 269816 326126
rect 269764 326062 269816 326068
rect 269672 177540 269724 177546
rect 269672 177482 269724 177488
rect 269580 3868 269632 3874
rect 269580 3810 269632 3816
rect 269776 3126 269804 326062
rect 269868 8498 269896 326182
rect 269960 87718 269988 326318
rect 269948 87712 270000 87718
rect 269948 87654 270000 87660
rect 270052 8702 270080 335378
rect 270040 8696 270092 8702
rect 270040 8638 270092 8644
rect 270144 8634 270172 337708
rect 270328 337708 270402 337736
rect 270328 336054 270356 337708
rect 270466 337634 270494 338028
rect 270558 337890 270586 338028
rect 270650 337958 270678 338028
rect 270742 337958 270770 338028
rect 270834 337963 270862 338028
rect 270638 337952 270690 337958
rect 270638 337894 270690 337900
rect 270730 337952 270782 337958
rect 270730 337894 270782 337900
rect 270820 337954 270876 337963
rect 270546 337884 270598 337890
rect 270820 337889 270876 337898
rect 270926 337906 270954 338028
rect 271064 338014 271124 338042
rect 270926 337878 271000 337906
rect 270546 337826 270598 337832
rect 270420 337606 270494 337634
rect 270316 336048 270368 336054
rect 270316 335990 270368 335996
rect 270420 335442 270448 337606
rect 270776 337544 270828 337550
rect 270776 337486 270828 337492
rect 270500 335912 270552 335918
rect 270500 335854 270552 335860
rect 270408 335436 270460 335442
rect 270408 335378 270460 335384
rect 270224 335164 270276 335170
rect 270224 335106 270276 335112
rect 270132 8628 270184 8634
rect 270132 8570 270184 8576
rect 269856 8492 269908 8498
rect 269856 8434 269908 8440
rect 270236 6361 270264 335106
rect 270512 334490 270540 335854
rect 270500 334484 270552 334490
rect 270500 334426 270552 334432
rect 270500 326528 270552 326534
rect 270500 326470 270552 326476
rect 270512 7002 270540 326470
rect 270788 89010 270816 337486
rect 270972 337210 271000 337878
rect 270960 337204 271012 337210
rect 270960 337146 271012 337152
rect 270868 336524 270920 336530
rect 270868 336466 270920 336472
rect 270880 336002 270908 336466
rect 270880 335974 271000 336002
rect 270868 333396 270920 333402
rect 270868 333338 270920 333344
rect 270880 326126 270908 333338
rect 270972 326602 271000 335974
rect 271064 335714 271092 338014
rect 271202 337804 271230 338028
rect 271294 337958 271322 338028
rect 271386 337958 271414 338028
rect 271282 337952 271334 337958
rect 271282 337894 271334 337900
rect 271374 337952 271426 337958
rect 271374 337894 271426 337900
rect 271478 337804 271506 338028
rect 271202 337776 271322 337804
rect 271294 337668 271322 337776
rect 271156 337640 271322 337668
rect 271432 337776 271506 337804
rect 271052 335708 271104 335714
rect 271052 335650 271104 335656
rect 271052 335368 271104 335374
rect 271052 335310 271104 335316
rect 270960 326596 271012 326602
rect 270960 326538 271012 326544
rect 270960 326460 271012 326466
rect 270960 326402 271012 326408
rect 270868 326120 270920 326126
rect 270868 326062 270920 326068
rect 270776 89004 270828 89010
rect 270776 88946 270828 88952
rect 270500 6996 270552 7002
rect 270500 6938 270552 6944
rect 270222 6352 270278 6361
rect 270222 6287 270278 6296
rect 270972 6225 271000 326402
rect 271064 177478 271092 335310
rect 271156 326466 271184 337640
rect 271328 335436 271380 335442
rect 271328 335378 271380 335384
rect 271340 331214 271368 335378
rect 271248 331186 271368 331214
rect 271144 326460 271196 326466
rect 271144 326402 271196 326408
rect 271248 326346 271276 331186
rect 271328 326596 271380 326602
rect 271328 326538 271380 326544
rect 271156 326318 271276 326346
rect 271052 177472 271104 177478
rect 271052 177414 271104 177420
rect 270958 6216 271014 6225
rect 270958 6151 271014 6160
rect 271156 3466 271184 326318
rect 271340 326210 271368 326538
rect 271432 326534 271460 337776
rect 271570 337736 271598 338028
rect 271662 337822 271690 338028
rect 271650 337816 271702 337822
rect 271650 337758 271702 337764
rect 271524 337708 271598 337736
rect 271524 336938 271552 337708
rect 271754 337634 271782 338028
rect 271708 337606 271782 337634
rect 271512 336932 271564 336938
rect 271512 336874 271564 336880
rect 271708 335374 271736 337606
rect 271846 337498 271874 338028
rect 271938 337634 271966 338028
rect 272030 337770 272058 338028
rect 272122 337890 272150 338028
rect 272306 337890 272334 338028
rect 272110 337884 272162 337890
rect 272110 337826 272162 337832
rect 272294 337884 272346 337890
rect 272294 337826 272346 337832
rect 272030 337742 272104 337770
rect 272076 337634 272104 337742
rect 272398 337736 272426 338028
rect 272490 337890 272518 338028
rect 272478 337884 272530 337890
rect 272478 337826 272530 337832
rect 272582 337822 272610 338028
rect 272674 337958 272702 338028
rect 272662 337952 272714 337958
rect 272766 337929 272794 338028
rect 272662 337894 272714 337900
rect 272752 337920 272808 337929
rect 272752 337855 272808 337864
rect 272858 337822 272886 338028
rect 272570 337816 272622 337822
rect 272570 337758 272622 337764
rect 272846 337816 272898 337822
rect 272846 337758 272898 337764
rect 272950 337770 272978 338028
rect 273042 337890 273070 338028
rect 273030 337884 273082 337890
rect 273030 337826 273082 337832
rect 272950 337742 273024 337770
rect 272352 337708 272426 337736
rect 271938 337606 272012 337634
rect 272076 337606 272196 337634
rect 271800 337470 271874 337498
rect 271800 336025 271828 337470
rect 271880 337408 271932 337414
rect 271880 337350 271932 337356
rect 271786 336016 271842 336025
rect 271786 335951 271842 335960
rect 271696 335368 271748 335374
rect 271696 335310 271748 335316
rect 271604 335300 271656 335306
rect 271604 335242 271656 335248
rect 271616 333554 271644 335242
rect 271892 334762 271920 337350
rect 271984 335866 272012 337606
rect 271984 335838 272104 335866
rect 271972 335368 272024 335374
rect 271972 335310 272024 335316
rect 271880 334756 271932 334762
rect 271880 334698 271932 334704
rect 271616 333526 271736 333554
rect 271604 333396 271656 333402
rect 271604 333338 271656 333344
rect 271512 333192 271564 333198
rect 271512 333134 271564 333140
rect 271420 326528 271472 326534
rect 271420 326470 271472 326476
rect 271420 326392 271472 326398
rect 271420 326334 271472 326340
rect 271248 326182 271368 326210
rect 271248 11762 271276 326182
rect 271328 326120 271380 326126
rect 271328 326062 271380 326068
rect 271236 11756 271288 11762
rect 271236 11698 271288 11704
rect 271236 5160 271288 5166
rect 271236 5102 271288 5108
rect 271144 3460 271196 3466
rect 271144 3402 271196 3408
rect 270040 3324 270092 3330
rect 270040 3266 270092 3272
rect 269764 3120 269816 3126
rect 269764 3062 269816 3068
rect 270052 480 270080 3266
rect 271248 480 271276 5102
rect 271340 3058 271368 326062
rect 271432 3194 271460 326334
rect 271524 16574 271552 333134
rect 271616 326398 271644 333338
rect 271708 333198 271736 333526
rect 271696 333192 271748 333198
rect 271696 333134 271748 333140
rect 271604 326392 271656 326398
rect 271604 326334 271656 326340
rect 271984 240038 272012 335310
rect 272076 334898 272104 335838
rect 272064 334892 272116 334898
rect 272064 334834 272116 334840
rect 272064 334756 272116 334762
rect 272064 334698 272116 334704
rect 271972 240032 272024 240038
rect 271972 239974 272024 239980
rect 272076 84862 272104 334698
rect 272168 330750 272196 337606
rect 272248 336116 272300 336122
rect 272248 336058 272300 336064
rect 272260 335617 272288 336058
rect 272246 335608 272302 335617
rect 272246 335543 272302 335552
rect 272352 335374 272380 337708
rect 272892 337680 272944 337686
rect 272892 337622 272944 337628
rect 272432 337612 272484 337618
rect 272432 337554 272484 337560
rect 272444 335889 272472 337554
rect 272524 337544 272576 337550
rect 272524 337486 272576 337492
rect 272800 337544 272852 337550
rect 272800 337486 272852 337492
rect 272430 335880 272486 335889
rect 272430 335815 272486 335824
rect 272340 335368 272392 335374
rect 272340 335310 272392 335316
rect 272156 330744 272208 330750
rect 272156 330686 272208 330692
rect 272064 84856 272116 84862
rect 272064 84798 272116 84804
rect 271524 16546 271644 16574
rect 271512 11756 271564 11762
rect 271512 11698 271564 11704
rect 271524 3330 271552 11698
rect 271616 8362 271644 16546
rect 272536 8838 272564 337486
rect 272616 335368 272668 335374
rect 272616 335310 272668 335316
rect 272628 8906 272656 335310
rect 272812 235346 272840 337486
rect 272904 333441 272932 337622
rect 272890 333432 272946 333441
rect 272890 333367 272946 333376
rect 272800 235340 272852 235346
rect 272800 235282 272852 235288
rect 272996 82142 273024 337742
rect 273134 337736 273162 338028
rect 273088 337708 273162 337736
rect 273226 337736 273254 338028
rect 273364 338014 273424 338042
rect 273226 337708 273300 337736
rect 273088 335374 273116 337708
rect 273272 337482 273300 337708
rect 273260 337476 273312 337482
rect 273260 337418 273312 337424
rect 273364 337362 273392 338014
rect 273502 337872 273530 338028
rect 273272 337334 273392 337362
rect 273456 337844 273530 337872
rect 273076 335368 273128 335374
rect 273076 335310 273128 335316
rect 273272 331430 273300 337334
rect 273352 337272 273404 337278
rect 273352 337214 273404 337220
rect 273364 333713 273392 337214
rect 273456 333849 273484 337844
rect 273594 337736 273622 338028
rect 273548 337708 273622 337736
rect 273686 337736 273714 338028
rect 273778 337890 273806 338028
rect 273766 337884 273818 337890
rect 273766 337826 273818 337832
rect 273870 337736 273898 338028
rect 273686 337708 273760 337736
rect 273548 335374 273576 337708
rect 273732 337142 273760 337708
rect 273824 337708 273898 337736
rect 273720 337136 273772 337142
rect 273720 337078 273772 337084
rect 273720 335640 273772 335646
rect 273720 335582 273772 335588
rect 273628 335572 273680 335578
rect 273628 335514 273680 335520
rect 273536 335368 273588 335374
rect 273536 335310 273588 335316
rect 273442 333840 273498 333849
rect 273442 333775 273498 333784
rect 273350 333704 273406 333713
rect 273350 333639 273406 333648
rect 273260 331424 273312 331430
rect 273260 331366 273312 331372
rect 272984 82136 273036 82142
rect 272984 82078 273036 82084
rect 272616 8900 272668 8906
rect 272616 8842 272668 8848
rect 272524 8832 272576 8838
rect 272524 8774 272576 8780
rect 271604 8356 271656 8362
rect 271604 8298 271656 8304
rect 273640 7138 273668 335514
rect 273732 335481 273760 335582
rect 273718 335472 273774 335481
rect 273718 335407 273774 335416
rect 273824 330682 273852 337708
rect 273962 337668 273990 338028
rect 274054 337822 274082 338028
rect 274042 337816 274094 337822
rect 274042 337758 274094 337764
rect 274146 337668 274174 338028
rect 274238 337890 274266 338028
rect 274330 337940 274358 338028
rect 274422 338008 274450 338028
rect 274560 338014 274620 338042
rect 274422 337980 274496 338008
rect 274330 337912 274404 337940
rect 274226 337884 274278 337890
rect 274226 337826 274278 337832
rect 274376 337770 274404 337912
rect 274468 337822 274496 337980
rect 274284 337742 274404 337770
rect 274456 337816 274508 337822
rect 274456 337758 274508 337764
rect 273962 337640 274036 337668
rect 274146 337640 274220 337668
rect 274008 335481 274036 337640
rect 274088 337544 274140 337550
rect 274088 337486 274140 337492
rect 273994 335472 274050 335481
rect 273994 335407 274050 335416
rect 273996 335368 274048 335374
rect 273996 335310 274048 335316
rect 273812 330676 273864 330682
rect 273812 330618 273864 330624
rect 273720 330336 273772 330342
rect 273720 330278 273772 330284
rect 273628 7132 273680 7138
rect 273628 7074 273680 7080
rect 273732 7070 273760 330278
rect 273904 330268 273956 330274
rect 273904 330210 273956 330216
rect 273916 8770 273944 330210
rect 274008 239630 274036 335310
rect 274100 330562 274128 337486
rect 274192 335578 274220 337640
rect 274180 335572 274232 335578
rect 274180 335514 274232 335520
rect 274284 335374 274312 337742
rect 274456 337680 274508 337686
rect 274456 337622 274508 337628
rect 274364 337612 274416 337618
rect 274364 337554 274416 337560
rect 274272 335368 274324 335374
rect 274272 335310 274324 335316
rect 274180 335300 274232 335306
rect 274180 335242 274232 335248
rect 274192 331214 274220 335242
rect 274270 335200 274326 335209
rect 274270 335135 274326 335144
rect 274284 331566 274312 335135
rect 274272 331560 274324 331566
rect 274272 331502 274324 331508
rect 274192 331186 274312 331214
rect 274100 330534 274220 330562
rect 274088 330200 274140 330206
rect 274088 330142 274140 330148
rect 273996 239624 274048 239630
rect 273996 239566 274048 239572
rect 274100 162178 274128 330142
rect 274192 239698 274220 330534
rect 274180 239692 274232 239698
rect 274180 239634 274232 239640
rect 274088 162172 274140 162178
rect 274088 162114 274140 162120
rect 274284 87650 274312 331186
rect 274272 87644 274324 87650
rect 274272 87586 274324 87592
rect 273904 8764 273956 8770
rect 273904 8706 273956 8712
rect 274376 7206 274404 337554
rect 274468 336569 274496 337622
rect 274454 336560 274510 336569
rect 274454 336495 274510 336504
rect 274560 334354 274588 338014
rect 274698 337872 274726 338028
rect 274652 337844 274726 337872
rect 274548 334348 274600 334354
rect 274548 334290 274600 334296
rect 274652 333577 274680 337844
rect 274790 337736 274818 338028
rect 274882 337890 274910 338028
rect 274870 337884 274922 337890
rect 274870 337826 274922 337832
rect 274790 337708 274864 337736
rect 274732 337612 274784 337618
rect 274732 337554 274784 337560
rect 274744 335458 274772 337554
rect 274836 335986 274864 337708
rect 274974 337668 275002 338028
rect 275066 337736 275094 338028
rect 275158 337890 275186 338028
rect 275250 337890 275278 338028
rect 275146 337884 275198 337890
rect 275146 337826 275198 337832
rect 275238 337884 275290 337890
rect 275238 337826 275290 337832
rect 275342 337770 275370 338028
rect 275204 337742 275370 337770
rect 275066 337708 275140 337736
rect 274974 337640 275048 337668
rect 274916 336116 274968 336122
rect 274916 336058 274968 336064
rect 274824 335980 274876 335986
rect 274824 335922 274876 335928
rect 274744 335430 274864 335458
rect 274732 335300 274784 335306
rect 274732 335242 274784 335248
rect 274638 333568 274694 333577
rect 274638 333503 274694 333512
rect 274744 239494 274772 335242
rect 274836 331362 274864 335430
rect 274824 331356 274876 331362
rect 274824 331298 274876 331304
rect 274928 325694 274956 336058
rect 275020 335578 275048 337640
rect 275112 335918 275140 337708
rect 275100 335912 275152 335918
rect 275100 335854 275152 335860
rect 275008 335572 275060 335578
rect 275008 335514 275060 335520
rect 275204 328454 275232 337742
rect 275434 337668 275462 338028
rect 275526 338008 275554 338028
rect 275664 338014 275724 338042
rect 275526 337980 275600 338008
rect 275282 337648 275338 337657
rect 275282 337583 275338 337592
rect 275388 337640 275462 337668
rect 275296 332246 275324 337583
rect 275284 332240 275336 332246
rect 275284 332182 275336 332188
rect 275388 331498 275416 337640
rect 275468 337544 275520 337550
rect 275468 337486 275520 337492
rect 275480 336433 275508 337486
rect 275466 336424 275522 336433
rect 275466 336359 275522 336368
rect 275572 335753 275600 337980
rect 275558 335744 275614 335753
rect 275558 335679 275614 335688
rect 275560 335572 275612 335578
rect 275560 335514 275612 335520
rect 275468 335368 275520 335374
rect 275468 335310 275520 335316
rect 275376 331492 275428 331498
rect 275376 331434 275428 331440
rect 275376 330676 275428 330682
rect 275376 330618 275428 330624
rect 275204 328426 275324 328454
rect 274928 325666 275140 325694
rect 274732 239488 274784 239494
rect 274732 239430 274784 239436
rect 274824 11688 274876 11694
rect 274824 11630 274876 11636
rect 274364 7200 274416 7206
rect 274364 7142 274416 7148
rect 273720 7064 273772 7070
rect 273720 7006 273772 7012
rect 272432 5092 272484 5098
rect 272432 5034 272484 5040
rect 271512 3324 271564 3330
rect 271512 3266 271564 3272
rect 271420 3188 271472 3194
rect 271420 3130 271472 3136
rect 271328 3052 271380 3058
rect 271328 2994 271380 3000
rect 272444 480 272472 5034
rect 273628 3188 273680 3194
rect 273628 3130 273680 3136
rect 273640 480 273668 3130
rect 274836 480 274864 11630
rect 275112 7410 275140 325666
rect 275296 316034 275324 328426
rect 275204 316006 275324 316034
rect 275100 7404 275152 7410
rect 275100 7346 275152 7352
rect 275204 7342 275232 316006
rect 275388 239426 275416 330618
rect 275376 239420 275428 239426
rect 275376 239362 275428 239368
rect 275480 239329 275508 335310
rect 275572 239562 275600 335514
rect 275664 330682 275692 338014
rect 275802 337872 275830 338028
rect 275756 337844 275830 337872
rect 275756 336122 275784 337844
rect 275894 337736 275922 338028
rect 275848 337708 275922 337736
rect 275848 336122 275876 337708
rect 275986 337668 276014 338028
rect 275940 337640 276014 337668
rect 275744 336116 275796 336122
rect 275744 336058 275796 336064
rect 275836 336116 275888 336122
rect 275836 336058 275888 336064
rect 275836 335980 275888 335986
rect 275836 335922 275888 335928
rect 275744 335912 275796 335918
rect 275744 335854 275796 335860
rect 275652 330676 275704 330682
rect 275652 330618 275704 330624
rect 275652 330540 275704 330546
rect 275652 330482 275704 330488
rect 275560 239556 275612 239562
rect 275560 239498 275612 239504
rect 275466 239320 275522 239329
rect 275466 239255 275522 239264
rect 275664 79354 275692 330482
rect 275652 79348 275704 79354
rect 275652 79290 275704 79296
rect 275192 7336 275244 7342
rect 275192 7278 275244 7284
rect 275756 7274 275784 335854
rect 275848 330546 275876 335922
rect 275940 335374 275968 337640
rect 276078 337634 276106 338028
rect 276170 337736 276198 338028
rect 276262 337804 276290 338028
rect 276354 337958 276382 338028
rect 276446 337963 276474 338028
rect 276342 337952 276394 337958
rect 276342 337894 276394 337900
rect 276432 337954 276488 337963
rect 276538 337958 276566 338028
rect 276432 337889 276488 337898
rect 276526 337952 276578 337958
rect 276526 337894 276578 337900
rect 276262 337776 276336 337804
rect 276170 337708 276244 337736
rect 276078 337606 276152 337634
rect 276020 336252 276072 336258
rect 276020 336194 276072 336200
rect 275928 335368 275980 335374
rect 275928 335310 275980 335316
rect 275836 330540 275888 330546
rect 275836 330482 275888 330488
rect 276032 8226 276060 336194
rect 276124 336122 276152 337606
rect 276216 336161 276244 337708
rect 276202 336152 276258 336161
rect 276112 336116 276164 336122
rect 276202 336087 276258 336096
rect 276112 336058 276164 336064
rect 276112 335912 276164 335918
rect 276112 335854 276164 335860
rect 276202 335880 276258 335889
rect 276020 8220 276072 8226
rect 276020 8162 276072 8168
rect 275744 7268 275796 7274
rect 275744 7210 275796 7216
rect 276124 5302 276152 335854
rect 276202 335815 276258 335824
rect 276216 325694 276244 335815
rect 276308 328454 276336 337776
rect 276478 337784 276534 337793
rect 276630 337736 276658 338028
rect 276478 337719 276534 337728
rect 276492 331634 276520 337719
rect 276584 337708 276658 337736
rect 276480 331628 276532 331634
rect 276480 331570 276532 331576
rect 276308 328426 276520 328454
rect 276216 325666 276428 325694
rect 276400 235414 276428 325666
rect 276388 235408 276440 235414
rect 276388 235350 276440 235356
rect 276492 83638 276520 328426
rect 276480 83632 276532 83638
rect 276480 83574 276532 83580
rect 276584 8294 276612 337708
rect 276722 337668 276750 338028
rect 276676 337640 276750 337668
rect 276860 338014 276920 338042
rect 276676 335170 276704 337640
rect 276756 337544 276808 337550
rect 276756 337486 276808 337492
rect 276664 335164 276716 335170
rect 276664 335106 276716 335112
rect 276664 334348 276716 334354
rect 276664 334290 276716 334296
rect 276572 8288 276624 8294
rect 276572 8230 276624 8236
rect 276112 5296 276164 5302
rect 276112 5238 276164 5244
rect 276020 5024 276072 5030
rect 276020 4966 276072 4972
rect 276032 480 276060 4966
rect 276676 3534 276704 334290
rect 276768 7546 276796 337486
rect 276860 335918 276888 338014
rect 276998 337940 277026 338028
rect 276952 337912 277026 337940
rect 276952 336258 276980 337912
rect 277090 337872 277118 338028
rect 277044 337844 277118 337872
rect 276940 336252 276992 336258
rect 276940 336194 276992 336200
rect 276938 336152 276994 336161
rect 276938 336087 276994 336096
rect 276848 335912 276900 335918
rect 276952 335889 276980 336087
rect 276848 335854 276900 335860
rect 276938 335880 276994 335889
rect 276938 335815 276994 335824
rect 277044 335458 277072 337844
rect 277182 337736 277210 338028
rect 276860 335430 277072 335458
rect 277136 337708 277210 337736
rect 277274 337736 277302 338028
rect 277366 337890 277394 338028
rect 277354 337884 277406 337890
rect 277354 337826 277406 337832
rect 277274 337708 277348 337736
rect 276860 334354 276888 335430
rect 276940 335368 276992 335374
rect 276940 335310 276992 335316
rect 277032 335368 277084 335374
rect 277032 335310 277084 335316
rect 276848 334348 276900 334354
rect 276848 334290 276900 334296
rect 276756 7540 276808 7546
rect 276756 7482 276808 7488
rect 276952 7478 276980 335310
rect 277044 8158 277072 335310
rect 277032 8152 277084 8158
rect 277032 8094 277084 8100
rect 276940 7472 276992 7478
rect 276940 7414 276992 7420
rect 277136 5234 277164 337708
rect 277216 337612 277268 337618
rect 277216 337554 277268 337560
rect 277228 335918 277256 337554
rect 277216 335912 277268 335918
rect 277216 335854 277268 335860
rect 277216 335776 277268 335782
rect 277216 335718 277268 335724
rect 277228 5370 277256 335718
rect 277320 335374 277348 337708
rect 277458 337668 277486 338028
rect 277550 337736 277578 338028
rect 277642 337929 277670 338028
rect 277628 337920 277684 337929
rect 277628 337855 277684 337864
rect 277734 337736 277762 338028
rect 277826 337770 277854 338028
rect 277918 337890 277946 338028
rect 278056 338014 278116 338042
rect 277906 337884 277958 337890
rect 277906 337826 277958 337832
rect 277950 337784 278006 337793
rect 277826 337742 277900 337770
rect 277550 337708 277624 337736
rect 277458 337640 277532 337668
rect 277400 335572 277452 335578
rect 277400 335514 277452 335520
rect 277308 335368 277360 335374
rect 277308 335310 277360 335316
rect 277308 335232 277360 335238
rect 277308 335174 277360 335180
rect 277320 332217 277348 335174
rect 277306 332208 277362 332217
rect 277306 332143 277362 332152
rect 277216 5364 277268 5370
rect 277216 5306 277268 5312
rect 277124 5228 277176 5234
rect 277124 5170 277176 5176
rect 277412 5030 277440 335514
rect 277504 335374 277532 337640
rect 277596 336122 277624 337708
rect 277688 337708 277762 337736
rect 277688 337600 277716 337708
rect 277688 337572 277808 337600
rect 277676 336252 277728 336258
rect 277676 336194 277728 336200
rect 277584 336116 277636 336122
rect 277584 336058 277636 336064
rect 277584 335912 277636 335918
rect 277584 335854 277636 335860
rect 277492 335368 277544 335374
rect 277492 335310 277544 335316
rect 277596 334490 277624 335854
rect 277584 334484 277636 334490
rect 277584 334426 277636 334432
rect 277688 316034 277716 336194
rect 277780 330614 277808 337572
rect 277872 335034 277900 337742
rect 277950 337719 278006 337728
rect 277964 335481 277992 337719
rect 277950 335472 278006 335481
rect 277950 335407 278006 335416
rect 277952 335368 278004 335374
rect 277952 335310 278004 335316
rect 277860 335028 277912 335034
rect 277860 334970 277912 334976
rect 277860 330744 277912 330750
rect 277860 330686 277912 330692
rect 277768 330608 277820 330614
rect 277768 330550 277820 330556
rect 277872 316034 277900 330686
rect 277596 316006 277716 316034
rect 277780 316006 277900 316034
rect 277596 7818 277624 316006
rect 277584 7812 277636 7818
rect 277584 7754 277636 7760
rect 277780 5166 277808 316006
rect 277964 239873 277992 335310
rect 278056 330750 278084 338014
rect 278194 337770 278222 338028
rect 278286 337958 278314 338028
rect 278274 337952 278326 337958
rect 278274 337894 278326 337900
rect 278194 337742 278268 337770
rect 278136 337612 278188 337618
rect 278136 337554 278188 337560
rect 278044 330744 278096 330750
rect 278044 330686 278096 330692
rect 278044 330608 278096 330614
rect 278044 330550 278096 330556
rect 277950 239864 278006 239873
rect 277950 239799 278006 239808
rect 278056 83570 278084 330550
rect 278044 83564 278096 83570
rect 278044 83506 278096 83512
rect 278148 7886 278176 337554
rect 278240 7954 278268 337742
rect 278378 337736 278406 338028
rect 278470 337890 278498 338028
rect 278458 337884 278510 337890
rect 278458 337826 278510 337832
rect 278562 337736 278590 338028
rect 278332 337708 278406 337736
rect 278516 337708 278590 337736
rect 278332 335578 278360 337708
rect 278516 336297 278544 337708
rect 278654 337634 278682 338028
rect 278608 337606 278682 337634
rect 278502 336288 278558 336297
rect 278502 336223 278558 336232
rect 278504 336116 278556 336122
rect 278504 336058 278556 336064
rect 278320 335572 278372 335578
rect 278320 335514 278372 335520
rect 278320 335028 278372 335034
rect 278320 334970 278372 334976
rect 278332 8022 278360 334970
rect 278516 331214 278544 336058
rect 278424 331186 278544 331214
rect 278424 8090 278452 331186
rect 278608 316034 278636 337606
rect 278746 337498 278774 338028
rect 278838 337668 278866 338028
rect 278930 337736 278958 338028
rect 279022 338008 279050 338028
rect 279160 338014 279220 338042
rect 279022 337980 279096 338008
rect 278930 337708 279004 337736
rect 278838 337640 278912 337668
rect 278700 337470 278774 337498
rect 278700 336258 278728 337470
rect 278780 337408 278832 337414
rect 278780 337350 278832 337356
rect 278688 336252 278740 336258
rect 278688 336194 278740 336200
rect 278686 336152 278742 336161
rect 278686 336087 278742 336096
rect 278700 335034 278728 336087
rect 278688 335028 278740 335034
rect 278688 334970 278740 334976
rect 278516 316006 278636 316034
rect 278412 8084 278464 8090
rect 278412 8026 278464 8032
rect 278320 8016 278372 8022
rect 278320 7958 278372 7964
rect 278228 7948 278280 7954
rect 278228 7890 278280 7896
rect 278136 7880 278188 7886
rect 278136 7822 278188 7828
rect 277768 5160 277820 5166
rect 277768 5102 277820 5108
rect 278516 5030 278544 316006
rect 278792 7614 278820 337350
rect 278884 337074 278912 337640
rect 278872 337068 278924 337074
rect 278872 337010 278924 337016
rect 278872 335776 278924 335782
rect 278872 335718 278924 335724
rect 278884 325694 278912 335718
rect 278976 330478 279004 337708
rect 279068 330750 279096 337980
rect 279160 336161 279188 338014
rect 279298 337634 279326 338028
rect 279390 337770 279418 338028
rect 279482 337958 279510 338028
rect 279574 337963 279602 338028
rect 279470 337952 279522 337958
rect 279470 337894 279522 337900
rect 279560 337954 279616 337963
rect 279666 337958 279694 338028
rect 279560 337889 279616 337898
rect 279654 337952 279706 337958
rect 279654 337894 279706 337900
rect 279758 337890 279786 338028
rect 279746 337884 279798 337890
rect 279746 337826 279798 337832
rect 279514 337784 279570 337793
rect 279390 337742 279464 337770
rect 279298 337606 279372 337634
rect 279240 337544 279292 337550
rect 279240 337486 279292 337492
rect 279146 336152 279202 336161
rect 279146 336087 279202 336096
rect 279148 335640 279200 335646
rect 279146 335608 279148 335617
rect 279200 335608 279202 335617
rect 279146 335543 279202 335552
rect 279252 334529 279280 337486
rect 279238 334520 279294 334529
rect 279238 334455 279294 334464
rect 279056 330744 279108 330750
rect 279056 330686 279108 330692
rect 278964 330472 279016 330478
rect 278964 330414 279016 330420
rect 279344 325694 279372 337606
rect 279436 335374 279464 337742
rect 279850 337770 279878 338028
rect 279514 337719 279570 337728
rect 279804 337742 279878 337770
rect 279942 337770 279970 338028
rect 280034 337890 280062 338028
rect 280022 337884 280074 337890
rect 280022 337826 280074 337832
rect 279942 337742 280016 337770
rect 279424 335368 279476 335374
rect 279424 335310 279476 335316
rect 279424 335164 279476 335170
rect 279424 335106 279476 335112
rect 279436 334665 279464 335106
rect 279422 334656 279478 334665
rect 279422 334591 279478 334600
rect 278884 325666 279004 325694
rect 279344 325666 279464 325694
rect 278780 7608 278832 7614
rect 278780 7550 278832 7556
rect 278976 5098 279004 325666
rect 279436 239601 279464 325666
rect 279422 239592 279478 239601
rect 279422 239527 279478 239536
rect 279528 239465 279556 337719
rect 279608 337680 279660 337686
rect 279606 337648 279608 337657
rect 279660 337648 279662 337657
rect 279606 337583 279662 337592
rect 279804 330834 279832 337742
rect 279884 337680 279936 337686
rect 279884 337622 279936 337628
rect 279896 335617 279924 337622
rect 279882 335608 279938 335617
rect 279882 335543 279938 335552
rect 279884 335368 279936 335374
rect 279884 335310 279936 335316
rect 279620 330806 279832 330834
rect 279514 239456 279570 239465
rect 279514 239391 279570 239400
rect 279620 83502 279648 330806
rect 279700 330744 279752 330750
rect 279700 330686 279752 330692
rect 279608 83496 279660 83502
rect 279608 83438 279660 83444
rect 279712 7750 279740 330686
rect 279896 330562 279924 335310
rect 279804 330534 279924 330562
rect 279700 7744 279752 7750
rect 279700 7686 279752 7692
rect 279804 7682 279832 330534
rect 279884 330472 279936 330478
rect 279884 330414 279936 330420
rect 279896 239737 279924 330414
rect 279882 239728 279938 239737
rect 279882 239663 279938 239672
rect 279988 7857 280016 337742
rect 280126 337736 280154 338028
rect 280080 337708 280154 337736
rect 280080 335782 280108 337708
rect 280218 337668 280246 338028
rect 280172 337640 280246 337668
rect 280356 338014 280416 338042
rect 280068 335776 280120 335782
rect 280068 335718 280120 335724
rect 280172 335374 280200 337640
rect 280356 336274 280384 338014
rect 280494 337929 280522 338028
rect 280480 337920 280536 337929
rect 280586 337890 280614 338028
rect 280678 337958 280706 338028
rect 280770 337963 280798 338028
rect 280666 337952 280718 337958
rect 280666 337894 280718 337900
rect 280756 337954 280812 337963
rect 280480 337855 280536 337864
rect 280574 337884 280626 337890
rect 280756 337889 280812 337898
rect 280862 337890 280890 338028
rect 280954 337890 280982 338028
rect 280574 337826 280626 337832
rect 280850 337884 280902 337890
rect 280850 337826 280902 337832
rect 280942 337884 280994 337890
rect 280942 337826 280994 337832
rect 280710 337784 280766 337793
rect 281046 337770 281074 338028
rect 281138 337890 281166 338028
rect 281126 337884 281178 337890
rect 281126 337826 281178 337832
rect 280710 337719 280766 337728
rect 280896 337748 280948 337754
rect 280264 336246 280384 336274
rect 280264 335918 280292 336246
rect 280344 336116 280396 336122
rect 280344 336058 280396 336064
rect 280252 335912 280304 335918
rect 280252 335854 280304 335860
rect 280160 335368 280212 335374
rect 280160 335310 280212 335316
rect 280066 334792 280122 334801
rect 280066 334727 280068 334736
rect 280120 334727 280122 334736
rect 280068 334698 280120 334704
rect 280160 334688 280212 334694
rect 280160 334630 280212 334636
rect 280356 334642 280384 336058
rect 280620 335776 280672 335782
rect 280620 335718 280672 335724
rect 280434 335472 280490 335481
rect 280434 335407 280490 335416
rect 280448 334744 280476 335407
rect 280448 334716 280568 334744
rect 280172 332314 280200 334630
rect 280356 334614 280476 334642
rect 280160 332308 280212 332314
rect 280160 332250 280212 332256
rect 280344 332308 280396 332314
rect 280344 332250 280396 332256
rect 280252 331288 280304 331294
rect 280252 331230 280304 331236
rect 279974 7848 280030 7857
rect 279974 7783 280030 7792
rect 279792 7676 279844 7682
rect 279792 7618 279844 7624
rect 278964 5092 279016 5098
rect 278964 5034 279016 5040
rect 277400 5024 277452 5030
rect 277400 4966 277452 4972
rect 278504 5024 278556 5030
rect 278504 4966 278556 4972
rect 280264 4962 280292 331230
rect 280356 330478 280384 332250
rect 280344 330472 280396 330478
rect 280344 330414 280396 330420
rect 280448 5273 280476 334614
rect 280540 235278 280568 334716
rect 280528 235272 280580 235278
rect 280528 235214 280580 235220
rect 280632 177342 280660 335718
rect 280724 177410 280752 337719
rect 280896 337690 280948 337696
rect 281000 337742 281074 337770
rect 280908 335345 280936 337690
rect 280894 335336 280950 335345
rect 280894 335271 280950 335280
rect 280804 334620 280856 334626
rect 280804 334562 280856 334568
rect 280712 177404 280764 177410
rect 280712 177346 280764 177352
rect 280620 177336 280672 177342
rect 280620 177278 280672 177284
rect 280434 5264 280490 5273
rect 280434 5199 280490 5208
rect 278320 4956 278372 4962
rect 278320 4898 278372 4904
rect 280252 4956 280304 4962
rect 280252 4898 280304 4904
rect 276664 3528 276716 3534
rect 276664 3470 276716 3476
rect 277124 3052 277176 3058
rect 277124 2994 277176 3000
rect 277136 480 277164 2994
rect 278332 480 278360 4898
rect 279516 4888 279568 4894
rect 279516 4830 279568 4836
rect 279528 480 279556 4830
rect 280816 3738 280844 334562
rect 281000 331294 281028 337742
rect 281230 337736 281258 338028
rect 281184 337708 281258 337736
rect 281080 337680 281132 337686
rect 281080 337622 281132 337628
rect 280988 331288 281040 331294
rect 280988 331230 281040 331236
rect 280988 330608 281040 330614
rect 280988 330550 281040 330556
rect 280896 330472 280948 330478
rect 280896 330414 280948 330420
rect 280804 3732 280856 3738
rect 280804 3674 280856 3680
rect 280712 3596 280764 3602
rect 280712 3538 280764 3544
rect 280724 480 280752 3538
rect 280908 3262 280936 330414
rect 281000 9314 281028 330550
rect 281092 9382 281120 337622
rect 281184 335866 281212 337708
rect 281322 337668 281350 338028
rect 281414 337906 281442 338028
rect 281552 338014 281612 338042
rect 281414 337878 281488 337906
rect 281552 337890 281580 338014
rect 281276 337640 281350 337668
rect 281276 336122 281304 337640
rect 281264 336116 281316 336122
rect 281264 336058 281316 336064
rect 281184 335838 281396 335866
rect 281172 335708 281224 335714
rect 281172 335650 281224 335656
rect 281080 9376 281132 9382
rect 281080 9318 281132 9324
rect 280988 9308 281040 9314
rect 280988 9250 281040 9256
rect 281184 7585 281212 335650
rect 281368 335458 281396 335838
rect 281460 335782 281488 337878
rect 281540 337884 281592 337890
rect 281540 337826 281592 337832
rect 281690 337736 281718 338028
rect 281782 337822 281810 338028
rect 281874 337958 281902 338028
rect 281862 337952 281914 337958
rect 281862 337894 281914 337900
rect 281770 337816 281822 337822
rect 281770 337758 281822 337764
rect 281552 337708 281718 337736
rect 281448 335776 281500 335782
rect 281448 335718 281500 335724
rect 281368 335430 281488 335458
rect 281356 335300 281408 335306
rect 281356 335242 281408 335248
rect 281368 316034 281396 335242
rect 281460 335209 281488 335430
rect 281446 335200 281502 335209
rect 281446 335135 281502 335144
rect 281552 332081 281580 337708
rect 281966 337668 281994 338028
rect 282058 337770 282086 338028
rect 282150 337890 282178 338028
rect 282138 337884 282190 337890
rect 282138 337826 282190 337832
rect 282058 337742 282132 337770
rect 281920 337640 281994 337668
rect 281632 337612 281684 337618
rect 281632 337554 281684 337560
rect 281644 335073 281672 337554
rect 281724 337544 281776 337550
rect 281724 337486 281776 337492
rect 281736 335458 281764 337486
rect 281736 335430 281856 335458
rect 281724 335368 281776 335374
rect 281724 335310 281776 335316
rect 281630 335064 281686 335073
rect 281630 334999 281686 335008
rect 281632 334688 281684 334694
rect 281632 334630 281684 334636
rect 281538 332072 281594 332081
rect 281538 332007 281594 332016
rect 281644 331214 281672 334630
rect 281552 331186 281672 331214
rect 281552 330478 281580 331186
rect 281540 330472 281592 330478
rect 281540 330414 281592 330420
rect 281276 316006 281396 316034
rect 281276 7721 281304 316006
rect 281262 7712 281318 7721
rect 281262 7647 281318 7656
rect 281170 7576 281226 7585
rect 281170 7511 281226 7520
rect 281736 5137 281764 335310
rect 281828 334694 281856 335430
rect 281816 334688 281868 334694
rect 281816 334630 281868 334636
rect 281920 316034 281948 337640
rect 282000 335776 282052 335782
rect 282000 335718 282052 335724
rect 281828 316006 281948 316034
rect 281722 5128 281778 5137
rect 281722 5063 281778 5072
rect 281828 4894 281856 316006
rect 282012 9042 282040 335718
rect 282104 9178 282132 337742
rect 282242 337736 282270 338028
rect 282196 337708 282270 337736
rect 282334 337736 282362 338028
rect 282426 337872 282454 338028
rect 282518 337940 282546 338028
rect 282656 338014 282716 338042
rect 282518 337912 282592 337940
rect 282426 337844 282500 337872
rect 282334 337708 282408 337736
rect 282196 335374 282224 337708
rect 282184 335368 282236 335374
rect 282184 335310 282236 335316
rect 282182 334792 282238 334801
rect 282182 334727 282238 334736
rect 282092 9172 282144 9178
rect 282092 9114 282144 9120
rect 282000 9036 282052 9042
rect 282000 8978 282052 8984
rect 281816 4888 281868 4894
rect 281816 4830 281868 4836
rect 281908 4820 281960 4826
rect 281908 4762 281960 4768
rect 280896 3256 280948 3262
rect 280896 3198 280948 3204
rect 281920 480 281948 4762
rect 282196 2854 282224 334727
rect 282380 330698 282408 337708
rect 282472 336938 282500 337844
rect 282460 336932 282512 336938
rect 282460 336874 282512 336880
rect 282380 330670 282500 330698
rect 282368 330540 282420 330546
rect 282368 330482 282420 330488
rect 282276 330472 282328 330478
rect 282276 330414 282328 330420
rect 282288 3505 282316 330414
rect 282380 9246 282408 330482
rect 282368 9240 282420 9246
rect 282368 9182 282420 9188
rect 282472 9110 282500 330670
rect 282460 9104 282512 9110
rect 282460 9046 282512 9052
rect 282564 5001 282592 337912
rect 282656 335782 282684 338014
rect 282794 337890 282822 338028
rect 282782 337884 282834 337890
rect 282782 337826 282834 337832
rect 282886 337770 282914 338028
rect 282748 337742 282914 337770
rect 282644 335776 282696 335782
rect 282644 335718 282696 335724
rect 282644 335640 282696 335646
rect 282642 335608 282644 335617
rect 282696 335608 282698 335617
rect 282642 335543 282698 335552
rect 282642 334656 282698 334665
rect 282642 334591 282698 334600
rect 282656 334490 282684 334591
rect 282644 334484 282696 334490
rect 282644 334426 282696 334432
rect 282748 331214 282776 337742
rect 282828 337680 282880 337686
rect 282978 337668 283006 338028
rect 283070 337770 283098 338028
rect 283162 337958 283190 338028
rect 283150 337952 283202 337958
rect 283150 337894 283202 337900
rect 283254 337770 283282 338028
rect 283346 337958 283374 338028
rect 283438 337958 283466 338028
rect 283334 337952 283386 337958
rect 283334 337894 283386 337900
rect 283426 337952 283478 337958
rect 283426 337894 283478 337900
rect 283530 337770 283558 338028
rect 283622 337872 283650 338028
rect 283714 337940 283742 338028
rect 283714 337912 283788 337940
rect 283622 337844 283696 337872
rect 283070 337742 283144 337770
rect 283254 337742 283420 337770
rect 283530 337742 283604 337770
rect 282978 337640 283052 337668
rect 282828 337622 282880 337628
rect 282840 334801 282868 337622
rect 282920 336796 282972 336802
rect 282920 336738 282972 336744
rect 282932 334937 282960 336738
rect 283024 335730 283052 337640
rect 283116 336938 283144 337742
rect 283196 337680 283248 337686
rect 283196 337622 283248 337628
rect 283288 337680 283340 337686
rect 283288 337622 283340 337628
rect 283104 336932 283156 336938
rect 283104 336874 283156 336880
rect 283208 336870 283236 337622
rect 283196 336864 283248 336870
rect 283196 336806 283248 336812
rect 283300 336802 283328 337622
rect 283288 336796 283340 336802
rect 283288 336738 283340 336744
rect 283392 336274 283420 337742
rect 283472 337680 283524 337686
rect 283472 337622 283524 337628
rect 283208 336246 283420 336274
rect 283024 335702 283144 335730
rect 283012 335640 283064 335646
rect 283010 335608 283012 335617
rect 283064 335608 283066 335617
rect 283010 335543 283066 335552
rect 283012 335368 283064 335374
rect 283012 335310 283064 335316
rect 282918 334928 282974 334937
rect 282918 334863 282974 334872
rect 282826 334792 282882 334801
rect 282826 334727 282882 334736
rect 283024 331214 283052 335310
rect 283116 331945 283144 335702
rect 283102 331936 283158 331945
rect 283102 331871 283158 331880
rect 283208 331809 283236 336246
rect 283378 336152 283434 336161
rect 283378 336087 283434 336096
rect 283286 335744 283342 335753
rect 283286 335679 283342 335688
rect 283194 331800 283250 331809
rect 283194 331735 283250 331744
rect 282748 331186 282868 331214
rect 282840 316034 282868 331186
rect 282932 331186 283052 331214
rect 282932 330546 282960 331186
rect 282920 330540 282972 330546
rect 282920 330482 282972 330488
rect 283300 321554 283328 335679
rect 283392 335617 283420 336087
rect 283378 335608 283434 335617
rect 283378 335543 283434 335552
rect 283484 326398 283512 337622
rect 283576 335374 283604 337742
rect 283564 335368 283616 335374
rect 283564 335310 283616 335316
rect 283668 334665 283696 337844
rect 283760 337600 283788 337912
rect 283898 337793 283926 338028
rect 283990 337929 284018 338028
rect 284082 337958 284110 338028
rect 284070 337952 284122 337958
rect 283976 337920 284032 337929
rect 284070 337894 284122 337900
rect 284174 337890 284202 338028
rect 283976 337855 284032 337864
rect 284162 337884 284214 337890
rect 284162 337826 284214 337832
rect 283884 337784 283940 337793
rect 283884 337719 283940 337728
rect 284114 337784 284170 337793
rect 284266 337770 284294 338028
rect 284114 337719 284170 337728
rect 284220 337742 284294 337770
rect 284358 337770 284386 338028
rect 284450 337890 284478 338028
rect 284438 337884 284490 337890
rect 284438 337826 284490 337832
rect 284542 337770 284570 338028
rect 284358 337742 284432 337770
rect 283760 337572 283880 337600
rect 283748 337476 283800 337482
rect 283748 337418 283800 337424
rect 283760 336161 283788 337418
rect 283746 336152 283802 336161
rect 283746 336087 283802 336096
rect 283746 335880 283802 335889
rect 283746 335815 283802 335824
rect 283654 334656 283710 334665
rect 283654 334591 283710 334600
rect 283760 331214 283788 335815
rect 283852 333305 283880 337572
rect 284024 335368 284076 335374
rect 284024 335310 284076 335316
rect 283838 333296 283894 333305
rect 283838 333231 283894 333240
rect 283668 331186 283788 331214
rect 283472 326392 283524 326398
rect 283472 326334 283524 326340
rect 283668 321554 283696 331186
rect 283840 326392 283892 326398
rect 283840 326334 283892 326340
rect 283300 321526 283604 321554
rect 283668 321526 283788 321554
rect 282656 316006 282868 316034
rect 282550 4992 282606 5001
rect 282550 4927 282606 4936
rect 282656 4865 282684 316006
rect 283576 9654 283604 321526
rect 283564 9648 283616 9654
rect 283564 9590 283616 9596
rect 283760 9586 283788 321526
rect 283748 9580 283800 9586
rect 283748 9522 283800 9528
rect 283852 8974 283880 326334
rect 284036 240106 284064 335310
rect 284024 240100 284076 240106
rect 284024 240042 284076 240048
rect 283840 8968 283892 8974
rect 284128 8945 284156 337719
rect 284220 335374 284248 337742
rect 284404 335442 284432 337742
rect 284496 337742 284570 337770
rect 284634 337770 284662 338028
rect 284726 337906 284754 338028
rect 284832 338014 285076 338042
rect 284726 337878 284892 337906
rect 284634 337742 284800 337770
rect 284392 335436 284444 335442
rect 284392 335378 284444 335384
rect 284496 335374 284524 337742
rect 284666 335744 284722 335753
rect 284666 335679 284722 335688
rect 284574 335472 284630 335481
rect 284574 335407 284630 335416
rect 284208 335368 284260 335374
rect 284208 335310 284260 335316
rect 284484 335368 284536 335374
rect 284484 335310 284536 335316
rect 284588 331401 284616 335407
rect 284574 331392 284630 331401
rect 284574 331327 284630 331336
rect 284680 331265 284708 335679
rect 284666 331256 284722 331265
rect 284666 331191 284722 331200
rect 284300 239828 284352 239834
rect 284300 239770 284352 239776
rect 284312 11762 284340 239770
rect 284772 236978 284800 337742
rect 284864 335578 284892 337878
rect 284944 337884 284996 337890
rect 284944 337826 284996 337832
rect 284852 335572 284904 335578
rect 284852 335514 284904 335520
rect 284852 335368 284904 335374
rect 284852 335310 284904 335316
rect 284864 300150 284892 335310
rect 284956 331702 284984 337826
rect 285048 335374 285076 338014
rect 285036 335368 285088 335374
rect 285036 335310 285088 335316
rect 285036 334008 285088 334014
rect 285036 333950 285088 333956
rect 284944 331696 284996 331702
rect 284944 331638 284996 331644
rect 285048 331514 285076 333950
rect 284956 331486 285076 331514
rect 284852 300144 284904 300150
rect 284852 300086 284904 300092
rect 284760 236972 284812 236978
rect 284760 236914 284812 236920
rect 284392 89072 284444 89078
rect 284392 89014 284444 89020
rect 284300 11756 284352 11762
rect 284300 11698 284352 11704
rect 283840 8910 283892 8916
rect 284114 8936 284170 8945
rect 284114 8871 284170 8880
rect 282642 4856 282698 4865
rect 282642 4791 282698 4800
rect 283104 4752 283156 4758
rect 283104 4694 283156 4700
rect 282274 3496 282330 3505
rect 282274 3431 282330 3440
rect 282184 2848 282236 2854
rect 282184 2790 282236 2796
rect 283116 480 283144 4694
rect 284404 3482 284432 89014
rect 284956 6914 284984 331486
rect 285034 331392 285090 331401
rect 285034 331327 285090 331336
rect 285048 9450 285076 331327
rect 285140 86970 285168 388311
rect 286322 388104 286378 388113
rect 286322 388039 286378 388048
rect 285770 337920 285826 337929
rect 285770 337855 285826 337864
rect 285586 337648 285642 337657
rect 285586 337583 285642 337592
rect 285404 335572 285456 335578
rect 285404 335514 285456 335520
rect 285312 335436 285364 335442
rect 285312 335378 285364 335384
rect 285218 331256 285274 331265
rect 285218 331191 285274 331200
rect 285128 86964 285180 86970
rect 285128 86906 285180 86912
rect 285232 9518 285260 331191
rect 285324 239970 285352 335378
rect 285312 239964 285364 239970
rect 285312 239906 285364 239912
rect 285416 237182 285444 335514
rect 285496 335368 285548 335374
rect 285496 335310 285548 335316
rect 285508 237250 285536 335310
rect 285600 330614 285628 337583
rect 285784 331906 285812 337855
rect 285680 331900 285732 331906
rect 285680 331842 285732 331848
rect 285772 331900 285824 331906
rect 285772 331842 285824 331848
rect 285588 330608 285640 330614
rect 285588 330550 285640 330556
rect 285496 237244 285548 237250
rect 285496 237186 285548 237192
rect 285404 237176 285456 237182
rect 285404 237118 285456 237124
rect 285692 16574 285720 331842
rect 286336 33114 286364 388039
rect 286428 353258 286456 388894
rect 286506 388240 286562 388249
rect 286506 388175 286562 388184
rect 286416 353252 286468 353258
rect 286416 353194 286468 353200
rect 286416 337952 286468 337958
rect 286416 337894 286468 337900
rect 286428 336297 286456 337894
rect 286414 336288 286470 336297
rect 286414 336223 286470 336232
rect 286416 335640 286468 335646
rect 286416 335582 286468 335588
rect 286324 33108 286376 33114
rect 286324 33050 286376 33056
rect 285692 16546 286364 16574
rect 285404 11756 285456 11762
rect 285404 11698 285456 11704
rect 285220 9512 285272 9518
rect 285220 9454 285272 9460
rect 285036 9444 285088 9450
rect 285036 9386 285088 9392
rect 284864 6886 284984 6914
rect 284864 4146 284892 6886
rect 284852 4140 284904 4146
rect 284852 4082 284904 4088
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 285416 480 285444 11698
rect 286336 2802 286364 16546
rect 286428 2922 286456 335582
rect 286520 73166 286548 388175
rect 286612 100706 286640 390050
rect 286692 388816 286744 388822
rect 286692 388758 286744 388764
rect 286704 126954 286732 388758
rect 286796 139398 286824 390186
rect 286876 388884 286928 388890
rect 286876 388826 286928 388832
rect 286888 153202 286916 388826
rect 286980 233238 287008 390254
rect 287610 387696 287666 387705
rect 287610 387631 287666 387640
rect 287624 387190 287652 387631
rect 287612 387184 287664 387190
rect 287612 387126 287664 387132
rect 287610 387016 287666 387025
rect 287610 386951 287666 386960
rect 287624 386510 287652 386951
rect 287612 386504 287664 386510
rect 287612 386446 287664 386452
rect 287518 386336 287574 386345
rect 287518 386271 287574 386280
rect 287532 385694 287560 386271
rect 287520 385688 287572 385694
rect 287520 385630 287572 385636
rect 287610 385656 287666 385665
rect 287610 385591 287666 385600
rect 287624 385422 287652 385591
rect 287612 385416 287664 385422
rect 287612 385358 287664 385364
rect 288346 385112 288402 385121
rect 288346 385047 288348 385056
rect 288400 385047 288402 385056
rect 288348 385018 288400 385024
rect 287794 384432 287850 384441
rect 287794 384367 287850 384376
rect 287610 383072 287666 383081
rect 287610 383007 287666 383016
rect 287624 382430 287652 383007
rect 287612 382424 287664 382430
rect 287612 382366 287664 382372
rect 287702 371376 287758 371385
rect 287702 371311 287758 371320
rect 287610 370152 287666 370161
rect 287610 370087 287666 370096
rect 287624 369986 287652 370087
rect 287612 369980 287664 369986
rect 287612 369922 287664 369928
rect 287610 368792 287666 368801
rect 287610 368727 287666 368736
rect 287624 368626 287652 368727
rect 287612 368620 287664 368626
rect 287612 368562 287664 368568
rect 287518 366888 287574 366897
rect 287518 366823 287574 366832
rect 287426 366208 287482 366217
rect 287426 366143 287482 366152
rect 287334 365528 287390 365537
rect 287334 365463 287390 365472
rect 287150 364304 287206 364313
rect 287150 364239 287206 364248
rect 287164 362982 287192 364239
rect 287152 362976 287204 362982
rect 287152 362918 287204 362924
rect 287348 358290 287376 365463
rect 287336 358284 287388 358290
rect 287336 358226 287388 358232
rect 287440 358222 287468 366143
rect 287428 358216 287480 358222
rect 287428 358158 287480 358164
rect 287532 358154 287560 366823
rect 287520 358148 287572 358154
rect 287520 358090 287572 358096
rect 287716 358086 287744 371311
rect 287704 358080 287756 358086
rect 287704 358022 287756 358028
rect 287610 357096 287666 357105
rect 287610 357031 287666 357040
rect 287426 356416 287482 356425
rect 287426 356351 287482 356360
rect 287440 356114 287468 356351
rect 287624 356318 287652 357031
rect 287612 356312 287664 356318
rect 287612 356254 287664 356260
rect 287428 356108 287480 356114
rect 287428 356050 287480 356056
rect 287702 354512 287758 354521
rect 287702 354447 287758 354456
rect 287610 353832 287666 353841
rect 287610 353767 287612 353776
rect 287664 353767 287666 353776
rect 287612 353738 287664 353744
rect 287716 350334 287744 354447
rect 287704 350328 287756 350334
rect 287704 350270 287756 350276
rect 287610 347304 287666 347313
rect 287610 347239 287666 347248
rect 287624 346458 287652 347239
rect 287612 346452 287664 346458
rect 287612 346394 287664 346400
rect 287334 346080 287390 346089
rect 287334 346015 287390 346024
rect 287348 345166 287376 346015
rect 287336 345160 287388 345166
rect 287336 345102 287388 345108
rect 287518 344176 287574 344185
rect 287518 344111 287574 344120
rect 287532 335850 287560 344111
rect 287610 342816 287666 342825
rect 287610 342751 287666 342760
rect 287624 335918 287652 342751
rect 287702 341456 287758 341465
rect 287702 341391 287758 341400
rect 287716 340950 287744 341391
rect 287704 340944 287756 340950
rect 287704 340886 287756 340892
rect 287612 335912 287664 335918
rect 287612 335854 287664 335860
rect 287520 335844 287572 335850
rect 287520 335786 287572 335792
rect 287704 334076 287756 334082
rect 287704 334018 287756 334024
rect 287060 238196 287112 238202
rect 287060 238138 287112 238144
rect 286968 233232 287020 233238
rect 286968 233174 287020 233180
rect 286876 153196 286928 153202
rect 286876 153138 286928 153144
rect 286784 139392 286836 139398
rect 286784 139334 286836 139340
rect 286692 126948 286744 126954
rect 286692 126890 286744 126896
rect 286600 100700 286652 100706
rect 286600 100642 286652 100648
rect 286508 73160 286560 73166
rect 286508 73102 286560 73108
rect 287072 16574 287100 238138
rect 287072 16546 287376 16574
rect 286416 2916 286468 2922
rect 286416 2858 286468 2864
rect 286336 2774 286640 2802
rect 286612 480 286640 2774
rect 287348 490 287376 16546
rect 287716 3602 287744 334018
rect 287808 239154 287836 384367
rect 288346 383752 288402 383761
rect 288346 383687 288348 383696
rect 288400 383687 288402 383696
rect 288348 383658 288400 383664
rect 288346 382392 288402 382401
rect 288346 382327 288348 382336
rect 288400 382327 288402 382336
rect 288348 382298 288400 382304
rect 288162 381848 288218 381857
rect 288162 381783 288218 381792
rect 288176 381002 288204 381783
rect 288346 381168 288402 381177
rect 288346 381103 288402 381112
rect 288164 380996 288216 381002
rect 288164 380938 288216 380944
rect 288360 380934 288388 381103
rect 288348 380928 288400 380934
rect 288348 380870 288400 380876
rect 288254 380488 288310 380497
rect 288254 380423 288310 380432
rect 288268 379574 288296 380423
rect 288346 379808 288402 379817
rect 288346 379743 288348 379752
rect 288400 379743 288402 379752
rect 288348 379714 288400 379720
rect 288256 379568 288308 379574
rect 288256 379510 288308 379516
rect 288254 379264 288310 379273
rect 288254 379199 288310 379208
rect 288268 378214 288296 379199
rect 288346 378584 288402 378593
rect 288346 378519 288402 378528
rect 288360 378282 288388 378519
rect 288348 378276 288400 378282
rect 288348 378218 288400 378224
rect 288256 378208 288308 378214
rect 288256 378150 288308 378156
rect 288254 377904 288310 377913
rect 288254 377839 288310 377848
rect 288268 376786 288296 377839
rect 288346 377224 288402 377233
rect 288346 377159 288402 377168
rect 288360 376854 288388 377159
rect 288348 376848 288400 376854
rect 288348 376790 288400 376796
rect 288256 376780 288308 376786
rect 288256 376722 288308 376728
rect 288346 376544 288402 376553
rect 288346 376479 288402 376488
rect 288162 376000 288218 376009
rect 288162 375935 288218 375944
rect 288176 375494 288204 375935
rect 288164 375488 288216 375494
rect 288164 375430 288216 375436
rect 288360 375426 288388 376479
rect 288348 375420 288400 375426
rect 288348 375362 288400 375368
rect 288346 375320 288402 375329
rect 288346 375255 288402 375264
rect 288162 374640 288218 374649
rect 288162 374575 288218 374584
rect 288176 374134 288204 374575
rect 288164 374128 288216 374134
rect 288164 374070 288216 374076
rect 288360 374066 288388 375255
rect 288348 374060 288400 374066
rect 288348 374002 288400 374008
rect 288254 373960 288310 373969
rect 288254 373895 288310 373904
rect 288162 373416 288218 373425
rect 288162 373351 288218 373360
rect 288176 372706 288204 373351
rect 288164 372700 288216 372706
rect 288164 372642 288216 372648
rect 288268 372638 288296 373895
rect 288348 372768 288400 372774
rect 288346 372736 288348 372745
rect 288400 372736 288402 372745
rect 288346 372671 288402 372680
rect 288256 372632 288308 372638
rect 288256 372574 288308 372580
rect 288254 372056 288310 372065
rect 288254 371991 288310 372000
rect 288268 371278 288296 371991
rect 288256 371272 288308 371278
rect 288256 371214 288308 371220
rect 288346 370696 288402 370705
rect 288346 370631 288402 370640
rect 288360 369918 288388 370631
rect 288348 369912 288400 369918
rect 288348 369854 288400 369860
rect 288254 369472 288310 369481
rect 288254 369407 288310 369416
rect 288268 368558 288296 369407
rect 288256 368552 288308 368558
rect 288256 368494 288308 368500
rect 288346 368112 288402 368121
rect 288346 368047 288402 368056
rect 287978 367568 288034 367577
rect 287978 367503 288034 367512
rect 287992 367198 288020 367503
rect 287980 367192 288032 367198
rect 287980 367134 288032 367140
rect 288360 367130 288388 368047
rect 288348 367124 288400 367130
rect 288348 367066 288400 367072
rect 288346 364848 288402 364857
rect 288346 364783 288402 364792
rect 288360 364410 288388 364783
rect 288348 364404 288400 364410
rect 288348 364346 288400 364352
rect 288162 363624 288218 363633
rect 288162 363559 288218 363568
rect 288176 363050 288204 363559
rect 288164 363044 288216 363050
rect 288164 362986 288216 362992
rect 288162 362944 288218 362953
rect 288162 362879 288218 362888
rect 288176 361622 288204 362879
rect 288254 362264 288310 362273
rect 288254 362199 288310 362208
rect 288268 361758 288296 362199
rect 288256 361752 288308 361758
rect 288256 361694 288308 361700
rect 288346 361720 288402 361729
rect 288346 361655 288348 361664
rect 288400 361655 288402 361664
rect 288348 361626 288400 361632
rect 288164 361616 288216 361622
rect 288164 361558 288216 361564
rect 288162 361040 288218 361049
rect 288162 360975 288218 360984
rect 288176 360330 288204 360975
rect 288346 360360 288402 360369
rect 288164 360324 288216 360330
rect 288346 360295 288402 360304
rect 288164 360266 288216 360272
rect 288360 360262 288388 360295
rect 288348 360256 288400 360262
rect 288348 360198 288400 360204
rect 288346 359680 288402 359689
rect 288346 359615 288402 359624
rect 288162 359000 288218 359009
rect 288162 358935 288218 358944
rect 288176 358358 288204 358935
rect 288360 358834 288388 359615
rect 288348 358828 288400 358834
rect 288348 358770 288400 358776
rect 288254 358456 288310 358465
rect 288254 358391 288310 358400
rect 288164 358352 288216 358358
rect 288164 358294 288216 358300
rect 288268 357542 288296 358391
rect 288346 357776 288402 357785
rect 288346 357711 288402 357720
rect 288256 357536 288308 357542
rect 288256 357478 288308 357484
rect 288360 357474 288388 357711
rect 288348 357468 288400 357474
rect 288348 357410 288400 357416
rect 288346 355872 288402 355881
rect 288346 355807 288402 355816
rect 287978 355192 288034 355201
rect 287978 355127 288034 355136
rect 287992 354822 288020 355127
rect 287980 354816 288032 354822
rect 287980 354758 288032 354764
rect 288360 354754 288388 355807
rect 288348 354748 288400 354754
rect 288348 354690 288400 354696
rect 287978 353152 288034 353161
rect 287978 353087 288034 353096
rect 287886 352608 287942 352617
rect 287886 352543 287942 352552
rect 287796 239148 287848 239154
rect 287796 239090 287848 239096
rect 287900 237318 287928 352543
rect 287992 350418 288020 353087
rect 288348 351960 288400 351966
rect 288346 351928 288348 351937
rect 288400 351928 288402 351937
rect 288346 351863 288402 351872
rect 288070 351248 288126 351257
rect 288070 351183 288126 351192
rect 288084 350606 288112 351183
rect 288348 350668 288400 350674
rect 288348 350610 288400 350616
rect 288072 350600 288124 350606
rect 288360 350577 288388 350610
rect 288072 350542 288124 350548
rect 288346 350568 288402 350577
rect 288346 350503 288402 350512
rect 287992 350390 288112 350418
rect 287980 350328 288032 350334
rect 287980 350270 288032 350276
rect 287992 238202 288020 350270
rect 288084 238270 288112 350390
rect 288346 350024 288402 350033
rect 288346 349959 288402 349968
rect 288254 349344 288310 349353
rect 288254 349279 288256 349288
rect 288308 349279 288310 349288
rect 288256 349250 288308 349256
rect 288360 349178 288388 349959
rect 288348 349172 288400 349178
rect 288348 349114 288400 349120
rect 288346 348664 288402 348673
rect 288346 348599 288402 348608
rect 288254 347984 288310 347993
rect 288254 347919 288256 347928
rect 288308 347919 288310 347928
rect 288256 347890 288308 347896
rect 288360 347818 288388 348599
rect 288348 347812 288400 347818
rect 288348 347754 288400 347760
rect 288346 346760 288402 346769
rect 288346 346695 288348 346704
rect 288400 346695 288402 346704
rect 288348 346666 288400 346672
rect 288346 345400 288402 345409
rect 288346 345335 288402 345344
rect 288360 345098 288388 345335
rect 288348 345092 288400 345098
rect 288348 345034 288400 345040
rect 288162 344720 288218 344729
rect 288162 344655 288218 344664
rect 288176 343738 288204 344655
rect 288164 343732 288216 343738
rect 288164 343674 288216 343680
rect 288346 343496 288402 343505
rect 288346 343431 288402 343440
rect 288360 342310 288388 343431
rect 288348 342304 288400 342310
rect 288348 342246 288400 342252
rect 288162 342136 288218 342145
rect 288162 342071 288218 342080
rect 288176 336002 288204 342071
rect 288348 341012 288400 341018
rect 288348 340954 288400 340960
rect 288360 340921 288388 340954
rect 288346 340912 288402 340921
rect 288346 340847 288402 340856
rect 288254 340232 288310 340241
rect 288254 340167 288310 340176
rect 288268 339522 288296 340167
rect 288348 339584 288400 339590
rect 288346 339552 288348 339561
rect 288400 339552 288402 339561
rect 288256 339516 288308 339522
rect 288346 339487 288402 339496
rect 288256 339458 288308 339464
rect 288254 338872 288310 338881
rect 288254 338807 288310 338816
rect 288268 338230 288296 338807
rect 288346 338328 288402 338337
rect 288346 338263 288402 338272
rect 288256 338224 288308 338230
rect 288256 338166 288308 338172
rect 288360 338162 288388 338263
rect 288348 338156 288400 338162
rect 288348 338098 288400 338104
rect 288176 335974 288388 336002
rect 288256 335912 288308 335918
rect 288256 335854 288308 335860
rect 288164 335844 288216 335850
rect 288164 335786 288216 335792
rect 288176 238882 288204 335786
rect 288164 238876 288216 238882
rect 288164 238818 288216 238824
rect 288268 238746 288296 335854
rect 288256 238740 288308 238746
rect 288256 238682 288308 238688
rect 288072 238264 288124 238270
rect 288072 238206 288124 238212
rect 287980 238196 288032 238202
rect 287980 238138 288032 238144
rect 288360 237998 288388 335974
rect 289004 320890 289032 390390
rect 289096 365702 289124 390458
rect 537484 390380 537536 390386
rect 537484 390322 537536 390328
rect 289728 390176 289780 390182
rect 289728 390118 289780 390124
rect 289636 390040 289688 390046
rect 289636 389982 289688 389988
rect 289084 365696 289136 365702
rect 289084 365638 289136 365644
rect 289084 335776 289136 335782
rect 289084 335718 289136 335724
rect 288992 320884 289044 320890
rect 288992 320826 289044 320832
rect 288348 237992 288400 237998
rect 288348 237934 288400 237940
rect 287888 237312 287940 237318
rect 287888 237254 287940 237260
rect 287704 3596 287756 3602
rect 287704 3538 287756 3544
rect 288992 3596 289044 3602
rect 288992 3538 289044 3544
rect 287624 598 287836 626
rect 287624 490 287652 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 462 287652 490
rect 287808 480 287836 598
rect 289004 480 289032 3538
rect 289096 3058 289124 335718
rect 289176 335708 289228 335714
rect 289176 335650 289228 335656
rect 289084 3052 289136 3058
rect 289084 2994 289136 3000
rect 289188 2990 289216 335650
rect 289268 335640 289320 335646
rect 289268 335582 289320 335588
rect 289280 3194 289308 335582
rect 289360 334144 289412 334150
rect 289360 334086 289412 334092
rect 289372 3602 289400 334086
rect 289544 331628 289596 331634
rect 289544 331570 289596 331576
rect 289452 331424 289504 331430
rect 289452 331366 289504 331372
rect 289464 4010 289492 331366
rect 289452 4004 289504 4010
rect 289452 3946 289504 3952
rect 289556 3806 289584 331570
rect 289648 179382 289676 389982
rect 289740 219434 289768 390118
rect 292212 389632 292264 389638
rect 292212 389574 292264 389580
rect 311162 389600 311218 389609
rect 292120 389564 292172 389570
rect 292120 389506 292172 389512
rect 292028 389428 292080 389434
rect 292028 389370 292080 389376
rect 290832 379772 290884 379778
rect 290832 379714 290884 379720
rect 290554 336560 290610 336569
rect 290554 336495 290610 336504
rect 290464 335368 290516 335374
rect 290464 335310 290516 335316
rect 289728 219428 289780 219434
rect 289728 219370 289780 219376
rect 289636 179376 289688 179382
rect 289636 179318 289688 179324
rect 290188 5500 290240 5506
rect 290188 5442 290240 5448
rect 289544 3800 289596 3806
rect 289544 3742 289596 3748
rect 289360 3596 289412 3602
rect 289360 3538 289412 3544
rect 289268 3188 289320 3194
rect 289268 3130 289320 3136
rect 289176 2984 289228 2990
rect 289176 2926 289228 2932
rect 290200 480 290228 5442
rect 290476 4078 290504 335310
rect 290568 5438 290596 336495
rect 290648 331560 290700 331566
rect 290648 331502 290700 331508
rect 290556 5432 290608 5438
rect 290556 5374 290608 5380
rect 290464 4072 290516 4078
rect 290464 4014 290516 4020
rect 290660 3670 290688 331502
rect 290740 331356 290792 331362
rect 290740 331298 290792 331304
rect 290752 3777 290780 331298
rect 290844 245614 290872 379714
rect 291844 335572 291896 335578
rect 291844 335514 291896 335520
rect 290924 331492 290976 331498
rect 290924 331434 290976 331440
rect 290832 245608 290884 245614
rect 290832 245550 290884 245556
rect 290738 3768 290794 3777
rect 290738 3703 290794 3712
rect 290648 3664 290700 3670
rect 290936 3641 290964 331434
rect 291200 331288 291252 331294
rect 291200 331230 291252 331236
rect 291212 16574 291240 331230
rect 291212 16546 291424 16574
rect 290648 3606 290700 3612
rect 290922 3632 290978 3641
rect 290922 3567 290978 3576
rect 291396 480 291424 16546
rect 291856 3942 291884 335514
rect 291936 335436 291988 335442
rect 291936 335378 291988 335384
rect 291948 4758 291976 335378
rect 292040 238105 292068 389370
rect 292132 238474 292160 389506
rect 292120 238468 292172 238474
rect 292120 238410 292172 238416
rect 292026 238096 292082 238105
rect 292026 238031 292082 238040
rect 292224 237833 292252 389574
rect 311162 389535 311218 389544
rect 298836 389496 298888 389502
rect 298836 389438 298888 389444
rect 294604 389360 294656 389366
rect 294604 389302 294656 389308
rect 293316 389224 293368 389230
rect 293316 389166 293368 389172
rect 293222 336424 293278 336433
rect 293222 336359 293278 336368
rect 292580 334212 292632 334218
rect 292580 334154 292632 334160
rect 292304 331696 292356 331702
rect 292304 331638 292356 331644
rect 292210 237824 292266 237833
rect 292210 237759 292266 237768
rect 292316 236638 292344 331638
rect 292396 300144 292448 300150
rect 292396 300086 292448 300092
rect 292304 236632 292356 236638
rect 292304 236574 292356 236580
rect 292408 236570 292436 300086
rect 292396 236564 292448 236570
rect 292396 236506 292448 236512
rect 291936 4752 291988 4758
rect 291936 4694 291988 4700
rect 291844 3936 291896 3942
rect 291844 3878 291896 3884
rect 292592 480 292620 334154
rect 293236 5506 293264 336359
rect 293328 237726 293356 389166
rect 293408 386504 293460 386510
rect 293408 386446 293460 386452
rect 293420 238377 293448 386446
rect 293500 385688 293552 385694
rect 293500 385630 293552 385636
rect 293406 238368 293462 238377
rect 293512 238338 293540 385630
rect 293592 385416 293644 385422
rect 293592 385358 293644 385364
rect 293604 238406 293632 385358
rect 293592 238400 293644 238406
rect 293592 238342 293644 238348
rect 293406 238303 293462 238312
rect 293500 238332 293552 238338
rect 293500 238274 293552 238280
rect 294616 237930 294644 389302
rect 294696 387184 294748 387190
rect 294696 387126 294748 387132
rect 294708 238241 294736 387126
rect 298744 386708 298796 386714
rect 298744 386650 298796 386656
rect 295984 386640 296036 386646
rect 295984 386582 296036 386588
rect 294880 382424 294932 382430
rect 294880 382366 294932 382372
rect 294788 382356 294840 382362
rect 294788 382298 294840 382304
rect 294694 238232 294750 238241
rect 294694 238167 294750 238176
rect 294604 237924 294656 237930
rect 294604 237866 294656 237872
rect 294800 237862 294828 382298
rect 294788 237856 294840 237862
rect 294788 237798 294840 237804
rect 294892 237794 294920 382366
rect 294972 346724 295024 346730
rect 294972 346666 295024 346672
rect 294880 237788 294932 237794
rect 294880 237730 294932 237736
rect 293316 237720 293368 237726
rect 293316 237662 293368 237668
rect 294984 236774 295012 346666
rect 295064 346452 295116 346458
rect 295064 346394 295116 346400
rect 295076 238542 295104 346394
rect 295156 343732 295208 343738
rect 295156 343674 295208 343680
rect 295168 238950 295196 343674
rect 295156 238944 295208 238950
rect 295156 238886 295208 238892
rect 295064 238536 295116 238542
rect 295064 238478 295116 238484
rect 294972 236768 295024 236774
rect 294972 236710 295024 236716
rect 295996 6866 296024 386582
rect 297456 357536 297508 357542
rect 297456 357478 297508 357484
rect 297364 357468 297416 357474
rect 297364 357410 297416 357416
rect 296260 356312 296312 356318
rect 296260 356254 296312 356260
rect 296168 356108 296220 356114
rect 296168 356050 296220 356056
rect 296076 335912 296128 335918
rect 296076 335854 296128 335860
rect 296088 16574 296116 335854
rect 296180 235822 296208 356050
rect 296272 235890 296300 356254
rect 296352 353796 296404 353802
rect 296352 353738 296404 353744
rect 296364 237114 296392 353738
rect 296444 349308 296496 349314
rect 296444 349250 296496 349256
rect 296352 237108 296404 237114
rect 296352 237050 296404 237056
rect 296456 236910 296484 349250
rect 296536 347948 296588 347954
rect 296536 347890 296588 347896
rect 296444 236904 296496 236910
rect 296444 236846 296496 236852
rect 296548 236706 296576 347890
rect 296628 339584 296680 339590
rect 296628 339526 296680 339532
rect 296536 236700 296588 236706
rect 296536 236642 296588 236648
rect 296260 235884 296312 235890
rect 296260 235826 296312 235832
rect 296168 235816 296220 235822
rect 296168 235758 296220 235764
rect 296640 235754 296668 339526
rect 297376 235958 297404 357410
rect 297468 237017 297496 357478
rect 297640 341012 297692 341018
rect 297640 340954 297692 340960
rect 297548 340944 297600 340950
rect 297548 340886 297600 340892
rect 297454 237008 297510 237017
rect 297454 236943 297510 236952
rect 297560 236434 297588 340886
rect 297548 236428 297600 236434
rect 297548 236370 297600 236376
rect 297652 236366 297680 340954
rect 297732 339516 297784 339522
rect 297732 339458 297784 339464
rect 297640 236360 297692 236366
rect 297640 236302 297692 236308
rect 297744 236298 297772 339458
rect 298100 331764 298152 331770
rect 298100 331706 298152 331712
rect 297732 236292 297784 236298
rect 297732 236234 297784 236240
rect 297364 235952 297416 235958
rect 297364 235894 297416 235900
rect 296628 235748 296680 235754
rect 296628 235690 296680 235696
rect 296088 16546 296208 16574
rect 294880 6860 294932 6866
rect 294880 6802 294932 6808
rect 295984 6860 296036 6866
rect 295984 6802 296036 6808
rect 293132 5500 293184 5506
rect 293132 5442 293184 5448
rect 293224 5500 293276 5506
rect 293224 5442 293276 5448
rect 293144 4758 293172 5442
rect 293132 4752 293184 4758
rect 293132 4694 293184 4700
rect 293684 4752 293736 4758
rect 293684 4694 293736 4700
rect 293696 480 293724 4694
rect 294892 480 294920 6802
rect 296180 4010 296208 16546
rect 297272 4208 297324 4214
rect 297272 4150 297324 4156
rect 296168 4004 296220 4010
rect 296168 3946 296220 3952
rect 296076 3596 296128 3602
rect 296076 3538 296128 3544
rect 296088 480 296116 3538
rect 297284 480 297312 4150
rect 298112 490 298140 331706
rect 298756 193186 298784 386650
rect 298848 236745 298876 389438
rect 299020 383716 299072 383722
rect 299020 383658 299072 383664
rect 298928 380996 298980 381002
rect 298928 380938 298980 380944
rect 298834 236736 298890 236745
rect 298834 236671 298890 236680
rect 298940 236230 298968 380938
rect 299032 236881 299060 383658
rect 300216 354816 300268 354822
rect 300216 354758 300268 354764
rect 299112 347812 299164 347818
rect 299112 347754 299164 347760
rect 299124 238678 299152 347754
rect 299296 345160 299348 345166
rect 299296 345102 299348 345108
rect 299204 342304 299256 342310
rect 299204 342246 299256 342252
rect 299112 238672 299164 238678
rect 299112 238614 299164 238620
rect 299018 236872 299074 236881
rect 299018 236807 299074 236816
rect 299216 236502 299244 342246
rect 299308 239018 299336 345102
rect 300124 335980 300176 335986
rect 300124 335922 300176 335928
rect 299296 239012 299348 239018
rect 299296 238954 299348 238960
rect 299204 236496 299256 236502
rect 299204 236438 299256 236444
rect 298928 236224 298980 236230
rect 298928 236166 298980 236172
rect 298744 193180 298796 193186
rect 298744 193122 298796 193128
rect 300136 4146 300164 335922
rect 300228 237046 300256 354758
rect 300400 351960 300452 351966
rect 300400 351902 300452 351908
rect 300308 350668 300360 350674
rect 300308 350610 300360 350616
rect 300216 237040 300268 237046
rect 300216 236982 300268 236988
rect 300320 236842 300348 350610
rect 300412 238814 300440 351902
rect 300492 349172 300544 349178
rect 300492 349114 300544 349120
rect 300400 238808 300452 238814
rect 300400 238750 300452 238756
rect 300504 238610 300532 349114
rect 300584 338224 300636 338230
rect 300584 338166 300636 338172
rect 300596 239086 300624 338166
rect 309782 336288 309838 336297
rect 309782 336223 309838 336232
rect 308402 336016 308458 336025
rect 308402 335951 308458 335960
rect 306380 332648 306432 332654
rect 306380 332590 306432 332596
rect 300860 331832 300912 331838
rect 300860 331774 300912 331780
rect 300584 239080 300636 239086
rect 300584 239022 300636 239028
rect 300492 238604 300544 238610
rect 300492 238546 300544 238552
rect 300308 236836 300360 236842
rect 300308 236778 300360 236784
rect 300872 16574 300900 331774
rect 302240 87848 302292 87854
rect 302240 87790 302292 87796
rect 302252 16574 302280 87790
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 300768 4276 300820 4282
rect 300768 4218 300820 4224
rect 299664 4140 299716 4146
rect 299664 4082 299716 4088
rect 300124 4140 300176 4146
rect 300124 4082 300176 4088
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 4082
rect 300780 480 300808 4218
rect 301516 490 301544 16546
rect 301792 598 302004 626
rect 301792 490 301820 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 462 301820 490
rect 301976 480 302004 598
rect 303172 480 303200 16546
rect 304356 4344 304408 4350
rect 304356 4286 304408 4292
rect 304368 480 304396 4286
rect 305552 3324 305604 3330
rect 305552 3266 305604 3272
rect 305564 480 305592 3266
rect 306392 490 306420 332590
rect 307760 332580 307812 332586
rect 307760 332522 307812 332528
rect 307772 3330 307800 332522
rect 307852 85128 307904 85134
rect 307852 85070 307904 85076
rect 307864 16574 307892 85070
rect 307864 16546 307984 16574
rect 307760 3324 307812 3330
rect 307760 3266 307812 3272
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 16546
rect 308416 3448 308444 335951
rect 309140 334280 309192 334286
rect 309140 334222 309192 334228
rect 309152 6914 309180 334222
rect 309796 16574 309824 336223
rect 311176 20670 311204 389535
rect 438124 385076 438176 385082
rect 438124 385018 438176 385024
rect 370504 379568 370556 379574
rect 370504 379510 370556 379516
rect 353944 378276 353996 378282
rect 353944 378218 353996 378224
rect 349804 376848 349856 376854
rect 349804 376790 349856 376796
rect 342904 375488 342956 375494
rect 342904 375430 342956 375436
rect 338764 374128 338816 374134
rect 338764 374070 338816 374076
rect 319442 336152 319498 336161
rect 319442 336087 319498 336096
rect 316132 332784 316184 332790
rect 316132 332726 316184 332732
rect 313280 332716 313332 332722
rect 313280 332658 313332 332664
rect 311900 332512 311952 332518
rect 311900 332454 311952 332460
rect 311164 20664 311216 20670
rect 311164 20606 311216 20612
rect 311912 16574 311940 332454
rect 313292 16574 313320 332658
rect 309796 16546 309916 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 309152 6886 309824 6914
rect 308416 3420 309180 3448
rect 309152 3330 309180 3420
rect 309048 3324 309100 3330
rect 309048 3266 309100 3272
rect 309140 3324 309192 3330
rect 309140 3266 309192 3272
rect 309060 480 309088 3266
rect 309796 490 309824 6886
rect 309888 3369 309916 16546
rect 311440 4412 311492 4418
rect 311440 4354 311492 4360
rect 309874 3360 309930 3369
rect 309874 3295 309930 3304
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 4354
rect 312188 490 312216 16546
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 16546
rect 316144 11762 316172 332726
rect 318800 332444 318852 332450
rect 318800 332386 318852 332392
rect 318812 16574 318840 332386
rect 318812 16546 319392 16574
rect 316132 11756 316184 11762
rect 316132 11698 316184 11704
rect 317328 11756 317380 11762
rect 317328 11698 317380 11704
rect 315028 4480 315080 4486
rect 315028 4422 315080 4428
rect 315040 480 315068 4422
rect 316224 3460 316276 3466
rect 316224 3402 316276 3408
rect 316236 480 316264 3402
rect 317340 480 317368 11698
rect 318524 4548 318576 4554
rect 318524 4490 318576 4496
rect 318536 480 318564 4490
rect 319364 3346 319392 16546
rect 319456 3466 319484 336087
rect 325700 334416 325752 334422
rect 325700 334358 325752 334364
rect 320180 80912 320232 80918
rect 320180 80854 320232 80860
rect 320192 16574 320220 80854
rect 325712 16574 325740 334358
rect 329840 332376 329892 332382
rect 329840 332318 329892 332324
rect 329852 16574 329880 332318
rect 338776 322862 338804 374070
rect 340144 374060 340196 374066
rect 340144 374002 340196 374008
rect 338764 322856 338816 322862
rect 338764 322798 338816 322804
rect 340156 322794 340184 374002
rect 340972 332920 341024 332926
rect 340972 332862 341024 332868
rect 340144 322788 340196 322794
rect 340144 322730 340196 322736
rect 332600 85060 332652 85066
rect 332600 85002 332652 85008
rect 320192 16546 320496 16574
rect 325712 16546 326384 16574
rect 329852 16546 330432 16574
rect 319444 3460 319496 3466
rect 319444 3402 319496 3408
rect 319364 3318 319760 3346
rect 319732 480 319760 3318
rect 320468 490 320496 16546
rect 324320 10804 324372 10810
rect 324320 10746 324372 10752
rect 322112 5568 322164 5574
rect 322112 5510 322164 5516
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 5510
rect 324332 2854 324360 10746
rect 324412 5636 324464 5642
rect 324412 5578 324464 5584
rect 323308 2848 323360 2854
rect 323308 2790 323360 2796
rect 324320 2848 324372 2854
rect 324320 2790 324372 2796
rect 323320 480 323348 2790
rect 324424 480 324452 5578
rect 325608 2848 325660 2854
rect 325608 2790 325660 2796
rect 325620 480 325648 2790
rect 326356 490 326384 16546
rect 328736 10736 328788 10742
rect 328736 10678 328788 10684
rect 328000 5704 328052 5710
rect 328000 5646 328052 5652
rect 326632 598 326844 626
rect 326632 490 326660 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 462 326660 490
rect 326816 480 326844 598
rect 328012 480 328040 5646
rect 328748 490 328776 10678
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 16546
rect 331588 5772 331640 5778
rect 331588 5714 331640 5720
rect 331600 480 331628 5714
rect 332612 2854 332640 85002
rect 340984 16590 341012 332862
rect 342916 322726 342944 375430
rect 345664 375420 345716 375426
rect 345664 375362 345716 375368
rect 342904 322720 342956 322726
rect 342904 322662 342956 322668
rect 345676 322658 345704 375362
rect 347780 336728 347832 336734
rect 347780 336670 347832 336676
rect 345664 322652 345716 322658
rect 345664 322594 345716 322600
rect 345020 80844 345072 80850
rect 345020 80786 345072 80792
rect 340972 16584 341024 16590
rect 340972 16526 341024 16532
rect 342168 16584 342220 16590
rect 345032 16574 345060 80786
rect 347792 16574 347820 336670
rect 349816 322590 349844 376790
rect 352656 376780 352708 376786
rect 352656 376722 352708 376728
rect 352564 345092 352616 345098
rect 352564 345034 352616 345040
rect 349804 322584 349856 322590
rect 349804 322526 349856 322532
rect 352576 237658 352604 345034
rect 352668 322454 352696 376722
rect 353956 322522 353984 378218
rect 356704 378208 356756 378214
rect 356704 378150 356756 378156
rect 354680 336660 354732 336666
rect 354680 336602 354732 336608
rect 353944 322516 353996 322522
rect 353944 322458 353996 322464
rect 352656 322448 352708 322454
rect 352656 322390 352708 322396
rect 352564 237652 352616 237658
rect 352564 237594 352616 237600
rect 349160 84992 349212 84998
rect 349160 84934 349212 84940
rect 349172 16574 349200 84934
rect 354692 16574 354720 336602
rect 356060 332852 356112 332858
rect 356060 332794 356112 332800
rect 356072 16574 356100 332794
rect 356716 322386 356744 378150
rect 363604 363044 363656 363050
rect 363604 362986 363656 362992
rect 360844 361752 360896 361758
rect 360844 361694 360896 361700
rect 359464 360324 359516 360330
rect 359464 360266 359516 360272
rect 358820 332988 358872 332994
rect 358820 332930 358872 332936
rect 357440 332308 357492 332314
rect 357440 332250 357492 332256
rect 356704 322380 356756 322386
rect 356704 322322 356756 322328
rect 345032 16546 345336 16574
rect 347792 16546 348096 16574
rect 349172 16546 349292 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 342168 16526 342220 16532
rect 332692 10668 332744 10674
rect 332692 10610 332744 10616
rect 332600 2848 332652 2854
rect 332600 2790 332652 2796
rect 332704 480 332732 10610
rect 336280 10600 336332 10606
rect 336280 10542 336332 10548
rect 335084 5840 335136 5846
rect 335084 5782 335136 5788
rect 333888 2848 333940 2854
rect 333888 2790 333940 2796
rect 333900 480 333928 2790
rect 335096 480 335124 5782
rect 336292 480 336320 10542
rect 338672 5908 338724 5914
rect 338672 5850 338724 5856
rect 337476 2916 337528 2922
rect 337476 2858 337528 2864
rect 337488 480 337516 2858
rect 338684 480 338712 5850
rect 339868 4616 339920 4622
rect 339868 4558 339920 4564
rect 339880 480 339908 4558
rect 340972 3120 341024 3126
rect 340972 3062 341024 3068
rect 340984 480 341012 3062
rect 342180 480 342208 16526
rect 343364 5976 343416 5982
rect 343364 5918 343416 5924
rect 343376 480 343404 5918
rect 344560 2984 344612 2990
rect 344560 2926 344612 2932
rect 344572 480 344600 2926
rect 345308 490 345336 16546
rect 346952 6044 347004 6050
rect 346952 5986 347004 5992
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 5986
rect 348068 480 348096 16546
rect 349264 480 349292 16546
rect 354036 6792 354088 6798
rect 354036 6734 354088 6740
rect 350448 6112 350500 6118
rect 350448 6054 350500 6060
rect 350460 480 350488 6054
rect 352840 4684 352892 4690
rect 352840 4626 352892 4632
rect 351644 3052 351696 3058
rect 351644 2994 351696 3000
rect 351656 480 351684 2994
rect 352852 480 352880 4626
rect 354048 480 354076 6734
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357452 3126 357480 332250
rect 358832 16574 358860 332930
rect 359476 322250 359504 360266
rect 360856 322318 360884 361694
rect 361580 336592 361632 336598
rect 361580 336534 361632 336540
rect 360844 322312 360896 322318
rect 360844 322254 360896 322260
rect 359464 322244 359516 322250
rect 359464 322186 359516 322192
rect 361592 16574 361620 336534
rect 362960 333056 363012 333062
rect 362960 332998 363012 333004
rect 362972 16574 363000 332998
rect 363616 322182 363644 362986
rect 367744 362976 367796 362982
rect 367744 362918 367796 362924
rect 363604 322176 363656 322182
rect 363604 322118 363656 322124
rect 367756 322114 367784 362918
rect 368480 336524 368532 336530
rect 368480 336466 368532 336472
rect 367744 322108 367796 322114
rect 367744 322050 367796 322056
rect 364340 239964 364392 239970
rect 364340 239906 364392 239912
rect 364352 236162 364380 239906
rect 364340 236156 364392 236162
rect 364340 236098 364392 236104
rect 365720 80776 365772 80782
rect 365720 80718 365772 80724
rect 358832 16546 359504 16574
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 357532 6724 357584 6730
rect 357532 6666 357584 6672
rect 357440 3120 357492 3126
rect 357440 3062 357492 3068
rect 357544 480 357572 6666
rect 358728 3120 358780 3126
rect 358728 3062 358780 3068
rect 358740 480 358768 3062
rect 359476 490 359504 16546
rect 361120 6656 361172 6662
rect 361120 6598 361172 6604
rect 359752 598 359964 626
rect 359752 490 359780 598
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 462 359780 490
rect 359936 480 359964 598
rect 361132 480 361160 6598
rect 361868 490 361896 16546
rect 362144 598 362356 626
rect 362144 490 362172 598
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 361868 462 362172 490
rect 362328 480 362356 598
rect 363524 480 363552 16546
rect 364616 6588 364668 6594
rect 364616 6530 364668 6536
rect 364628 480 364656 6530
rect 365732 3126 365760 80718
rect 368492 16574 368520 336466
rect 370516 248402 370544 379510
rect 372620 336456 372672 336462
rect 372620 336398 372672 336404
rect 370504 248396 370556 248402
rect 370504 248338 370556 248344
rect 369860 84924 369912 84930
rect 369860 84866 369912 84872
rect 369872 16574 369900 84866
rect 372632 16574 372660 336398
rect 375380 336388 375432 336394
rect 375380 336330 375432 336336
rect 375392 16574 375420 336330
rect 382280 336320 382332 336326
rect 382280 336262 382332 336268
rect 380900 333124 380952 333130
rect 380900 333066 380952 333072
rect 380912 16574 380940 333066
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 372632 16546 372936 16574
rect 375392 16546 376064 16574
rect 380912 16546 381216 16574
rect 365812 8356 365864 8362
rect 365812 8298 365864 8304
rect 365720 3120 365772 3126
rect 365720 3062 365772 3068
rect 365824 480 365852 8298
rect 368204 6520 368256 6526
rect 368204 6462 368256 6468
rect 367008 3120 367060 3126
rect 367008 3062 367060 3068
rect 367020 480 367048 3062
rect 368216 480 368244 6462
rect 369412 480 369440 16546
rect 370148 490 370176 16546
rect 371240 10532 371292 10538
rect 371240 10474 371292 10480
rect 370424 598 370636 626
rect 370424 490 370452 598
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 462 370452 490
rect 370608 480 370636 598
rect 371252 490 371280 10474
rect 371528 598 371740 626
rect 371528 490 371556 598
rect 370566 -960 370678 480
rect 371252 462 371556 490
rect 371712 480 371740 598
rect 372908 480 372936 16546
rect 374000 10464 374052 10470
rect 374000 10406 374052 10412
rect 374012 3126 374040 10406
rect 374092 6452 374144 6458
rect 374092 6394 374144 6400
rect 374000 3120 374052 3126
rect 374000 3062 374052 3068
rect 374104 480 374132 6394
rect 375288 3120 375340 3126
rect 375288 3062 375340 3068
rect 375300 480 375328 3062
rect 376036 490 376064 16546
rect 378416 10396 378468 10402
rect 378416 10338 378468 10344
rect 377680 6384 377732 6390
rect 377680 6326 377732 6332
rect 376312 598 376524 626
rect 376312 490 376340 598
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 462 376340 490
rect 376496 480 376524 598
rect 377692 480 377720 6326
rect 378428 490 378456 10338
rect 379980 8424 380032 8430
rect 379980 8366 380032 8372
rect 378704 598 378916 626
rect 378704 490 378732 598
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 462 378732 490
rect 378888 480 378916 598
rect 379992 480 380020 8366
rect 381188 480 381216 16546
rect 382292 3126 382320 336262
rect 397460 336252 397512 336258
rect 397460 336194 397512 336200
rect 396724 335300 396776 335306
rect 396724 335242 396776 335248
rect 387800 334552 387852 334558
rect 387800 334494 387852 334500
rect 383660 333940 383712 333946
rect 383660 333882 383712 333888
rect 383672 16574 383700 333882
rect 385040 80708 385092 80714
rect 385040 80650 385092 80656
rect 385052 16574 385080 80650
rect 383672 16546 384344 16574
rect 385052 16546 386000 16574
rect 382372 10328 382424 10334
rect 382372 10270 382424 10276
rect 382280 3120 382332 3126
rect 382280 3062 382332 3068
rect 382384 480 382412 10270
rect 383568 3120 383620 3126
rect 383568 3062 383620 3068
rect 383580 480 383608 3062
rect 384316 490 384344 16546
rect 384592 598 384804 626
rect 384592 490 384620 598
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 462 384620 490
rect 384776 480 384804 598
rect 385972 480 386000 16546
rect 387156 8492 387208 8498
rect 387156 8434 387208 8440
rect 387168 480 387196 8434
rect 387812 490 387840 334494
rect 393964 334484 394016 334490
rect 393964 334426 394016 334432
rect 391204 334348 391256 334354
rect 391204 334290 391256 334296
rect 390652 333192 390704 333198
rect 390652 333134 390704 333140
rect 389180 87780 389232 87786
rect 389180 87722 389232 87728
rect 389192 16574 389220 87722
rect 390664 16574 390692 333134
rect 389192 16546 389496 16574
rect 390664 16546 391152 16574
rect 388088 598 388300 626
rect 388088 490 388116 598
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 462 388116 490
rect 388272 480 388300 598
rect 389468 480 389496 16546
rect 390652 3188 390704 3194
rect 390652 3130 390704 3136
rect 390664 480 390692 3130
rect 391124 2938 391152 16546
rect 391216 3058 391244 334290
rect 393044 6316 393096 6322
rect 393044 6258 393096 6264
rect 391204 3052 391256 3058
rect 391204 2994 391256 3000
rect 391124 2910 391888 2938
rect 391860 480 391888 2910
rect 393056 480 393084 6258
rect 393976 3194 394004 334426
rect 394700 333872 394752 333878
rect 394700 333814 394752 333820
rect 394712 16574 394740 333814
rect 394712 16546 395384 16574
rect 394240 3256 394292 3262
rect 394240 3198 394292 3204
rect 393964 3188 394016 3194
rect 393964 3130 394016 3136
rect 394252 480 394280 3198
rect 395356 480 395384 16546
rect 396540 6248 396592 6254
rect 396540 6190 396592 6196
rect 396552 480 396580 6190
rect 396736 3262 396764 335242
rect 397472 16574 397500 336194
rect 404360 336184 404412 336190
rect 404360 336126 404412 336132
rect 403624 335232 403676 335238
rect 403624 335174 403676 335180
rect 398840 333804 398892 333810
rect 398840 333746 398892 333752
rect 398852 16574 398880 333746
rect 400862 332208 400918 332217
rect 400862 332143 400918 332152
rect 397472 16546 397776 16574
rect 398852 16546 398972 16574
rect 396724 3256 396776 3262
rect 396724 3198 396776 3204
rect 397748 480 397776 16546
rect 398944 480 398972 16546
rect 400128 6180 400180 6186
rect 400128 6122 400180 6128
rect 400140 480 400168 6122
rect 400876 3126 400904 332143
rect 402980 177608 403032 177614
rect 402980 177550 403032 177556
rect 402992 16574 403020 177550
rect 402992 16546 403572 16574
rect 402520 8560 402572 8566
rect 402520 8502 402572 8508
rect 401324 3392 401376 3398
rect 401324 3334 401376 3340
rect 400864 3120 400916 3126
rect 400864 3062 400916 3068
rect 401336 480 401364 3334
rect 402532 480 402560 8502
rect 403544 3210 403572 16546
rect 403636 3398 403664 335174
rect 403624 3392 403676 3398
rect 403624 3334 403676 3340
rect 403544 3182 403664 3210
rect 403636 480 403664 3182
rect 404372 490 404400 336126
rect 411260 336116 411312 336122
rect 411260 336058 411312 336064
rect 405740 335096 405792 335102
rect 405740 335038 405792 335044
rect 405752 16574 405780 335038
rect 407762 334520 407818 334529
rect 407762 334455 407818 334464
rect 407212 87712 407264 87718
rect 407212 87654 407264 87660
rect 405752 16546 406056 16574
rect 404648 598 404860 626
rect 404648 490 404676 598
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 462 404676 490
rect 404832 480 404860 598
rect 406028 480 406056 16546
rect 407224 480 407252 87654
rect 407776 4026 407804 334455
rect 409142 333840 409198 333849
rect 409142 333775 409198 333784
rect 408500 333736 408552 333742
rect 408500 333678 408552 333684
rect 408512 6914 408540 333678
rect 409156 16574 409184 333775
rect 411272 16574 411300 336058
rect 418160 336048 418212 336054
rect 418160 335990 418212 335996
rect 414662 333704 414718 333713
rect 412640 333668 412692 333674
rect 414662 333639 414718 333648
rect 412640 333610 412692 333616
rect 409156 16546 409276 16574
rect 411272 16546 411944 16574
rect 408512 6886 409184 6914
rect 407776 3998 408540 4026
rect 408512 3874 408540 3998
rect 408408 3868 408460 3874
rect 408408 3810 408460 3816
rect 408500 3868 408552 3874
rect 408500 3810 408552 3816
rect 408420 480 408448 3810
rect 409156 490 409184 6886
rect 409248 2922 409276 16546
rect 410798 6488 410854 6497
rect 410798 6423 410854 6432
rect 409236 2916 409288 2922
rect 409236 2858 409288 2864
rect 409432 598 409644 626
rect 409432 490 409460 598
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 462 409460 490
rect 409616 480 409644 598
rect 410812 480 410840 6423
rect 411916 480 411944 16546
rect 412652 490 412680 333610
rect 414294 6352 414350 6361
rect 414294 6287 414350 6296
rect 412928 598 413140 626
rect 412928 490 412956 598
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 462 412956 490
rect 413112 480 413140 598
rect 414308 480 414336 6287
rect 414676 2854 414704 333639
rect 415400 333600 415452 333606
rect 415400 333542 415452 333548
rect 417422 333568 417478 333577
rect 415412 2990 415440 333542
rect 417422 333503 417478 333512
rect 416780 177540 416832 177546
rect 416780 177482 416832 177488
rect 415492 8628 415544 8634
rect 415492 8570 415544 8576
rect 415400 2984 415452 2990
rect 415400 2926 415452 2932
rect 414664 2848 414716 2854
rect 414664 2790 414716 2796
rect 415504 480 415532 8570
rect 416792 6914 416820 177482
rect 417436 16574 417464 333503
rect 418172 16574 418200 335990
rect 433984 335164 434036 335170
rect 433984 335106 434036 335112
rect 423680 333532 423732 333538
rect 423680 333474 423732 333480
rect 422944 330676 422996 330682
rect 422944 330618 422996 330624
rect 420920 89004 420972 89010
rect 420920 88946 420972 88952
rect 417436 16546 417556 16574
rect 418172 16546 418568 16574
rect 416792 6886 417464 6914
rect 416688 2984 416740 2990
rect 416688 2926 416740 2932
rect 416700 480 416728 2926
rect 417436 490 417464 6886
rect 417528 2990 417556 16546
rect 417516 2984 417568 2990
rect 417516 2926 417568 2932
rect 417712 598 417924 626
rect 417712 490 417740 598
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 462 417740 490
rect 417896 480 417924 598
rect 418540 490 418568 16546
rect 420184 8696 420236 8702
rect 420184 8638 420236 8644
rect 418816 598 419028 626
rect 418816 490 418844 598
rect 417854 -960 417966 480
rect 418540 462 418844 490
rect 419000 480 419028 598
rect 420196 480 420224 8638
rect 420932 490 420960 88946
rect 422956 4078 422984 330618
rect 423692 6914 423720 333474
rect 430580 333464 430632 333470
rect 430580 333406 430632 333412
rect 426440 333396 426492 333402
rect 426440 333338 426492 333344
rect 423772 332240 423824 332246
rect 423772 332182 423824 332188
rect 423784 11762 423812 332182
rect 426452 16574 426480 333338
rect 430592 16574 430620 333406
rect 433340 333328 433392 333334
rect 433340 333270 433392 333276
rect 433352 16574 433380 333270
rect 426452 16546 426848 16574
rect 430592 16546 430896 16574
rect 433352 16546 433932 16574
rect 423772 11756 423824 11762
rect 423772 11698 423824 11704
rect 424968 11756 425020 11762
rect 424968 11698 425020 11704
rect 423692 6886 423812 6914
rect 422576 4072 422628 4078
rect 422576 4014 422628 4020
rect 422944 4072 422996 4078
rect 422944 4014 422996 4020
rect 421208 598 421420 626
rect 421208 490 421236 598
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 462 421236 490
rect 421392 480 421420 598
rect 422588 480 422616 4014
rect 423784 480 423812 6886
rect 424980 480 425008 11698
rect 426164 3936 426216 3942
rect 426164 3878 426216 3884
rect 426176 480 426204 3878
rect 426820 490 426848 16546
rect 428462 6216 428518 6225
rect 428462 6151 428518 6160
rect 427096 598 427308 626
rect 427096 490 427124 598
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 462 427124 490
rect 427280 480 427308 598
rect 428476 480 428504 6151
rect 429660 4004 429712 4010
rect 429660 3946 429712 3952
rect 429672 480 429700 3946
rect 430868 480 430896 16546
rect 432052 6996 432104 7002
rect 432052 6938 432104 6944
rect 432064 480 432092 6938
rect 433248 4140 433300 4146
rect 433248 4082 433300 4088
rect 433260 480 433288 4082
rect 433904 626 433932 16546
rect 433996 4078 434024 335106
rect 434076 335028 434128 335034
rect 434076 334970 434128 334976
rect 433984 4072 434036 4078
rect 433984 4014 434036 4020
rect 434088 3942 434116 334970
rect 434168 334960 434220 334966
rect 434168 334902 434220 334908
rect 434180 4146 434208 334902
rect 437480 334892 437532 334898
rect 437480 334834 437532 334840
rect 436744 333260 436796 333266
rect 436744 333202 436796 333208
rect 436756 265713 436784 333202
rect 437020 332172 437072 332178
rect 437020 332114 437072 332120
rect 436928 332104 436980 332110
rect 436928 332046 436980 332052
rect 436836 332036 436888 332042
rect 436836 331978 436888 331984
rect 436848 267481 436876 331978
rect 436940 271998 436968 332046
rect 436928 271992 436980 271998
rect 436928 271934 436980 271940
rect 436928 271856 436980 271862
rect 436928 271798 436980 271804
rect 436940 271289 436968 271798
rect 436926 271280 436982 271289
rect 436926 271215 436982 271224
rect 437032 270065 437060 332114
rect 437112 327752 437164 327758
rect 437112 327694 437164 327700
rect 437124 273057 437152 327694
rect 437388 278792 437440 278798
rect 437388 278734 437440 278740
rect 437400 274145 437428 278734
rect 437386 274136 437442 274145
rect 437386 274071 437442 274080
rect 437110 273048 437166 273057
rect 437110 272983 437166 272992
rect 437112 271992 437164 271998
rect 437112 271934 437164 271940
rect 437018 270056 437074 270065
rect 437018 269991 437074 270000
rect 436928 269068 436980 269074
rect 436928 269010 436980 269016
rect 436940 268433 436968 269010
rect 436926 268424 436982 268433
rect 436926 268359 436982 268368
rect 436834 267472 436890 267481
rect 436834 267407 436890 267416
rect 436848 266830 436876 267407
rect 436836 266824 436888 266830
rect 436836 266766 436888 266772
rect 436742 265704 436798 265713
rect 436742 265639 436798 265648
rect 436756 258074 436784 265639
rect 436940 262970 436968 268359
rect 437032 267734 437060 269991
rect 437124 269074 437152 271934
rect 437112 269068 437164 269074
rect 437112 269010 437164 269016
rect 437032 267706 437336 267734
rect 437204 266824 437256 266830
rect 437204 266766 437256 266772
rect 436940 262942 437152 262970
rect 436756 258046 437060 258074
rect 436100 248396 436152 248402
rect 436100 248338 436152 248344
rect 436112 247353 436140 248338
rect 436098 247344 436154 247353
rect 436098 247279 436154 247288
rect 436100 245608 436152 245614
rect 436098 245576 436100 245585
rect 436152 245576 436154 245585
rect 436098 245511 436154 245520
rect 437032 239358 437060 258046
rect 437124 239970 437152 262942
rect 437112 239964 437164 239970
rect 437112 239906 437164 239912
rect 437020 239352 437072 239358
rect 437020 239294 437072 239300
rect 437216 237697 437244 266766
rect 437308 240038 437336 267706
rect 437296 240032 437348 240038
rect 437296 239974 437348 239980
rect 437400 239766 437428 274071
rect 437388 239760 437440 239766
rect 437388 239702 437440 239708
rect 437202 237688 437258 237697
rect 437202 237623 437258 237632
rect 434720 177472 434772 177478
rect 434720 177414 434772 177420
rect 434732 16574 434760 177414
rect 434732 16546 435128 16574
rect 434168 4140 434220 4146
rect 434168 4082 434220 4088
rect 434076 3936 434128 3942
rect 434076 3878 434128 3884
rect 433904 598 434024 626
rect 433996 490 434024 598
rect 434272 598 434484 626
rect 434272 490 434300 598
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 462 434300 490
rect 434456 480 434484 598
rect 435100 490 435128 16546
rect 436744 3324 436796 3330
rect 436744 3266 436796 3272
rect 435376 598 435588 626
rect 435376 490 435404 598
rect 434414 -960 434526 480
rect 435100 462 435404 490
rect 435560 480 435588 598
rect 436756 480 436784 3266
rect 437492 490 437520 334834
rect 438136 237454 438164 385018
rect 537116 380928 537168 380934
rect 537116 380870 537168 380876
rect 453304 372768 453356 372774
rect 453304 372710 453356 372716
rect 450544 371272 450596 371278
rect 450544 371214 450596 371220
rect 440976 367192 441028 367198
rect 440976 367134 441028 367140
rect 440884 367124 440936 367130
rect 440884 367066 440936 367072
rect 438216 354748 438268 354754
rect 438216 354690 438268 354696
rect 438228 237590 438256 354690
rect 439688 350600 439740 350606
rect 439688 350542 439740 350548
rect 439504 337000 439556 337006
rect 439504 336942 439556 336948
rect 438766 273048 438822 273057
rect 438766 272983 438822 272992
rect 438674 271280 438730 271289
rect 438674 271215 438730 271224
rect 438584 240100 438636 240106
rect 438584 240042 438636 240048
rect 438216 237584 438268 237590
rect 438216 237526 438268 237532
rect 438124 237448 438176 237454
rect 438124 237390 438176 237396
rect 438596 237386 438624 240042
rect 438688 239222 438716 271215
rect 438780 239290 438808 272983
rect 439412 240780 439464 240786
rect 439412 240722 439464 240728
rect 438768 239284 438820 239290
rect 438768 239226 438820 239232
rect 438676 239216 438728 239222
rect 438676 239158 438728 239164
rect 438584 237380 438636 237386
rect 438584 237322 438636 237328
rect 439424 236609 439452 240722
rect 439410 236600 439466 236609
rect 439410 236535 439466 236544
rect 439516 4010 439544 336942
rect 439594 333432 439650 333441
rect 439594 333367 439650 333376
rect 439136 4004 439188 4010
rect 439136 3946 439188 3952
rect 439504 4004 439556 4010
rect 439504 3946 439556 3952
rect 437768 598 437980 626
rect 437768 490 437796 598
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437492 462 437796 490
rect 437952 480 437980 598
rect 439148 480 439176 3946
rect 439608 3330 439636 333367
rect 439700 237522 439728 350542
rect 439780 338156 439832 338162
rect 439780 338098 439832 338104
rect 439792 239834 439820 338098
rect 440896 322046 440924 367066
rect 440884 322040 440936 322046
rect 440884 321982 440936 321988
rect 440988 321978 441016 367134
rect 449164 358828 449216 358834
rect 449164 358770 449216 358776
rect 449176 322930 449204 358770
rect 449164 322924 449216 322930
rect 449164 322866 449216 322872
rect 440976 321972 441028 321978
rect 440976 321914 441028 321920
rect 450556 321910 450584 371214
rect 450544 321904 450596 321910
rect 450544 321846 450596 321852
rect 453316 321774 453344 372710
rect 454684 372700 454736 372706
rect 454684 372642 454736 372648
rect 454696 321842 454724 372642
rect 496820 372632 496872 372638
rect 496820 372574 496872 372580
rect 488540 369980 488592 369986
rect 488540 369922 488592 369928
rect 485044 368620 485096 368626
rect 485044 368562 485096 368568
rect 478880 364404 478932 364410
rect 478880 364346 478932 364352
rect 472072 361684 472124 361690
rect 472072 361626 472124 361632
rect 470600 360256 470652 360262
rect 470600 360198 470652 360204
rect 467840 358352 467892 358358
rect 467840 358294 467892 358300
rect 467852 322561 467880 358294
rect 469404 322924 469456 322930
rect 469404 322866 469456 322872
rect 467838 322552 467894 322561
rect 467838 322487 467894 322496
rect 454684 321836 454736 321842
rect 454684 321778 454736 321784
rect 453304 321768 453356 321774
rect 453304 321710 453356 321716
rect 469416 321609 469444 322866
rect 470612 322833 470640 360198
rect 470598 322824 470654 322833
rect 470598 322759 470654 322768
rect 470506 322688 470562 322697
rect 470506 322623 470562 322632
rect 469402 321600 469458 321609
rect 469402 321535 469458 321544
rect 470520 319977 470548 322623
rect 472084 322561 472112 361626
rect 474740 361616 474792 361622
rect 474740 361558 474792 361564
rect 474752 322561 474780 361558
rect 478892 322561 478920 364346
rect 480260 358284 480312 358290
rect 480260 358226 480312 358232
rect 480272 322561 480300 358226
rect 481640 358216 481692 358222
rect 481640 358158 481692 358164
rect 481652 322561 481680 358158
rect 483020 358148 483072 358154
rect 483020 358090 483072 358096
rect 483032 322561 483060 358090
rect 485056 322930 485084 368562
rect 486424 368552 486476 368558
rect 486424 368494 486476 368500
rect 485044 322924 485096 322930
rect 485044 322866 485096 322872
rect 486332 322924 486384 322930
rect 486332 322866 486384 322872
rect 486344 322561 486372 322866
rect 472070 322552 472126 322561
rect 472070 322487 472126 322496
rect 474738 322552 474794 322561
rect 474738 322487 474794 322496
rect 478878 322552 478934 322561
rect 478878 322487 478934 322496
rect 480258 322552 480314 322561
rect 480258 322487 480314 322496
rect 481638 322552 481694 322561
rect 481638 322487 481694 322496
rect 483018 322552 483074 322561
rect 483018 322487 483074 322496
rect 486330 322552 486386 322561
rect 486330 322487 486386 322496
rect 474556 322312 474608 322318
rect 474556 322254 474608 322260
rect 471980 322244 472032 322250
rect 471980 322186 472032 322192
rect 471992 321609 472020 322186
rect 474568 321609 474596 322254
rect 476764 322176 476816 322182
rect 476764 322118 476816 322124
rect 476776 321609 476804 322118
rect 478236 322108 478288 322114
rect 478236 322050 478288 322056
rect 478248 321609 478276 322050
rect 485412 322040 485464 322046
rect 485412 321982 485464 321988
rect 484400 321972 484452 321978
rect 484400 321914 484452 321920
rect 484412 321609 484440 321914
rect 485424 321609 485452 321982
rect 486436 321638 486464 368494
rect 488552 322561 488580 369922
rect 489920 369912 489972 369918
rect 489920 369854 489972 369860
rect 489932 322561 489960 369854
rect 491300 358080 491352 358086
rect 491300 358022 491352 358028
rect 491312 322561 491340 358022
rect 496832 322561 496860 372574
rect 536840 334824 536892 334830
rect 536840 334766 536892 334772
rect 519544 331968 519596 331974
rect 519544 331910 519596 331916
rect 498200 322856 498252 322862
rect 498200 322798 498252 322804
rect 488538 322552 488594 322561
rect 488538 322487 488594 322496
rect 489918 322552 489974 322561
rect 489918 322487 489974 322496
rect 491298 322552 491354 322561
rect 491298 322487 491354 322496
rect 496818 322552 496874 322561
rect 496818 322487 496874 322496
rect 492772 321904 492824 321910
rect 492772 321846 492824 321852
rect 486424 321632 486476 321638
rect 471978 321600 472034 321609
rect 471978 321535 472034 321544
rect 474554 321600 474610 321609
rect 474554 321535 474610 321544
rect 476762 321600 476818 321609
rect 476762 321535 476818 321544
rect 478234 321600 478290 321609
rect 478234 321535 478290 321544
rect 484398 321600 484454 321609
rect 484398 321535 484454 321544
rect 485410 321600 485466 321609
rect 488172 321632 488224 321638
rect 486424 321574 486476 321580
rect 488170 321600 488172 321609
rect 492784 321609 492812 321846
rect 495532 321836 495584 321842
rect 495532 321778 495584 321784
rect 494244 321768 494296 321774
rect 494244 321710 494296 321716
rect 494256 321609 494284 321710
rect 495544 321609 495572 321778
rect 498212 321609 498240 322798
rect 499212 322788 499264 322794
rect 499212 322730 499264 322736
rect 499224 321609 499252 322730
rect 500684 322720 500736 322726
rect 500684 322662 500736 322668
rect 500696 321609 500724 322662
rect 501236 322652 501288 322658
rect 501236 322594 501288 322600
rect 501248 321609 501276 322594
rect 503260 322584 503312 322590
rect 503260 322526 503312 322532
rect 503272 321609 503300 322526
rect 505468 322516 505520 322522
rect 505468 322458 505520 322464
rect 503812 322448 503864 322454
rect 503812 322390 503864 322396
rect 503824 321609 503852 322390
rect 505480 321609 505508 322458
rect 519556 322425 519584 331910
rect 519542 322416 519598 322425
rect 506940 322380 506992 322386
rect 519542 322351 519598 322360
rect 506940 322322 506992 322328
rect 506952 321609 506980 322322
rect 519556 322250 519584 322351
rect 519544 322244 519596 322250
rect 519544 322186 519596 322192
rect 530032 321632 530084 321638
rect 488224 321600 488226 321609
rect 485410 321535 485466 321544
rect 488170 321535 488226 321544
rect 492770 321600 492826 321609
rect 492770 321535 492826 321544
rect 494242 321600 494298 321609
rect 494242 321535 494298 321544
rect 495530 321600 495586 321609
rect 495530 321535 495586 321544
rect 498198 321600 498254 321609
rect 498198 321535 498254 321544
rect 499210 321600 499266 321609
rect 499210 321535 499266 321544
rect 500682 321600 500738 321609
rect 500682 321535 500738 321544
rect 501234 321600 501290 321609
rect 501234 321535 501290 321544
rect 503258 321600 503314 321609
rect 503258 321535 503314 321544
rect 503810 321600 503866 321609
rect 503810 321535 503866 321544
rect 505466 321600 505522 321609
rect 505466 321535 505522 321544
rect 506938 321600 506994 321609
rect 506938 321535 506994 321544
rect 530030 321600 530032 321609
rect 530084 321600 530086 321609
rect 530030 321535 530086 321544
rect 470506 319968 470562 319977
rect 470506 319903 470562 319912
rect 439872 240032 439924 240038
rect 439872 239974 439924 239980
rect 439780 239828 439832 239834
rect 439780 239770 439832 239776
rect 439884 239306 439912 239974
rect 441436 239896 441488 239902
rect 502338 239864 502394 239873
rect 441488 239844 441660 239850
rect 441436 239838 441660 239844
rect 441448 239822 441660 239838
rect 439884 239278 441568 239306
rect 441540 239222 441568 239278
rect 441528 239216 441580 239222
rect 441528 239158 441580 239164
rect 439688 237516 439740 237522
rect 439688 237458 439740 237464
rect 440240 235408 440292 235414
rect 440240 235350 440292 235356
rect 440252 4214 440280 235350
rect 441632 16574 441660 239822
rect 467840 239828 467892 239834
rect 502338 239799 502394 239808
rect 523130 239864 523186 239873
rect 523130 239799 523186 239808
rect 467840 239770 467892 239776
rect 459560 239692 459612 239698
rect 459560 239634 459612 239640
rect 452106 239184 452162 239193
rect 446404 239148 446456 239154
rect 446404 239090 446456 239096
rect 447048 239148 447100 239154
rect 452106 239119 452162 239128
rect 447048 239090 447100 239096
rect 446416 236473 446444 239090
rect 447060 237289 447088 239090
rect 451646 238912 451702 238921
rect 451646 238847 451702 238856
rect 451660 238626 451688 238847
rect 452120 238785 452148 239119
rect 456798 239048 456854 239057
rect 456798 238983 456854 238992
rect 456812 238898 456840 238983
rect 457074 238912 457130 238921
rect 456812 238870 457074 238898
rect 457074 238847 457130 238856
rect 452106 238776 452162 238785
rect 452290 238776 452346 238785
rect 452106 238711 452162 238720
rect 452212 238734 452290 238762
rect 452212 238626 452240 238734
rect 452290 238711 452346 238720
rect 451660 238598 452240 238626
rect 459572 237561 459600 239634
rect 465172 239624 465224 239630
rect 465172 239566 465224 239572
rect 465080 238128 465132 238134
rect 465080 238070 465132 238076
rect 465092 237969 465120 238070
rect 461582 237960 461638 237969
rect 461582 237895 461638 237904
rect 463698 237960 463754 237969
rect 463698 237895 463754 237904
rect 465078 237960 465134 237969
rect 465078 237895 465134 237904
rect 459558 237552 459614 237561
rect 459558 237487 459614 237496
rect 447046 237280 447102 237289
rect 447046 237215 447102 237224
rect 460938 237280 460994 237289
rect 460938 237215 460994 237224
rect 446402 236464 446458 236473
rect 446402 236399 446458 236408
rect 460952 236230 460980 237215
rect 461596 236230 461624 237895
rect 463712 237726 463740 237895
rect 463700 237720 463752 237726
rect 463700 237662 463752 237668
rect 460940 236224 460992 236230
rect 460940 236166 460992 236172
rect 461584 236224 461636 236230
rect 461584 236166 461636 236172
rect 462320 236088 462372 236094
rect 462320 236030 462372 236036
rect 462410 236056 462466 236065
rect 445760 235340 445812 235346
rect 445760 235282 445812 235288
rect 444380 162172 444432 162178
rect 444380 162114 444432 162120
rect 444392 16574 444420 162114
rect 441632 16546 442672 16574
rect 444392 16546 445064 16574
rect 440332 8764 440384 8770
rect 440332 8706 440384 8712
rect 440240 4208 440292 4214
rect 440240 4150 440292 4156
rect 439596 3324 439648 3330
rect 439596 3266 439648 3272
rect 440344 480 440372 8706
rect 441528 4208 441580 4214
rect 441528 4150 441580 4156
rect 441540 480 441568 4150
rect 442644 480 442672 16546
rect 443828 3732 443880 3738
rect 443828 3674 443880 3680
rect 443840 480 443868 3674
rect 445036 480 445064 16546
rect 445772 490 445800 235282
rect 456800 87644 456852 87650
rect 456800 87586 456852 87592
rect 452660 84856 452712 84862
rect 452660 84798 452712 84804
rect 448612 82136 448664 82142
rect 448612 82078 448664 82084
rect 448624 13326 448652 82078
rect 452672 16574 452700 84798
rect 456812 16574 456840 87586
rect 452672 16546 453344 16574
rect 456812 16546 456932 16574
rect 448612 13320 448664 13326
rect 448612 13262 448664 13268
rect 449808 13320 449860 13326
rect 449808 13262 449860 13268
rect 447416 3800 447468 3806
rect 447416 3742 447468 3748
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 3742
rect 448612 3324 448664 3330
rect 448612 3266 448664 3272
rect 448624 480 448652 3266
rect 449820 480 449848 13262
rect 452108 8900 452160 8906
rect 452108 8842 452160 8848
rect 450912 8832 450964 8838
rect 450912 8774 450964 8780
rect 450924 480 450952 8774
rect 452120 480 452148 8842
rect 453316 480 453344 16546
rect 454500 3664 454552 3670
rect 454500 3606 454552 3612
rect 454512 480 454540 3606
rect 455696 2916 455748 2922
rect 455696 2858 455748 2864
rect 455708 480 455736 2858
rect 456904 480 456932 16546
rect 460388 7064 460440 7070
rect 460388 7006 460440 7012
rect 458088 4752 458140 4758
rect 458088 4694 458140 4700
rect 458100 480 458128 4694
rect 459192 2848 459244 2854
rect 459192 2790 459244 2796
rect 459204 480 459232 2790
rect 460400 480 460428 7006
rect 461584 3596 461636 3602
rect 461584 3538 461636 3544
rect 461596 480 461624 3538
rect 462332 490 462360 236030
rect 462410 235991 462412 236000
rect 462464 235991 462466 236000
rect 462412 235962 462464 235968
rect 465184 219434 465212 239566
rect 467852 239193 467880 239770
rect 472072 239760 472124 239766
rect 472072 239702 472124 239708
rect 467838 239184 467894 239193
rect 467838 239119 467894 239128
rect 469218 239184 469274 239193
rect 469218 239119 469274 239128
rect 469232 239086 469260 239119
rect 469220 239080 469272 239086
rect 469220 239022 469272 239028
rect 470690 238096 470746 238105
rect 468300 238060 468352 238066
rect 470690 238031 470746 238040
rect 471794 238096 471850 238105
rect 471794 238031 471850 238040
rect 468300 238002 468352 238008
rect 468312 237969 468340 238002
rect 467194 237960 467250 237969
rect 467194 237895 467250 237904
rect 468298 237960 468354 237969
rect 468298 237895 468354 237904
rect 467208 237862 467236 237895
rect 467196 237856 467248 237862
rect 467196 237798 467248 237804
rect 470704 237794 470732 238031
rect 471808 237930 471836 238031
rect 471796 237924 471848 237930
rect 471796 237866 471848 237872
rect 470692 237788 470744 237794
rect 470692 237730 470744 237736
rect 472084 237386 472112 239702
rect 473360 239556 473412 239562
rect 473360 239498 473412 239504
rect 471980 237380 472032 237386
rect 471980 237322 472032 237328
rect 472072 237380 472124 237386
rect 472072 237322 472124 237328
rect 471992 237289 472020 237322
rect 469218 237280 469274 237289
rect 469218 237215 469274 237224
rect 471978 237280 472034 237289
rect 471978 237215 472034 237224
rect 469232 235754 469260 237215
rect 472070 236600 472126 236609
rect 472070 236535 472126 236544
rect 472084 236366 472112 236535
rect 472072 236360 472124 236366
rect 471978 236328 472034 236337
rect 472072 236302 472124 236308
rect 471978 236263 471980 236272
rect 472032 236263 472034 236272
rect 471980 236234 472032 236240
rect 469220 235748 469272 235754
rect 469220 235690 469272 235696
rect 465092 219406 465212 219434
rect 465092 16574 465120 219406
rect 470600 79348 470652 79354
rect 470600 79290 470652 79296
rect 465092 16546 465856 16574
rect 463976 7132 464028 7138
rect 463976 7074 464028 7080
rect 462608 598 462820 626
rect 462608 490 462636 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462332 462 462636 490
rect 462792 480 462820 598
rect 463988 480 464016 7074
rect 465172 5500 465224 5506
rect 465172 5442 465224 5448
rect 465184 480 465212 5442
rect 465828 490 465856 16546
rect 467472 7200 467524 7206
rect 467472 7142 467524 7148
rect 466104 598 466316 626
rect 466104 490 466132 598
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 462 466132 490
rect 466288 480 466316 598
rect 467484 480 467512 7142
rect 468668 3528 468720 3534
rect 468668 3470 468720 3476
rect 468680 480 468708 3470
rect 469864 2984 469916 2990
rect 469864 2926 469916 2932
rect 469876 480 469904 2926
rect 470612 490 470640 79290
rect 473372 16574 473400 239498
rect 476120 239488 476172 239494
rect 476120 239430 476172 239436
rect 475658 238096 475714 238105
rect 475658 238031 475714 238040
rect 475672 237998 475700 238031
rect 475660 237992 475712 237998
rect 475660 237934 475712 237940
rect 473450 236600 473506 236609
rect 473450 236535 473506 236544
rect 473464 236434 473492 236535
rect 473452 236428 473504 236434
rect 473452 236370 473504 236376
rect 476132 16574 476160 239430
rect 481732 239420 481784 239426
rect 481732 239362 481784 239368
rect 480442 239048 480498 239057
rect 480442 238983 480498 238992
rect 480456 238950 480484 238983
rect 480444 238944 480496 238950
rect 479154 238912 479210 238921
rect 480444 238886 480496 238892
rect 479154 238847 479156 238856
rect 479208 238847 479210 238856
rect 479156 238818 479208 238824
rect 476762 238776 476818 238785
rect 476762 238711 476764 238720
rect 476816 238711 476818 238720
rect 477590 238776 477646 238785
rect 477590 238711 477646 238720
rect 476764 238682 476816 238688
rect 477498 236600 477554 236609
rect 477498 236535 477554 236544
rect 477512 236502 477540 236535
rect 477500 236496 477552 236502
rect 477500 236438 477552 236444
rect 477604 236162 477632 238711
rect 481640 237652 481692 237658
rect 481640 237594 481692 237600
rect 481652 237289 481680 237594
rect 481638 237280 481694 237289
rect 481638 237215 481694 237224
rect 480258 236736 480314 236745
rect 480258 236671 480314 236680
rect 480272 236638 480300 236671
rect 480260 236632 480312 236638
rect 480260 236574 480312 236580
rect 480534 236600 480590 236609
rect 480534 236535 480536 236544
rect 480588 236535 480590 236544
rect 480536 236506 480588 236512
rect 477592 236156 477644 236162
rect 477592 236098 477644 236104
rect 481744 219434 481772 239362
rect 484582 239320 484638 239329
rect 484582 239255 484638 239264
rect 483018 239048 483074 239057
rect 483018 238983 483020 238992
rect 483072 238983 483074 238992
rect 483020 238954 483072 238960
rect 483662 238504 483718 238513
rect 483662 238439 483718 238448
rect 483676 238105 483704 238439
rect 483662 238096 483718 238105
rect 483662 238031 483718 238040
rect 481916 237448 481968 237454
rect 481916 237390 481968 237396
rect 481928 237289 481956 237390
rect 481914 237280 481970 237289
rect 481914 237215 481970 237224
rect 483018 237144 483074 237153
rect 483018 237079 483074 237088
rect 483032 236978 483060 237079
rect 483020 236972 483072 236978
rect 483020 236914 483072 236920
rect 484398 236872 484454 236881
rect 484398 236807 484454 236816
rect 484412 236774 484440 236807
rect 484400 236768 484452 236774
rect 484400 236710 484452 236716
rect 481652 219406 481772 219434
rect 481652 16574 481680 219406
rect 484596 16574 484624 239255
rect 494242 238912 494298 238921
rect 494242 238847 494298 238856
rect 494256 238814 494284 238847
rect 494244 238808 494296 238814
rect 494244 238750 494296 238756
rect 487804 238672 487856 238678
rect 487804 238614 487856 238620
rect 490562 238640 490618 238649
rect 485412 238536 485464 238542
rect 484858 238504 484914 238513
rect 484858 238439 484860 238448
rect 484912 238439 484914 238448
rect 485410 238504 485412 238513
rect 487816 238513 487844 238614
rect 490562 238575 490564 238584
rect 490616 238575 490618 238584
rect 490564 238546 490616 238552
rect 485464 238504 485466 238513
rect 485410 238439 485466 238448
rect 487802 238504 487858 238513
rect 487802 238439 487858 238448
rect 491666 238504 491722 238513
rect 491666 238439 491722 238448
rect 484860 238410 484912 238416
rect 491680 238406 491708 238439
rect 491668 238400 491720 238406
rect 491668 238342 491720 238348
rect 492770 238368 492826 238377
rect 492770 238303 492772 238312
rect 492824 238303 492826 238312
rect 496818 238368 496874 238377
rect 496818 238303 496874 238312
rect 492772 238274 492824 238280
rect 496832 238270 496860 238303
rect 496820 238264 496872 238270
rect 496820 238206 496872 238212
rect 499210 238232 499266 238241
rect 499210 238167 499212 238176
rect 499264 238167 499266 238176
rect 499212 238138 499264 238144
rect 500960 237584 501012 237590
rect 500960 237526 501012 237532
rect 492680 237516 492732 237522
rect 492680 237458 492732 237464
rect 492692 237289 492720 237458
rect 495440 237312 495492 237318
rect 487158 237280 487214 237289
rect 487158 237215 487214 237224
rect 492678 237280 492734 237289
rect 492678 237215 492734 237224
rect 493322 237280 493378 237289
rect 493322 237215 493324 237224
rect 487172 237182 487200 237215
rect 493376 237215 493378 237224
rect 495438 237280 495440 237289
rect 500972 237289 501000 237526
rect 495492 237280 495494 237289
rect 495438 237215 495494 237224
rect 500958 237280 501014 237289
rect 500958 237215 501014 237224
rect 493324 237186 493376 237192
rect 487160 237176 487212 237182
rect 487160 237118 487212 237124
rect 488538 237144 488594 237153
rect 488538 237079 488594 237088
rect 496818 237144 496874 237153
rect 496818 237079 496820 237088
rect 488552 236910 488580 237079
rect 496872 237079 496874 237088
rect 499854 237144 499910 237153
rect 499854 237079 499910 237088
rect 496820 237050 496872 237056
rect 499868 237046 499896 237079
rect 499856 237040 499908 237046
rect 499856 236982 499908 236988
rect 488540 236904 488592 236910
rect 488540 236846 488592 236852
rect 491298 236872 491354 236881
rect 491298 236807 491300 236816
rect 491352 236807 491354 236816
rect 491300 236778 491352 236784
rect 485778 236736 485834 236745
rect 485778 236671 485780 236680
rect 485832 236671 485834 236680
rect 485780 236642 485832 236648
rect 485778 236464 485834 236473
rect 485778 236399 485834 236408
rect 485792 236230 485820 236399
rect 485780 236224 485832 236230
rect 485780 236166 485832 236172
rect 488540 83632 488592 83638
rect 488540 83574 488592 83580
rect 488552 16574 488580 83574
rect 502352 16574 502380 239799
rect 520278 239728 520334 239737
rect 520278 239663 520334 239672
rect 503718 236736 503774 236745
rect 503718 236671 503774 236680
rect 502430 236056 502486 236065
rect 502430 235991 502486 236000
rect 502444 235822 502472 235991
rect 503732 235890 503760 236671
rect 505098 236328 505154 236337
rect 505098 236263 505154 236272
rect 505112 235958 505140 236263
rect 505100 235952 505152 235958
rect 505100 235894 505152 235900
rect 503720 235884 503772 235890
rect 503720 235826 503772 235832
rect 502432 235816 502484 235822
rect 502432 235758 502484 235764
rect 505100 235272 505152 235278
rect 505100 235214 505152 235220
rect 505112 16574 505140 235214
rect 506480 83564 506532 83570
rect 506480 83506 506532 83512
rect 473372 16546 473492 16574
rect 476132 16546 476528 16574
rect 481652 16546 481772 16574
rect 484596 16546 484808 16574
rect 488552 16546 488856 16574
rect 502352 16546 503024 16574
rect 505112 16546 505416 16574
rect 472254 3768 472310 3777
rect 472254 3703 472310 3712
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 3703
rect 473464 480 473492 16546
rect 474556 7268 474608 7274
rect 474556 7210 474608 7216
rect 474568 480 474596 7210
rect 475752 5432 475804 5438
rect 475752 5374 475804 5380
rect 475764 480 475792 5374
rect 476500 490 476528 16546
rect 480536 9648 480588 9654
rect 480536 9590 480588 9596
rect 478144 7336 478196 7342
rect 478144 7278 478196 7284
rect 476776 598 476988 626
rect 476776 490 476804 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 462 476804 490
rect 476960 480 476988 598
rect 478156 480 478184 7278
rect 479338 3632 479394 3641
rect 479338 3567 479394 3576
rect 479352 480 479380 3567
rect 480548 480 480576 9590
rect 481744 480 481772 16546
rect 482836 7404 482888 7410
rect 482836 7346 482888 7352
rect 482848 480 482876 7346
rect 484030 3496 484086 3505
rect 484030 3431 484086 3440
rect 484044 480 484072 3431
rect 484780 490 484808 16546
rect 487620 9580 487672 9586
rect 487620 9522 487672 9528
rect 486424 7472 486476 7478
rect 486424 7414 486476 7420
rect 485056 598 485268 626
rect 485056 490 485084 598
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 462 485084 490
rect 485240 480 485268 598
rect 486436 480 486464 7414
rect 487632 480 487660 9522
rect 488828 480 488856 16546
rect 493508 8288 493560 8294
rect 493508 8230 493560 8236
rect 489920 7540 489972 7546
rect 489920 7482 489972 7488
rect 489932 480 489960 7482
rect 492312 5364 492364 5370
rect 492312 5306 492364 5312
rect 491116 3052 491168 3058
rect 491116 2994 491168 3000
rect 491128 480 491156 2994
rect 492324 480 492352 5306
rect 493520 480 493548 8230
rect 497096 8220 497148 8226
rect 497096 8162 497148 8168
rect 495900 5296 495952 5302
rect 495900 5238 495952 5244
rect 494704 3188 494756 3194
rect 494704 3130 494756 3136
rect 494716 480 494744 3130
rect 495912 480 495940 5238
rect 497108 480 497136 8162
rect 500592 8152 500644 8158
rect 500592 8094 500644 8100
rect 499396 5228 499448 5234
rect 499396 5170 499448 5176
rect 498200 3256 498252 3262
rect 498200 3198 498252 3204
rect 498212 480 498240 3198
rect 499408 480 499436 5170
rect 500604 480 500632 8094
rect 501788 3120 501840 3126
rect 501788 3062 501840 3068
rect 501800 480 501828 3062
rect 502996 480 503024 16546
rect 504180 8084 504232 8090
rect 504180 8026 504232 8032
rect 504192 480 504220 8026
rect 505388 480 505416 16546
rect 506492 480 506520 83506
rect 507676 8016 507728 8022
rect 507676 7958 507728 7964
rect 507688 480 507716 7958
rect 511264 7948 511316 7954
rect 511264 7890 511316 7896
rect 510068 5160 510120 5166
rect 510068 5102 510120 5108
rect 508872 4140 508924 4146
rect 508872 4082 508924 4088
rect 508884 480 508912 4082
rect 510080 480 510108 5102
rect 511276 480 511304 7890
rect 514760 7880 514812 7886
rect 514760 7822 514812 7828
rect 513564 5092 513616 5098
rect 513564 5034 513616 5040
rect 512460 4072 512512 4078
rect 512460 4014 512512 4020
rect 512472 480 512500 4014
rect 513576 480 513604 5034
rect 514772 480 514800 7822
rect 518348 7812 518400 7818
rect 518348 7754 518400 7760
rect 517152 5024 517204 5030
rect 517152 4966 517204 4972
rect 515956 3936 516008 3942
rect 515956 3878 516008 3884
rect 515968 480 515996 3878
rect 517164 480 517192 4966
rect 518360 480 518388 7754
rect 519544 4004 519596 4010
rect 519544 3946 519596 3952
rect 519556 480 519584 3946
rect 520292 490 520320 239663
rect 522670 239592 522726 239601
rect 522670 239527 522726 239536
rect 522854 239592 522910 239601
rect 522854 239527 522910 239536
rect 522684 239290 522712 239527
rect 522868 239358 522896 239527
rect 522856 239352 522908 239358
rect 522856 239294 522908 239300
rect 522672 239284 522724 239290
rect 522672 239226 522724 239232
rect 523144 239222 523172 239799
rect 523222 239456 523278 239465
rect 523222 239391 523278 239400
rect 523132 239216 523184 239222
rect 523132 239158 523184 239164
rect 523040 237380 523092 237386
rect 523040 237322 523092 237328
rect 523052 237289 523080 237322
rect 523038 237280 523094 237289
rect 523038 237215 523094 237224
rect 523236 16574 523264 239391
rect 527178 239320 527234 239329
rect 527178 239255 527234 239264
rect 527192 16574 527220 239255
rect 531320 83496 531372 83502
rect 531320 83438 531372 83444
rect 523236 16546 523816 16574
rect 527192 16546 527864 16574
rect 523040 9512 523092 9518
rect 523040 9454 523092 9460
rect 521844 7744 521896 7750
rect 521844 7686 521896 7692
rect 520568 598 520780 626
rect 520568 490 520596 598
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 462 520596 490
rect 520752 480 520780 598
rect 521856 480 521884 7686
rect 523052 480 523080 9454
rect 523788 490 523816 16546
rect 525432 7676 525484 7682
rect 525432 7618 525484 7624
rect 524064 598 524276 626
rect 524064 490 524092 598
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523788 462 524092 490
rect 524248 480 524276 598
rect 525444 480 525472 7618
rect 526628 3392 526680 3398
rect 526628 3334 526680 3340
rect 526640 480 526668 3334
rect 527836 480 527864 16546
rect 530124 9444 530176 9450
rect 530124 9386 530176 9392
rect 529020 7608 529072 7614
rect 529020 7550 529072 7556
rect 529032 480 529060 7550
rect 530136 480 530164 9386
rect 531332 480 531360 83438
rect 536852 16574 536880 334766
rect 536932 322244 536984 322250
rect 536932 322186 536984 322192
rect 536944 239698 536972 322186
rect 537024 321632 537076 321638
rect 537024 321574 537076 321580
rect 536932 239692 536984 239698
rect 536932 239634 536984 239640
rect 537036 239154 537064 321574
rect 537128 316577 537156 380870
rect 537114 316568 537170 316577
rect 537114 316503 537170 316512
rect 537496 259418 537524 390322
rect 537576 389292 537628 389298
rect 537576 389234 537628 389240
rect 537588 273222 537616 389234
rect 580354 389192 580410 389201
rect 580354 389127 580410 389136
rect 580172 388272 580224 388278
rect 580172 388214 580224 388220
rect 580184 378457 580212 388214
rect 580264 386436 580316 386442
rect 580264 386378 580316 386384
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 568580 336932 568632 336938
rect 568580 336874 568632 336880
rect 543738 335336 543794 335345
rect 543738 335271 543794 335280
rect 539600 334756 539652 334762
rect 539600 334698 539652 334704
rect 538220 330608 538272 330614
rect 538220 330550 538272 330556
rect 537576 273216 537628 273222
rect 537576 273158 537628 273164
rect 537484 259412 537536 259418
rect 537484 259354 537536 259360
rect 537024 239148 537076 239154
rect 537024 239090 537076 239096
rect 538232 16574 538260 330550
rect 538310 256592 538366 256601
rect 538310 256527 538366 256536
rect 538324 239902 538352 256527
rect 538402 254960 538458 254969
rect 538402 254895 538458 254904
rect 538312 239896 538364 239902
rect 538312 239838 538364 239844
rect 538416 237697 538444 254895
rect 538494 253600 538550 253609
rect 538494 253535 538550 253544
rect 538508 239970 538536 253535
rect 538496 239964 538548 239970
rect 538496 239906 538548 239912
rect 538402 237688 538458 237697
rect 538402 237623 538458 237632
rect 539612 16574 539640 334698
rect 540980 177404 541032 177410
rect 540980 177346 541032 177352
rect 540992 16574 541020 177346
rect 543752 16574 543780 335271
rect 547878 335200 547934 335209
rect 547878 335135 547934 335144
rect 536852 16546 537248 16574
rect 538232 16546 538444 16574
rect 539612 16546 540376 16574
rect 540992 16546 542032 16574
rect 543752 16546 544424 16574
rect 532514 7848 532570 7857
rect 532514 7783 532570 7792
rect 532528 480 532556 7783
rect 536102 7712 536158 7721
rect 536102 7647 536158 7656
rect 534908 4956 534960 4962
rect 534908 4898 534960 4904
rect 533712 3868 533764 3874
rect 533712 3810 533764 3816
rect 533724 480 533752 3810
rect 534920 480 534948 4898
rect 536116 480 536144 7647
rect 537220 480 537248 16546
rect 538416 480 538444 16546
rect 539598 7576 539654 7585
rect 539598 7511 539654 7520
rect 539612 480 539640 7511
rect 540348 490 540376 16546
rect 540624 598 540836 626
rect 540624 490 540652 598
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540348 462 540652 490
rect 540808 480 540836 598
rect 542004 480 542032 16546
rect 543188 9376 543240 9382
rect 543188 9318 543240 9324
rect 543200 480 543228 9318
rect 544396 480 544424 16546
rect 546684 9308 546736 9314
rect 546684 9250 546736 9256
rect 545488 4888 545540 4894
rect 545488 4830 545540 4836
rect 545500 480 545528 4830
rect 546696 480 546724 9250
rect 547892 480 547920 335135
rect 557538 335064 557594 335073
rect 557538 334999 557594 335008
rect 550640 334688 550692 334694
rect 550640 334630 550692 334636
rect 549260 177336 549312 177342
rect 549260 177278 549312 177284
rect 549272 16574 549300 177278
rect 550652 16574 550680 334630
rect 554780 334620 554832 334626
rect 554780 334562 554832 334568
rect 552018 332072 552074 332081
rect 552018 332007 552074 332016
rect 552032 16574 552060 332007
rect 554792 16574 554820 334562
rect 557552 16574 557580 334999
rect 561678 334928 561734 334937
rect 561678 334863 561734 334872
rect 561692 16574 561720 334863
rect 564438 334792 564494 334801
rect 564438 334727 564494 334736
rect 564452 16574 564480 334727
rect 567198 331936 567254 331945
rect 567198 331871 567254 331880
rect 567212 16574 567240 331871
rect 568592 16574 568620 336874
rect 569960 336864 570012 336870
rect 569960 336806 570012 336812
rect 569972 16574 570000 336806
rect 572720 336796 572772 336802
rect 572720 336738 572772 336744
rect 571338 331800 571394 331809
rect 571338 331735 571394 331744
rect 571352 16574 571380 331735
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 554792 16546 555004 16574
rect 557552 16546 558592 16574
rect 561692 16546 562088 16574
rect 564452 16546 565216 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 571352 16546 571564 16574
rect 549074 5264 549130 5273
rect 549074 5199 549130 5208
rect 549088 480 549116 5199
rect 550284 480 550312 16546
rect 551020 490 551048 16546
rect 551296 598 551508 626
rect 551296 490 551324 598
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 462 551324 490
rect 551480 480 551508 598
rect 552676 480 552704 16546
rect 553768 9240 553820 9246
rect 553768 9182 553820 9188
rect 553780 480 553808 9182
rect 554976 480 555004 16546
rect 557356 9172 557408 9178
rect 557356 9114 557408 9120
rect 556160 4820 556212 4826
rect 556160 4762 556212 4768
rect 556172 480 556200 4762
rect 557368 480 557396 9114
rect 558564 480 558592 16546
rect 560852 9104 560904 9110
rect 560852 9046 560904 9052
rect 559746 5128 559802 5137
rect 559746 5063 559802 5072
rect 559760 480 559788 5063
rect 560864 480 560892 9046
rect 562060 480 562088 16546
rect 564440 9036 564492 9042
rect 564440 8978 564492 8984
rect 563242 4992 563298 5001
rect 563242 4927 563298 4936
rect 563256 480 563284 4927
rect 564452 480 564480 8978
rect 565188 490 565216 16546
rect 566830 4856 566886 4865
rect 566830 4791 566886 4800
rect 565464 598 565676 626
rect 565464 490 565492 598
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565188 462 565492 490
rect 565648 480 565676 598
rect 566844 480 566872 4791
rect 567580 490 567608 16546
rect 567856 598 568068 626
rect 567856 490 567884 598
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 462 567884 490
rect 568040 480 568068 598
rect 568684 490 568712 16546
rect 568960 598 569172 626
rect 568960 490 568988 598
rect 567998 -960 568110 480
rect 568684 462 568988 490
rect 569144 480 569172 598
rect 570340 480 570368 16546
rect 571536 480 571564 16546
rect 572732 480 572760 336738
rect 575478 334656 575534 334665
rect 575478 334591 575534 334600
rect 574100 330540 574152 330546
rect 574100 330482 574152 330488
rect 574112 16574 574140 330482
rect 575492 16574 575520 334591
rect 576858 333296 576914 333305
rect 576858 333231 576914 333240
rect 576872 16574 576900 333231
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 579988 219428 580040 219434
rect 579988 219370 580040 219376
rect 580000 219065 580028 219370
rect 579986 219056 580042 219065
rect 579986 218991 580042 219000
rect 579620 193180 579672 193186
rect 579620 193122 579672 193128
rect 579632 192545 579660 193122
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 579620 179376 579672 179382
rect 579620 179318 579672 179324
rect 579632 179217 579660 179318
rect 579618 179208 579674 179217
rect 579618 179143 579674 179152
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 579620 126948 579672 126954
rect 579620 126890 579672 126896
rect 579632 126041 579660 126890
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 579620 86964 579672 86970
rect 579620 86906 579672 86912
rect 579632 86193 579660 86906
rect 579618 86184 579674 86193
rect 579618 86119 579674 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580276 46345 580304 386378
rect 580368 59673 580396 389127
rect 580908 388204 580960 388210
rect 580908 388146 580960 388152
rect 580816 388136 580868 388142
rect 580816 388078 580868 388084
rect 580724 388068 580776 388074
rect 580724 388010 580776 388016
rect 580632 388000 580684 388006
rect 580632 387942 580684 387948
rect 580540 387932 580592 387938
rect 580540 387874 580592 387880
rect 580448 387864 580500 387870
rect 580448 387806 580500 387812
rect 580460 112849 580488 387806
rect 580552 165889 580580 387874
rect 580644 205737 580672 387942
rect 580736 245585 580764 388010
rect 580828 298761 580856 388078
rect 580920 325281 580948 388146
rect 581000 331900 581052 331906
rect 581000 331842 581052 331848
rect 580906 325272 580962 325281
rect 580906 325207 580962 325216
rect 580908 320884 580960 320890
rect 580908 320826 580960 320832
rect 580920 312089 580948 320826
rect 580906 312080 580962 312089
rect 580906 312015 580962 312024
rect 580814 298752 580870 298761
rect 580814 298687 580870 298696
rect 580722 245576 580778 245585
rect 580722 245511 580778 245520
rect 580630 205728 580686 205737
rect 580630 205663 580686 205672
rect 580538 165880 580594 165889
rect 580538 165815 580594 165824
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580354 59664 580410 59673
rect 580354 59599 580410 59608
rect 580262 46336 580318 46345
rect 580262 46271 580318 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 576872 16546 576992 16574
rect 573916 8968 573968 8974
rect 573916 8910 573968 8916
rect 573928 480 573956 8910
rect 575124 480 575152 16546
rect 575860 490 575888 16546
rect 576136 598 576348 626
rect 576136 490 576164 598
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 462 576164 490
rect 576320 480 576348 598
rect 576964 490 576992 16546
rect 578606 8936 578662 8945
rect 578606 8871 578662 8880
rect 577240 598 577452 626
rect 577240 490 577268 598
rect 576278 -960 576390 480
rect 576964 462 577268 490
rect 577424 480 577452 598
rect 578620 480 578648 8871
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581012 480 581040 331842
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 582194 3360 582250 3369
rect 582194 3295 582250 3304
rect 582208 480 582236 3295
rect 583404 480 583432 3402
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 3146 410488 3202 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3422 387912 3478 387968
rect 3330 371320 3386 371376
rect 2778 358436 2780 358456
rect 2780 358436 2832 358456
rect 2832 358436 2834 358456
rect 2778 358400 2834 358436
rect 2778 345344 2834 345400
rect 2686 333376 2742 333432
rect 18 333240 74 333296
rect 3330 306212 3332 306232
rect 3332 306212 3384 306232
rect 3384 306212 3386 306232
rect 3330 306176 3386 306212
rect 2778 254088 2834 254144
rect 2778 241032 2834 241088
rect 2962 201864 3018 201920
rect 2778 188808 2834 188864
rect 3146 149776 3202 149832
rect 2778 136720 2834 136776
rect 3238 97552 3294 97608
rect 2778 84632 2834 84688
rect 2962 58520 3018 58576
rect 2778 45500 2780 45520
rect 2780 45500 2832 45520
rect 2832 45500 2834 45520
rect 2778 45464 2834 45500
rect 4802 389272 4858 389328
rect 4066 319232 4122 319288
rect 3974 293120 4030 293176
rect 3882 267144 3938 267200
rect 3790 214920 3846 214976
rect 3698 162832 3754 162888
rect 3606 110608 3662 110664
rect 3514 71576 3570 71632
rect 3422 32408 3478 32464
rect 2962 19352 3018 19408
rect 2778 6468 2780 6488
rect 2780 6468 2832 6488
rect 2832 6468 2834 6488
rect 2778 6432 2834 6468
rect 2870 4800 2926 4856
rect 6182 389408 6238 389464
rect 236274 389544 236330 389600
rect 235584 388048 235640 388104
rect 237194 389136 237250 389192
rect 236872 388184 236928 388240
rect 237930 388320 237986 388376
rect 270222 389836 270278 389872
rect 270222 389816 270224 389836
rect 270224 389816 270276 389836
rect 270276 389816 270278 389836
rect 271602 389816 271658 389872
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 281906 389408 281962 389464
rect 281538 389272 281594 389328
rect 281078 387912 281134 387968
rect 285126 388320 285182 388376
rect 233054 385192 233110 385248
rect 232962 379616 233018 379672
rect 232870 374040 232926 374096
rect 232778 368464 232834 368520
rect 232686 357312 232742 357368
rect 232594 346160 232650 346216
rect 232502 340720 232558 340776
rect 68926 336640 68982 336696
rect 62026 336504 62082 336560
rect 19338 335552 19394 335608
rect 11058 335416 11114 335472
rect 16578 334600 16634 334656
rect 15934 3304 15990 3360
rect 28814 335960 28870 336016
rect 26238 334736 26294 334792
rect 25318 3440 25374 3496
rect 37186 336232 37242 336288
rect 35806 336096 35862 336152
rect 53746 336368 53802 336424
rect 52366 333648 52422 333704
rect 48226 333512 48282 333568
rect 55126 333784 55182 333840
rect 56046 6160 56102 6216
rect 92386 334872 92442 334928
rect 86866 6296 86922 6352
rect 90362 6432 90418 6488
rect 93950 6568 94006 6624
rect 136546 335280 136602 335336
rect 133786 335144 133842 335200
rect 129646 335008 129702 335064
rect 128174 4936 128230 4992
rect 131762 5072 131818 5128
rect 144826 334464 144882 334520
rect 137650 5208 137706 5264
rect 226246 4156 226248 4176
rect 226248 4156 226300 4176
rect 226300 4156 226302 4176
rect 226246 4120 226302 4156
rect 234526 362888 234582 362944
rect 234434 351736 234490 351792
rect 233054 238584 233110 238640
rect 232962 238448 233018 238504
rect 232870 237904 232926 237960
rect 227718 4156 227720 4176
rect 227720 4156 227772 4176
rect 227772 4156 227774 4176
rect 227718 4120 227774 4156
rect 232042 3984 232098 4040
rect 234434 237088 234490 237144
rect 234710 333240 234766 333296
rect 234526 236272 234582 236328
rect 234434 4664 234490 4720
rect 234066 3984 234122 4040
rect 235078 333376 235134 333432
rect 235584 337864 235640 337920
rect 235630 337728 235686 337784
rect 235538 335416 235594 335472
rect 236274 335688 236330 335744
rect 235906 335416 235962 335472
rect 235906 334600 235962 334656
rect 235446 238856 235502 238912
rect 234802 4800 234858 4856
rect 236734 335552 236790 335608
rect 236642 334736 236698 334792
rect 236090 240080 236146 240136
rect 235722 4664 235778 4720
rect 237010 337592 237066 337648
rect 237010 336640 237066 336696
rect 236826 240080 236882 240136
rect 237010 238992 237066 239048
rect 236826 238720 236882 238776
rect 236826 3440 236882 3496
rect 237470 337728 237526 337784
rect 237378 335960 237434 336016
rect 237286 335824 237342 335880
rect 238252 337864 238308 337920
rect 237654 335824 237710 335880
rect 237930 336232 237986 336288
rect 237838 336096 237894 336152
rect 238022 335552 238078 335608
rect 237930 334056 237986 334112
rect 238574 334872 238630 334928
rect 239034 335552 239090 335608
rect 238942 333512 238998 333568
rect 239218 333648 239274 333704
rect 239494 336368 239550 336424
rect 239586 333784 239642 333840
rect 240368 337864 240424 337920
rect 240046 336504 240102 336560
rect 238942 6160 238998 6216
rect 240414 337728 240470 337784
rect 240690 337592 240746 337648
rect 236642 3304 236698 3360
rect 241978 337592 242034 337648
rect 241702 6568 241758 6624
rect 241794 6432 241850 6488
rect 242760 337762 242816 337818
rect 241886 6296 241942 6352
rect 243358 335824 243414 335880
rect 244968 337898 245024 337954
rect 243726 337592 243782 337648
rect 244968 337728 245024 337784
rect 245704 337898 245760 337954
rect 245888 337898 245944 337954
rect 245842 337592 245898 337648
rect 246210 335144 246266 335200
rect 245842 5072 245898 5128
rect 246578 335280 246634 335336
rect 246486 5208 246542 5264
rect 247038 334464 247094 334520
rect 247406 337728 247462 337784
rect 247774 337728 247830 337784
rect 248280 337898 248336 337954
rect 248004 337728 248060 337784
rect 249154 334056 249210 334112
rect 250488 337898 250544 337954
rect 250672 337898 250728 337954
rect 246578 4936 246634 4992
rect 250442 337728 250498 337784
rect 251592 337898 251648 337954
rect 251270 337592 251326 337648
rect 251546 337728 251602 337784
rect 251960 337898 252016 337954
rect 253478 337456 253534 337512
rect 254168 337898 254224 337954
rect 254214 337592 254270 337648
rect 254398 326440 254454 326496
rect 254214 326168 254270 326224
rect 255640 337830 255696 337886
rect 256146 337728 256202 337784
rect 255318 335416 255374 335472
rect 256376 337728 256432 337784
rect 257296 337864 257352 337920
rect 257664 337898 257720 337954
rect 257342 337728 257398 337784
rect 256238 239128 256294 239184
rect 257434 337592 257490 337648
rect 261896 337898 261952 337954
rect 261942 337728 261998 337784
rect 263368 337864 263424 337920
rect 263414 337728 263470 337784
rect 263736 337898 263792 337954
rect 264472 337864 264528 337920
rect 264334 337592 264390 337648
rect 268336 337830 268392 337886
rect 268474 337592 268530 337648
rect 268382 333240 268438 333296
rect 269118 335724 269120 335744
rect 269120 335724 269172 335744
rect 269172 335724 269174 335744
rect 269118 335688 269174 335724
rect 269118 333512 269174 333568
rect 269394 6432 269450 6488
rect 270820 337898 270876 337954
rect 270222 6296 270278 6352
rect 270958 6160 271014 6216
rect 272752 337864 272808 337920
rect 271786 335960 271842 336016
rect 272246 335552 272302 335608
rect 272430 335824 272486 335880
rect 272890 333376 272946 333432
rect 273442 333784 273498 333840
rect 273350 333648 273406 333704
rect 273718 335416 273774 335472
rect 273994 335416 274050 335472
rect 274270 335144 274326 335200
rect 274454 336504 274510 336560
rect 274638 333512 274694 333568
rect 275282 337592 275338 337648
rect 275466 336368 275522 336424
rect 275558 335688 275614 335744
rect 275466 239264 275522 239320
rect 276432 337898 276488 337954
rect 276202 336096 276258 336152
rect 276202 335824 276258 335880
rect 276478 337728 276534 337784
rect 276938 336096 276994 336152
rect 276938 335824 276994 335880
rect 277628 337864 277684 337920
rect 277306 332152 277362 332208
rect 277950 337728 278006 337784
rect 277950 335416 278006 335472
rect 277950 239808 278006 239864
rect 278502 336232 278558 336288
rect 278686 336096 278742 336152
rect 279560 337898 279616 337954
rect 279146 336096 279202 336152
rect 279146 335588 279148 335608
rect 279148 335588 279200 335608
rect 279200 335588 279202 335608
rect 279146 335552 279202 335588
rect 279238 334464 279294 334520
rect 279514 337728 279570 337784
rect 279422 334600 279478 334656
rect 279422 239536 279478 239592
rect 279606 337628 279608 337648
rect 279608 337628 279660 337648
rect 279660 337628 279662 337648
rect 279606 337592 279662 337628
rect 279882 335552 279938 335608
rect 279514 239400 279570 239456
rect 279882 239672 279938 239728
rect 280480 337864 280536 337920
rect 280756 337898 280812 337954
rect 280710 337728 280766 337784
rect 280066 334756 280122 334792
rect 280066 334736 280068 334756
rect 280068 334736 280120 334756
rect 280120 334736 280122 334756
rect 280434 335416 280490 335472
rect 279974 7792 280030 7848
rect 280894 335280 280950 335336
rect 280434 5208 280490 5264
rect 281446 335144 281502 335200
rect 281630 335008 281686 335064
rect 281538 332016 281594 332072
rect 281262 7656 281318 7712
rect 281170 7520 281226 7576
rect 281722 5072 281778 5128
rect 282182 334736 282238 334792
rect 282642 335588 282644 335608
rect 282644 335588 282696 335608
rect 282696 335588 282698 335608
rect 282642 335552 282698 335588
rect 282642 334600 282698 334656
rect 283010 335588 283012 335608
rect 283012 335588 283064 335608
rect 283064 335588 283066 335608
rect 283010 335552 283066 335588
rect 282918 334872 282974 334928
rect 282826 334736 282882 334792
rect 283102 331880 283158 331936
rect 283378 336096 283434 336152
rect 283286 335688 283342 335744
rect 283194 331744 283250 331800
rect 283378 335552 283434 335608
rect 283976 337864 284032 337920
rect 283884 337728 283940 337784
rect 284114 337728 284170 337784
rect 283746 336096 283802 336152
rect 283746 335824 283802 335880
rect 283654 334600 283710 334656
rect 283838 333240 283894 333296
rect 282550 4936 282606 4992
rect 284666 335688 284722 335744
rect 284574 335416 284630 335472
rect 284574 331336 284630 331392
rect 284666 331200 284722 331256
rect 284114 8880 284170 8936
rect 282642 4800 282698 4856
rect 282274 3440 282330 3496
rect 285034 331336 285090 331392
rect 286322 388048 286378 388104
rect 285770 337864 285826 337920
rect 285586 337592 285642 337648
rect 285218 331200 285274 331256
rect 286506 388184 286562 388240
rect 286414 336232 286470 336288
rect 287610 387640 287666 387696
rect 287610 386960 287666 387016
rect 287518 386280 287574 386336
rect 287610 385600 287666 385656
rect 288346 385076 288402 385112
rect 288346 385056 288348 385076
rect 288348 385056 288400 385076
rect 288400 385056 288402 385076
rect 287794 384376 287850 384432
rect 287610 383016 287666 383072
rect 287702 371320 287758 371376
rect 287610 370096 287666 370152
rect 287610 368736 287666 368792
rect 287518 366832 287574 366888
rect 287426 366152 287482 366208
rect 287334 365472 287390 365528
rect 287150 364248 287206 364304
rect 287610 357040 287666 357096
rect 287426 356360 287482 356416
rect 287702 354456 287758 354512
rect 287610 353796 287666 353832
rect 287610 353776 287612 353796
rect 287612 353776 287664 353796
rect 287664 353776 287666 353796
rect 287610 347248 287666 347304
rect 287334 346024 287390 346080
rect 287518 344120 287574 344176
rect 287610 342760 287666 342816
rect 287702 341400 287758 341456
rect 288346 383716 288402 383752
rect 288346 383696 288348 383716
rect 288348 383696 288400 383716
rect 288400 383696 288402 383716
rect 288346 382356 288402 382392
rect 288346 382336 288348 382356
rect 288348 382336 288400 382356
rect 288400 382336 288402 382356
rect 288162 381792 288218 381848
rect 288346 381112 288402 381168
rect 288254 380432 288310 380488
rect 288346 379772 288402 379808
rect 288346 379752 288348 379772
rect 288348 379752 288400 379772
rect 288400 379752 288402 379772
rect 288254 379208 288310 379264
rect 288346 378528 288402 378584
rect 288254 377848 288310 377904
rect 288346 377168 288402 377224
rect 288346 376488 288402 376544
rect 288162 375944 288218 376000
rect 288346 375264 288402 375320
rect 288162 374584 288218 374640
rect 288254 373904 288310 373960
rect 288162 373360 288218 373416
rect 288346 372716 288348 372736
rect 288348 372716 288400 372736
rect 288400 372716 288402 372736
rect 288346 372680 288402 372716
rect 288254 372000 288310 372056
rect 288346 370640 288402 370696
rect 288254 369416 288310 369472
rect 288346 368056 288402 368112
rect 287978 367512 288034 367568
rect 288346 364792 288402 364848
rect 288162 363568 288218 363624
rect 288162 362888 288218 362944
rect 288254 362208 288310 362264
rect 288346 361684 288402 361720
rect 288346 361664 288348 361684
rect 288348 361664 288400 361684
rect 288400 361664 288402 361684
rect 288162 360984 288218 361040
rect 288346 360304 288402 360360
rect 288346 359624 288402 359680
rect 288162 358944 288218 359000
rect 288254 358400 288310 358456
rect 288346 357720 288402 357776
rect 288346 355816 288402 355872
rect 287978 355136 288034 355192
rect 287978 353096 288034 353152
rect 287886 352552 287942 352608
rect 288346 351908 288348 351928
rect 288348 351908 288400 351928
rect 288400 351908 288402 351928
rect 288346 351872 288402 351908
rect 288070 351192 288126 351248
rect 288346 350512 288402 350568
rect 288346 349968 288402 350024
rect 288254 349308 288310 349344
rect 288254 349288 288256 349308
rect 288256 349288 288308 349308
rect 288308 349288 288310 349308
rect 288346 348608 288402 348664
rect 288254 347948 288310 347984
rect 288254 347928 288256 347948
rect 288256 347928 288308 347948
rect 288308 347928 288310 347948
rect 288346 346724 288402 346760
rect 288346 346704 288348 346724
rect 288348 346704 288400 346724
rect 288400 346704 288402 346724
rect 288346 345344 288402 345400
rect 288162 344664 288218 344720
rect 288346 343440 288402 343496
rect 288162 342080 288218 342136
rect 288346 340856 288402 340912
rect 288254 340176 288310 340232
rect 288346 339532 288348 339552
rect 288348 339532 288400 339552
rect 288400 339532 288402 339552
rect 288346 339496 288402 339532
rect 288254 338816 288310 338872
rect 288346 338272 288402 338328
rect 290554 336504 290610 336560
rect 290738 3712 290794 3768
rect 290922 3576 290978 3632
rect 292026 238040 292082 238096
rect 311162 389544 311218 389600
rect 293222 336368 293278 336424
rect 292210 237768 292266 237824
rect 293406 238312 293462 238368
rect 294694 238176 294750 238232
rect 297454 236952 297510 237008
rect 298834 236680 298890 236736
rect 299018 236816 299074 236872
rect 309782 336232 309838 336288
rect 308402 335960 308458 336016
rect 319442 336096 319498 336152
rect 309874 3304 309930 3360
rect 400862 332152 400918 332208
rect 407762 334464 407818 334520
rect 409142 333784 409198 333840
rect 414662 333648 414718 333704
rect 410798 6432 410854 6488
rect 414294 6296 414350 6352
rect 417422 333512 417478 333568
rect 428462 6160 428518 6216
rect 436926 271224 436982 271280
rect 437386 274080 437442 274136
rect 437110 272992 437166 273048
rect 437018 270000 437074 270056
rect 436926 268368 436982 268424
rect 436834 267416 436890 267472
rect 436742 265648 436798 265704
rect 436098 247288 436154 247344
rect 436098 245556 436100 245576
rect 436100 245556 436152 245576
rect 436152 245556 436154 245576
rect 436098 245520 436154 245556
rect 437202 237632 437258 237688
rect 438766 272992 438822 273048
rect 438674 271224 438730 271280
rect 439410 236544 439466 236600
rect 439594 333376 439650 333432
rect 467838 322496 467894 322552
rect 470598 322768 470654 322824
rect 470506 322632 470562 322688
rect 469402 321544 469458 321600
rect 472070 322496 472126 322552
rect 474738 322496 474794 322552
rect 478878 322496 478934 322552
rect 480258 322496 480314 322552
rect 481638 322496 481694 322552
rect 483018 322496 483074 322552
rect 486330 322496 486386 322552
rect 488538 322496 488594 322552
rect 489918 322496 489974 322552
rect 491298 322496 491354 322552
rect 496818 322496 496874 322552
rect 471978 321544 472034 321600
rect 474554 321544 474610 321600
rect 476762 321544 476818 321600
rect 478234 321544 478290 321600
rect 484398 321544 484454 321600
rect 485410 321544 485466 321600
rect 519542 322360 519598 322416
rect 488170 321580 488172 321600
rect 488172 321580 488224 321600
rect 488224 321580 488226 321600
rect 488170 321544 488226 321580
rect 492770 321544 492826 321600
rect 494242 321544 494298 321600
rect 495530 321544 495586 321600
rect 498198 321544 498254 321600
rect 499210 321544 499266 321600
rect 500682 321544 500738 321600
rect 501234 321544 501290 321600
rect 503258 321544 503314 321600
rect 503810 321544 503866 321600
rect 505466 321544 505522 321600
rect 506938 321544 506994 321600
rect 530030 321580 530032 321600
rect 530032 321580 530084 321600
rect 530084 321580 530086 321600
rect 530030 321544 530086 321580
rect 470506 319912 470562 319968
rect 502338 239808 502394 239864
rect 523130 239808 523186 239864
rect 452106 239128 452162 239184
rect 451646 238856 451702 238912
rect 456798 238992 456854 239048
rect 457074 238856 457130 238912
rect 452106 238720 452162 238776
rect 452290 238720 452346 238776
rect 461582 237904 461638 237960
rect 463698 237904 463754 237960
rect 465078 237904 465134 237960
rect 459558 237496 459614 237552
rect 447046 237224 447102 237280
rect 460938 237224 460994 237280
rect 446402 236408 446458 236464
rect 462410 236020 462466 236056
rect 462410 236000 462412 236020
rect 462412 236000 462464 236020
rect 462464 236000 462466 236020
rect 467838 239128 467894 239184
rect 469218 239128 469274 239184
rect 470690 238040 470746 238096
rect 471794 238040 471850 238096
rect 467194 237904 467250 237960
rect 468298 237904 468354 237960
rect 469218 237224 469274 237280
rect 471978 237224 472034 237280
rect 472070 236544 472126 236600
rect 471978 236292 472034 236328
rect 471978 236272 471980 236292
rect 471980 236272 472032 236292
rect 472032 236272 472034 236292
rect 475658 238040 475714 238096
rect 473450 236544 473506 236600
rect 480442 238992 480498 239048
rect 479154 238876 479210 238912
rect 479154 238856 479156 238876
rect 479156 238856 479208 238876
rect 479208 238856 479210 238876
rect 476762 238740 476818 238776
rect 476762 238720 476764 238740
rect 476764 238720 476816 238740
rect 476816 238720 476818 238740
rect 477590 238720 477646 238776
rect 477498 236544 477554 236600
rect 481638 237224 481694 237280
rect 480258 236680 480314 236736
rect 480534 236564 480590 236600
rect 480534 236544 480536 236564
rect 480536 236544 480588 236564
rect 480588 236544 480590 236564
rect 484582 239264 484638 239320
rect 483018 239012 483074 239048
rect 483018 238992 483020 239012
rect 483020 238992 483072 239012
rect 483072 238992 483074 239012
rect 483662 238448 483718 238504
rect 483662 238040 483718 238096
rect 481914 237224 481970 237280
rect 483018 237088 483074 237144
rect 484398 236816 484454 236872
rect 494242 238856 494298 238912
rect 484858 238468 484914 238504
rect 484858 238448 484860 238468
rect 484860 238448 484912 238468
rect 484912 238448 484914 238468
rect 490562 238604 490618 238640
rect 490562 238584 490564 238604
rect 490564 238584 490616 238604
rect 490616 238584 490618 238604
rect 485410 238484 485412 238504
rect 485412 238484 485464 238504
rect 485464 238484 485466 238504
rect 485410 238448 485466 238484
rect 487802 238448 487858 238504
rect 491666 238448 491722 238504
rect 492770 238332 492826 238368
rect 492770 238312 492772 238332
rect 492772 238312 492824 238332
rect 492824 238312 492826 238332
rect 496818 238312 496874 238368
rect 499210 238196 499266 238232
rect 499210 238176 499212 238196
rect 499212 238176 499264 238196
rect 499264 238176 499266 238196
rect 487158 237224 487214 237280
rect 492678 237224 492734 237280
rect 493322 237244 493378 237280
rect 493322 237224 493324 237244
rect 493324 237224 493376 237244
rect 493376 237224 493378 237244
rect 495438 237260 495440 237280
rect 495440 237260 495492 237280
rect 495492 237260 495494 237280
rect 495438 237224 495494 237260
rect 500958 237224 501014 237280
rect 488538 237088 488594 237144
rect 496818 237108 496874 237144
rect 496818 237088 496820 237108
rect 496820 237088 496872 237108
rect 496872 237088 496874 237108
rect 499854 237088 499910 237144
rect 491298 236836 491354 236872
rect 491298 236816 491300 236836
rect 491300 236816 491352 236836
rect 491352 236816 491354 236836
rect 485778 236700 485834 236736
rect 485778 236680 485780 236700
rect 485780 236680 485832 236700
rect 485832 236680 485834 236700
rect 485778 236408 485834 236464
rect 520278 239672 520334 239728
rect 503718 236680 503774 236736
rect 502430 236000 502486 236056
rect 505098 236272 505154 236328
rect 472254 3712 472310 3768
rect 479338 3576 479394 3632
rect 484030 3440 484086 3496
rect 522670 239536 522726 239592
rect 522854 239536 522910 239592
rect 523222 239400 523278 239456
rect 523038 237224 523094 237280
rect 527178 239264 527234 239320
rect 537114 316512 537170 316568
rect 580354 389136 580410 389192
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 543738 335280 543794 335336
rect 538310 256536 538366 256592
rect 538402 254904 538458 254960
rect 538494 253544 538550 253600
rect 538402 237632 538458 237688
rect 547878 335144 547934 335200
rect 532514 7792 532570 7848
rect 536102 7656 536158 7712
rect 539598 7520 539654 7576
rect 557538 335008 557594 335064
rect 552018 332016 552074 332072
rect 561678 334872 561734 334928
rect 564438 334736 564494 334792
rect 567198 331880 567254 331936
rect 571338 331744 571394 331800
rect 549074 5208 549130 5264
rect 559746 5072 559802 5128
rect 563242 4936 563298 4992
rect 566830 4800 566886 4856
rect 575478 334600 575534 334656
rect 576858 333240 576914 333296
rect 580170 272176 580226 272232
rect 579802 258848 579858 258904
rect 579986 232328 580042 232384
rect 579986 219000 580042 219056
rect 579618 192480 579674 192536
rect 579618 179152 579674 179208
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 579618 125976 579674 126032
rect 580170 99456 580226 99512
rect 579618 86128 579674 86184
rect 580170 72936 580226 72992
rect 580906 325216 580962 325272
rect 580906 312024 580962 312080
rect 580814 298696 580870 298752
rect 580722 245520 580778 245576
rect 580630 205672 580686 205728
rect 580538 165824 580594 165880
rect 580446 112784 580502 112840
rect 580354 59608 580410 59664
rect 580262 46280 580318 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 578606 8880 578662 8936
rect 580170 6568 580226 6624
rect 582194 3304 582250 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 583520 391628 584960 391868
rect 270217 389874 270283 389877
rect 271597 389874 271663 389877
rect 270217 389872 271663 389874
rect 270217 389816 270222 389872
rect 270278 389816 271602 389872
rect 271658 389816 271663 389872
rect 270217 389814 271663 389816
rect 270217 389811 270283 389814
rect 271597 389811 271663 389814
rect 236269 389602 236335 389605
rect 311157 389602 311223 389605
rect 236269 389600 311223 389602
rect 236269 389544 236274 389600
rect 236330 389544 311162 389600
rect 311218 389544 311223 389600
rect 236269 389542 311223 389544
rect 236269 389539 236335 389542
rect 311157 389539 311223 389542
rect 6177 389466 6243 389469
rect 281901 389466 281967 389469
rect 6177 389464 281967 389466
rect 6177 389408 6182 389464
rect 6238 389408 281906 389464
rect 281962 389408 281967 389464
rect 6177 389406 281967 389408
rect 6177 389403 6243 389406
rect 281901 389403 281967 389406
rect 4797 389330 4863 389333
rect 281533 389330 281599 389333
rect 4797 389328 281599 389330
rect 4797 389272 4802 389328
rect 4858 389272 281538 389328
rect 281594 389272 281599 389328
rect 4797 389270 281599 389272
rect 4797 389267 4863 389270
rect 281533 389267 281599 389270
rect 237189 389194 237255 389197
rect 580349 389194 580415 389197
rect 237189 389192 580415 389194
rect 237189 389136 237194 389192
rect 237250 389136 580354 389192
rect 580410 389136 580415 389192
rect 237189 389134 580415 389136
rect 237189 389131 237255 389134
rect 580349 389131 580415 389134
rect 237925 388378 237991 388381
rect 285121 388378 285187 388381
rect 237925 388376 285187 388378
rect 237925 388320 237930 388376
rect 237986 388320 285126 388376
rect 285182 388320 285187 388376
rect 237925 388318 285187 388320
rect 237925 388315 237991 388318
rect 285121 388315 285187 388318
rect 236867 388242 236933 388245
rect 286501 388242 286567 388245
rect 236867 388240 286567 388242
rect 236867 388184 236872 388240
rect 236928 388184 286506 388240
rect 286562 388184 286567 388240
rect 236867 388182 286567 388184
rect 236867 388179 236933 388182
rect 286501 388179 286567 388182
rect 235579 388106 235645 388109
rect 286317 388106 286383 388109
rect 235579 388104 286383 388106
rect 235579 388048 235584 388104
rect 235640 388048 286322 388104
rect 286378 388048 286383 388104
rect 235579 388046 286383 388048
rect 235579 388043 235645 388046
rect 286317 388043 286383 388046
rect 3417 387970 3483 387973
rect 281073 387970 281139 387973
rect 3417 387968 281139 387970
rect 3417 387912 3422 387968
rect 3478 387912 281078 387968
rect 281134 387912 281139 387968
rect 3417 387910 281139 387912
rect 3417 387907 3483 387910
rect 281073 387907 281139 387910
rect 287605 387698 287671 387701
rect 284924 387696 287671 387698
rect 284924 387640 287610 387696
rect 287666 387640 287671 387696
rect 284924 387638 287671 387640
rect 287605 387635 287671 387638
rect 287605 387018 287671 387021
rect 284924 387016 287671 387018
rect 284924 386960 287610 387016
rect 287666 386960 287671 387016
rect 284924 386958 287671 386960
rect 287605 386955 287671 386958
rect 287513 386338 287579 386341
rect 284924 386336 287579 386338
rect 284924 386280 287518 386336
rect 287574 386280 287579 386336
rect 284924 386278 287579 386280
rect 287513 386275 287579 386278
rect 287605 385658 287671 385661
rect 284924 385656 287671 385658
rect 284924 385600 287610 385656
rect 287666 385600 287671 385656
rect 284924 385598 287671 385600
rect 287605 385595 287671 385598
rect 233049 385250 233115 385253
rect 233049 385248 235060 385250
rect 233049 385192 233054 385248
rect 233110 385192 235060 385248
rect 233049 385190 235060 385192
rect 233049 385187 233115 385190
rect 288341 385114 288407 385117
rect 284924 385112 288407 385114
rect 284924 385056 288346 385112
rect 288402 385056 288407 385112
rect 284924 385054 288407 385056
rect 288341 385051 288407 385054
rect -960 384284 480 384524
rect 287789 384434 287855 384437
rect 284924 384432 287855 384434
rect 284924 384376 287794 384432
rect 287850 384376 287855 384432
rect 284924 384374 287855 384376
rect 287789 384371 287855 384374
rect 288341 383754 288407 383757
rect 284924 383752 288407 383754
rect 284924 383696 288346 383752
rect 288402 383696 288407 383752
rect 284924 383694 288407 383696
rect 288341 383691 288407 383694
rect 287605 383074 287671 383077
rect 284924 383072 287671 383074
rect 284924 383016 287610 383072
rect 287666 383016 287671 383072
rect 284924 383014 287671 383016
rect 287605 383011 287671 383014
rect 288341 382394 288407 382397
rect 284924 382392 288407 382394
rect 284924 382336 288346 382392
rect 288402 382336 288407 382392
rect 284924 382334 288407 382336
rect 288341 382331 288407 382334
rect 288157 381850 288223 381853
rect 284924 381848 288223 381850
rect 284924 381792 288162 381848
rect 288218 381792 288223 381848
rect 284924 381790 288223 381792
rect 288157 381787 288223 381790
rect 288341 381170 288407 381173
rect 284924 381168 288407 381170
rect 284924 381112 288346 381168
rect 288402 381112 288407 381168
rect 284924 381110 288407 381112
rect 288341 381107 288407 381110
rect 288249 380490 288315 380493
rect 284924 380488 288315 380490
rect 284924 380432 288254 380488
rect 288310 380432 288315 380488
rect 284924 380430 288315 380432
rect 288249 380427 288315 380430
rect 288341 379810 288407 379813
rect 284924 379808 288407 379810
rect 284924 379752 288346 379808
rect 288402 379752 288407 379808
rect 284924 379750 288407 379752
rect 288341 379747 288407 379750
rect 232957 379674 233023 379677
rect 232957 379672 235060 379674
rect 232957 379616 232962 379672
rect 233018 379616 235060 379672
rect 232957 379614 235060 379616
rect 232957 379611 233023 379614
rect 288249 379266 288315 379269
rect 284924 379264 288315 379266
rect 284924 379208 288254 379264
rect 288310 379208 288315 379264
rect 284924 379206 288315 379208
rect 288249 379203 288315 379206
rect 288341 378586 288407 378589
rect 284924 378584 288407 378586
rect 284924 378528 288346 378584
rect 288402 378528 288407 378584
rect 284924 378526 288407 378528
rect 288341 378523 288407 378526
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 288249 377906 288315 377909
rect 284924 377904 288315 377906
rect 284924 377848 288254 377904
rect 288310 377848 288315 377904
rect 284924 377846 288315 377848
rect 288249 377843 288315 377846
rect 288341 377226 288407 377229
rect 284924 377224 288407 377226
rect 284924 377168 288346 377224
rect 288402 377168 288407 377224
rect 284924 377166 288407 377168
rect 288341 377163 288407 377166
rect 288341 376546 288407 376549
rect 284924 376544 288407 376546
rect 284924 376488 288346 376544
rect 288402 376488 288407 376544
rect 284924 376486 288407 376488
rect 288341 376483 288407 376486
rect 288157 376002 288223 376005
rect 284924 376000 288223 376002
rect 284924 375944 288162 376000
rect 288218 375944 288223 376000
rect 284924 375942 288223 375944
rect 288157 375939 288223 375942
rect 288341 375322 288407 375325
rect 284924 375320 288407 375322
rect 284924 375264 288346 375320
rect 288402 375264 288407 375320
rect 284924 375262 288407 375264
rect 288341 375259 288407 375262
rect 288157 374642 288223 374645
rect 284924 374640 288223 374642
rect 284924 374584 288162 374640
rect 288218 374584 288223 374640
rect 284924 374582 288223 374584
rect 288157 374579 288223 374582
rect 232865 374098 232931 374101
rect 232865 374096 235060 374098
rect 232865 374040 232870 374096
rect 232926 374040 235060 374096
rect 232865 374038 235060 374040
rect 232865 374035 232931 374038
rect 288249 373962 288315 373965
rect 284924 373960 288315 373962
rect 284924 373904 288254 373960
rect 288310 373904 288315 373960
rect 284924 373902 288315 373904
rect 288249 373899 288315 373902
rect 288157 373418 288223 373421
rect 284924 373416 288223 373418
rect 284924 373360 288162 373416
rect 288218 373360 288223 373416
rect 284924 373358 288223 373360
rect 288157 373355 288223 373358
rect 288341 372738 288407 372741
rect 284924 372736 288407 372738
rect 284924 372680 288346 372736
rect 288402 372680 288407 372736
rect 284924 372678 288407 372680
rect 288341 372675 288407 372678
rect 288249 372058 288315 372061
rect 284924 372056 288315 372058
rect 284924 372000 288254 372056
rect 288310 372000 288315 372056
rect 284924 371998 288315 372000
rect 288249 371995 288315 371998
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect 287697 371378 287763 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect 284924 371376 287763 371378
rect 284924 371320 287702 371376
rect 287758 371320 287763 371376
rect 284924 371318 287763 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 287697 371315 287763 371318
rect 288341 370698 288407 370701
rect 284924 370696 288407 370698
rect 284924 370640 288346 370696
rect 288402 370640 288407 370696
rect 284924 370638 288407 370640
rect 288341 370635 288407 370638
rect 287605 370154 287671 370157
rect 284924 370152 287671 370154
rect 284924 370096 287610 370152
rect 287666 370096 287671 370152
rect 284924 370094 287671 370096
rect 287605 370091 287671 370094
rect 288249 369474 288315 369477
rect 284924 369472 288315 369474
rect 284924 369416 288254 369472
rect 288310 369416 288315 369472
rect 284924 369414 288315 369416
rect 288249 369411 288315 369414
rect 287605 368794 287671 368797
rect 284924 368792 287671 368794
rect 284924 368736 287610 368792
rect 287666 368736 287671 368792
rect 284924 368734 287671 368736
rect 287605 368731 287671 368734
rect 232773 368522 232839 368525
rect 232773 368520 235060 368522
rect 232773 368464 232778 368520
rect 232834 368464 235060 368520
rect 232773 368462 235060 368464
rect 232773 368459 232839 368462
rect 288341 368114 288407 368117
rect 284924 368112 288407 368114
rect 284924 368056 288346 368112
rect 288402 368056 288407 368112
rect 284924 368054 288407 368056
rect 288341 368051 288407 368054
rect 287973 367570 288039 367573
rect 284924 367568 288039 367570
rect 284924 367512 287978 367568
rect 288034 367512 288039 367568
rect 284924 367510 288039 367512
rect 287973 367507 288039 367510
rect 287513 366890 287579 366893
rect 284924 366888 287579 366890
rect 284924 366832 287518 366888
rect 287574 366832 287579 366888
rect 284924 366830 287579 366832
rect 287513 366827 287579 366830
rect 287421 366210 287487 366213
rect 284924 366208 287487 366210
rect 284924 366152 287426 366208
rect 287482 366152 287487 366208
rect 284924 366150 287487 366152
rect 287421 366147 287487 366150
rect 287329 365530 287395 365533
rect 284924 365528 287395 365530
rect 284924 365472 287334 365528
rect 287390 365472 287395 365528
rect 284924 365470 287395 365472
rect 287329 365467 287395 365470
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 288341 364850 288407 364853
rect 284924 364848 288407 364850
rect 284924 364792 288346 364848
rect 288402 364792 288407 364848
rect 284924 364790 288407 364792
rect 288341 364787 288407 364790
rect 287145 364306 287211 364309
rect 284924 364304 287211 364306
rect 284924 364248 287150 364304
rect 287206 364248 287211 364304
rect 284924 364246 287211 364248
rect 287145 364243 287211 364246
rect 288157 363626 288223 363629
rect 284924 363624 288223 363626
rect 284924 363568 288162 363624
rect 288218 363568 288223 363624
rect 284924 363566 288223 363568
rect 288157 363563 288223 363566
rect 234521 362946 234587 362949
rect 288157 362946 288223 362949
rect 234521 362944 235060 362946
rect 234521 362888 234526 362944
rect 234582 362888 235060 362944
rect 234521 362886 235060 362888
rect 284924 362944 288223 362946
rect 284924 362888 288162 362944
rect 288218 362888 288223 362944
rect 284924 362886 288223 362888
rect 234521 362883 234587 362886
rect 288157 362883 288223 362886
rect 288249 362266 288315 362269
rect 284924 362264 288315 362266
rect 284924 362208 288254 362264
rect 288310 362208 288315 362264
rect 284924 362206 288315 362208
rect 288249 362203 288315 362206
rect 288341 361722 288407 361725
rect 284924 361720 288407 361722
rect 284924 361664 288346 361720
rect 288402 361664 288407 361720
rect 284924 361662 288407 361664
rect 288341 361659 288407 361662
rect 288157 361042 288223 361045
rect 284924 361040 288223 361042
rect 284924 360984 288162 361040
rect 288218 360984 288223 361040
rect 284924 360982 288223 360984
rect 288157 360979 288223 360982
rect 288341 360362 288407 360365
rect 284924 360360 288407 360362
rect 284924 360304 288346 360360
rect 288402 360304 288407 360360
rect 284924 360302 288407 360304
rect 288341 360299 288407 360302
rect 288341 359682 288407 359685
rect 284924 359680 288407 359682
rect 284924 359624 288346 359680
rect 288402 359624 288407 359680
rect 284924 359622 288407 359624
rect 288341 359619 288407 359622
rect 288157 359002 288223 359005
rect 284924 359000 288223 359002
rect 284924 358944 288162 359000
rect 288218 358944 288223 359000
rect 284924 358942 288223 358944
rect 288157 358939 288223 358942
rect -960 358458 480 358548
rect 2773 358458 2839 358461
rect 288249 358458 288315 358461
rect -960 358456 2839 358458
rect -960 358400 2778 358456
rect 2834 358400 2839 358456
rect -960 358398 2839 358400
rect 284924 358456 288315 358458
rect 284924 358400 288254 358456
rect 288310 358400 288315 358456
rect 284924 358398 288315 358400
rect -960 358308 480 358398
rect 2773 358395 2839 358398
rect 288249 358395 288315 358398
rect 288341 357778 288407 357781
rect 284924 357776 288407 357778
rect 284924 357720 288346 357776
rect 288402 357720 288407 357776
rect 284924 357718 288407 357720
rect 288341 357715 288407 357718
rect 232681 357370 232747 357373
rect 232681 357368 235060 357370
rect 232681 357312 232686 357368
rect 232742 357312 235060 357368
rect 232681 357310 235060 357312
rect 232681 357307 232747 357310
rect 287605 357098 287671 357101
rect 284924 357096 287671 357098
rect 284924 357040 287610 357096
rect 287666 357040 287671 357096
rect 284924 357038 287671 357040
rect 287605 357035 287671 357038
rect 287421 356418 287487 356421
rect 284924 356416 287487 356418
rect 284924 356360 287426 356416
rect 287482 356360 287487 356416
rect 284924 356358 287487 356360
rect 287421 356355 287487 356358
rect 288341 355874 288407 355877
rect 284924 355872 288407 355874
rect 284924 355816 288346 355872
rect 288402 355816 288407 355872
rect 284924 355814 288407 355816
rect 288341 355811 288407 355814
rect 287973 355194 288039 355197
rect 284924 355192 288039 355194
rect 284924 355136 287978 355192
rect 288034 355136 288039 355192
rect 284924 355134 288039 355136
rect 287973 355131 288039 355134
rect 287697 354514 287763 354517
rect 284924 354512 287763 354514
rect 284924 354456 287702 354512
rect 287758 354456 287763 354512
rect 284924 354454 287763 354456
rect 287697 354451 287763 354454
rect 287605 353834 287671 353837
rect 284924 353832 287671 353834
rect 284924 353776 287610 353832
rect 287666 353776 287671 353832
rect 284924 353774 287671 353776
rect 287605 353771 287671 353774
rect 287973 353154 288039 353157
rect 284924 353152 288039 353154
rect 284924 353096 287978 353152
rect 288034 353096 288039 353152
rect 284924 353094 288039 353096
rect 287973 353091 288039 353094
rect 287881 352610 287947 352613
rect 284924 352608 287947 352610
rect 284924 352552 287886 352608
rect 287942 352552 287947 352608
rect 284924 352550 287947 352552
rect 287881 352547 287947 352550
rect 288341 351930 288407 351933
rect 284924 351928 288407 351930
rect 284924 351872 288346 351928
rect 288402 351872 288407 351928
rect 284924 351870 288407 351872
rect 288341 351867 288407 351870
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 234429 351794 234495 351797
rect 234429 351792 235060 351794
rect 234429 351736 234434 351792
rect 234490 351736 235060 351792
rect 583520 351780 584960 351870
rect 234429 351734 235060 351736
rect 234429 351731 234495 351734
rect 288065 351250 288131 351253
rect 284924 351248 288131 351250
rect 284924 351192 288070 351248
rect 288126 351192 288131 351248
rect 284924 351190 288131 351192
rect 288065 351187 288131 351190
rect 288341 350570 288407 350573
rect 284924 350568 288407 350570
rect 284924 350512 288346 350568
rect 288402 350512 288407 350568
rect 284924 350510 288407 350512
rect 288341 350507 288407 350510
rect 288341 350026 288407 350029
rect 284924 350024 288407 350026
rect 284924 349968 288346 350024
rect 288402 349968 288407 350024
rect 284924 349966 288407 349968
rect 288341 349963 288407 349966
rect 288249 349346 288315 349349
rect 284924 349344 288315 349346
rect 284924 349288 288254 349344
rect 288310 349288 288315 349344
rect 284924 349286 288315 349288
rect 288249 349283 288315 349286
rect 288341 348666 288407 348669
rect 284924 348664 288407 348666
rect 284924 348608 288346 348664
rect 288402 348608 288407 348664
rect 284924 348606 288407 348608
rect 288341 348603 288407 348606
rect 288249 347986 288315 347989
rect 284924 347984 288315 347986
rect 284924 347928 288254 347984
rect 288310 347928 288315 347984
rect 284924 347926 288315 347928
rect 288249 347923 288315 347926
rect 287605 347306 287671 347309
rect 284924 347304 287671 347306
rect 284924 347248 287610 347304
rect 287666 347248 287671 347304
rect 284924 347246 287671 347248
rect 287605 347243 287671 347246
rect 288341 346762 288407 346765
rect 284924 346760 288407 346762
rect 284924 346704 288346 346760
rect 288402 346704 288407 346760
rect 284924 346702 288407 346704
rect 288341 346699 288407 346702
rect 232589 346218 232655 346221
rect 232589 346216 235060 346218
rect 232589 346160 232594 346216
rect 232650 346160 235060 346216
rect 232589 346158 235060 346160
rect 232589 346155 232655 346158
rect 287329 346082 287395 346085
rect 284924 346080 287395 346082
rect 284924 346024 287334 346080
rect 287390 346024 287395 346080
rect 284924 346022 287395 346024
rect 287329 346019 287395 346022
rect -960 345402 480 345492
rect 2773 345402 2839 345405
rect 288341 345402 288407 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect 284924 345400 288407 345402
rect 284924 345344 288346 345400
rect 288402 345344 288407 345400
rect 284924 345342 288407 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 288341 345339 288407 345342
rect 288157 344722 288223 344725
rect 284924 344720 288223 344722
rect 284924 344664 288162 344720
rect 288218 344664 288223 344720
rect 284924 344662 288223 344664
rect 288157 344659 288223 344662
rect 287513 344178 287579 344181
rect 284924 344176 287579 344178
rect 284924 344120 287518 344176
rect 287574 344120 287579 344176
rect 284924 344118 287579 344120
rect 287513 344115 287579 344118
rect 288341 343498 288407 343501
rect 284924 343496 288407 343498
rect 284924 343440 288346 343496
rect 288402 343440 288407 343496
rect 284924 343438 288407 343440
rect 288341 343435 288407 343438
rect 287605 342818 287671 342821
rect 284924 342816 287671 342818
rect 284924 342760 287610 342816
rect 287666 342760 287671 342816
rect 284924 342758 287671 342760
rect 287605 342755 287671 342758
rect 288157 342138 288223 342141
rect 284924 342136 288223 342138
rect 284924 342080 288162 342136
rect 288218 342080 288223 342136
rect 284924 342078 288223 342080
rect 288157 342075 288223 342078
rect 287697 341458 287763 341461
rect 284924 341456 287763 341458
rect 284924 341400 287702 341456
rect 287758 341400 287763 341456
rect 284924 341398 287763 341400
rect 287697 341395 287763 341398
rect 288341 340914 288407 340917
rect 284924 340912 288407 340914
rect 284924 340856 288346 340912
rect 288402 340856 288407 340912
rect 284924 340854 288407 340856
rect 288341 340851 288407 340854
rect 232497 340778 232563 340781
rect 232497 340776 235060 340778
rect 232497 340720 232502 340776
rect 232558 340720 235060 340776
rect 232497 340718 235060 340720
rect 232497 340715 232563 340718
rect 288249 340234 288315 340237
rect 284924 340232 288315 340234
rect 284924 340176 288254 340232
rect 288310 340176 288315 340232
rect 284924 340174 288315 340176
rect 288249 340171 288315 340174
rect 288341 339554 288407 339557
rect 284924 339552 288407 339554
rect 284924 339496 288346 339552
rect 288402 339496 288407 339552
rect 284924 339494 288407 339496
rect 288341 339491 288407 339494
rect 288249 338874 288315 338877
rect 284924 338872 288315 338874
rect 284924 338816 288254 338872
rect 288310 338816 288315 338872
rect 284924 338814 288315 338816
rect 288249 338811 288315 338814
rect 583520 338452 584960 338692
rect 288341 338330 288407 338333
rect 284924 338328 288407 338330
rect 284924 338272 288346 338328
rect 288402 338272 288407 338328
rect 284924 338270 288407 338272
rect 288341 338267 288407 338270
rect 244963 337954 245029 337959
rect 235579 337920 235645 337925
rect 238247 337922 238313 337925
rect 235579 337864 235584 337920
rect 235640 337864 235645 337920
rect 235579 337859 235645 337864
rect 237606 337920 238313 337922
rect 237606 337864 238252 337920
rect 238308 337864 238313 337920
rect 237606 337862 238313 337864
rect 235582 337789 235642 337859
rect 235582 337784 235691 337789
rect 235582 337728 235630 337784
rect 235686 337728 235691 337784
rect 235582 337726 235691 337728
rect 235625 337723 235691 337726
rect 237465 337786 237531 337789
rect 237606 337786 237666 337862
rect 238247 337859 238313 337862
rect 240363 337920 240429 337925
rect 240363 337864 240368 337920
rect 240424 337864 240429 337920
rect 244963 337898 244968 337954
rect 245024 337898 245029 337954
rect 244963 337893 245029 337898
rect 245699 337954 245765 337959
rect 245699 337898 245704 337954
rect 245760 337898 245765 337954
rect 245883 337956 245949 337959
rect 245883 337954 246006 337956
rect 245883 337924 245888 337954
rect 245944 337924 246006 337954
rect 245699 337893 245765 337898
rect 240363 337859 240429 337864
rect 237465 337784 237666 337786
rect 237465 337728 237470 337784
rect 237526 337728 237666 337784
rect 237465 337726 237666 337728
rect 240366 337789 240426 337859
rect 242755 337818 242821 337823
rect 240366 337784 240475 337789
rect 240366 337728 240414 337784
rect 240470 337728 240475 337784
rect 242755 337762 242760 337818
rect 242816 337762 242821 337818
rect 244966 337789 245026 337893
rect 242755 337757 242821 337762
rect 244963 337784 245029 337789
rect 240366 337726 240475 337728
rect 237465 337723 237531 337726
rect 240409 337723 240475 337726
rect 237005 337650 237071 337653
rect 240685 337650 240751 337653
rect 237005 337648 240751 337650
rect 237005 337592 237010 337648
rect 237066 337592 240690 337648
rect 240746 337592 240751 337648
rect 237005 337590 240751 337592
rect 237005 337587 237071 337590
rect 240685 337587 240751 337590
rect 241973 337650 242039 337653
rect 242758 337650 242818 337757
rect 244963 337728 244968 337784
rect 245024 337728 245029 337784
rect 244963 337723 245029 337728
rect 241973 337648 242818 337650
rect 241973 337592 241978 337648
rect 242034 337592 242818 337648
rect 241973 337590 242818 337592
rect 243721 337650 243787 337653
rect 245702 337650 245762 337893
rect 245878 337860 245884 337924
rect 245948 337896 246006 337924
rect 248275 337954 248341 337959
rect 248275 337922 248280 337954
rect 247542 337898 248280 337922
rect 248336 337898 248341 337954
rect 245948 337860 245954 337896
rect 247542 337893 248341 337898
rect 250483 337954 250549 337959
rect 250483 337898 250488 337954
rect 250544 337898 250549 337954
rect 250483 337893 250549 337898
rect 250667 337954 250733 337959
rect 250667 337898 250672 337954
rect 250728 337898 250733 337954
rect 250667 337893 250733 337898
rect 251587 337954 251653 337959
rect 251587 337898 251592 337954
rect 251648 337898 251653 337954
rect 251587 337893 251653 337898
rect 251955 337954 252021 337959
rect 251955 337898 251960 337954
rect 252016 337898 252021 337954
rect 251955 337893 252021 337898
rect 254163 337954 254229 337959
rect 254163 337898 254168 337954
rect 254224 337898 254229 337954
rect 257659 337954 257725 337959
rect 254163 337893 254229 337898
rect 257291 337920 257357 337925
rect 247542 337862 248338 337893
rect 247401 337786 247467 337789
rect 247542 337786 247602 337862
rect 250486 337789 250546 337893
rect 247401 337784 247602 337786
rect 247401 337728 247406 337784
rect 247462 337728 247602 337784
rect 247401 337726 247602 337728
rect 247769 337786 247835 337789
rect 247999 337786 248065 337789
rect 247769 337784 248065 337786
rect 247769 337728 247774 337784
rect 247830 337728 248004 337784
rect 248060 337728 248065 337784
rect 247769 337726 248065 337728
rect 247401 337723 247467 337726
rect 247769 337723 247835 337726
rect 247999 337723 248065 337726
rect 250437 337784 250546 337789
rect 250437 337728 250442 337784
rect 250498 337728 250546 337784
rect 250437 337726 250546 337728
rect 250437 337723 250503 337726
rect 243721 337648 245762 337650
rect 243721 337592 243726 337648
rect 243782 337592 245762 337648
rect 243721 337590 245762 337592
rect 245837 337650 245903 337653
rect 250670 337650 250730 337893
rect 251590 337789 251650 337893
rect 251541 337784 251650 337789
rect 251541 337728 251546 337784
rect 251602 337728 251650 337784
rect 251541 337726 251650 337728
rect 251541 337723 251607 337726
rect 245837 337648 250730 337650
rect 245837 337592 245842 337648
rect 245898 337592 250730 337648
rect 245837 337590 250730 337592
rect 251265 337650 251331 337653
rect 251958 337650 252018 337893
rect 251265 337648 252018 337650
rect 251265 337592 251270 337648
rect 251326 337592 252018 337648
rect 251265 337590 252018 337592
rect 254166 337653 254226 337893
rect 255635 337886 255701 337891
rect 255635 337830 255640 337886
rect 255696 337830 255701 337886
rect 257291 337864 257296 337920
rect 257352 337864 257357 337920
rect 257659 337898 257664 337954
rect 257720 337898 257725 337954
rect 257659 337893 257725 337898
rect 261891 337954 261957 337959
rect 261891 337898 261896 337954
rect 261952 337898 261957 337954
rect 263731 337956 263797 337959
rect 270815 337956 270881 337959
rect 263731 337954 263854 337956
rect 261891 337893 261957 337898
rect 263363 337920 263429 337925
rect 263731 337924 263736 337954
rect 263792 337924 263854 337954
rect 270815 337954 270924 337956
rect 257291 337859 257357 337864
rect 255635 337825 255701 337830
rect 254166 337648 254275 337653
rect 254166 337592 254214 337648
rect 254270 337592 254275 337648
rect 254166 337590 254275 337592
rect 241973 337587 242039 337590
rect 243721 337587 243787 337590
rect 245837 337587 245903 337590
rect 251265 337587 251331 337590
rect 254209 337587 254275 337590
rect 253473 337514 253539 337517
rect 255638 337514 255698 337825
rect 257294 337789 257354 337859
rect 256141 337786 256207 337789
rect 256371 337786 256437 337789
rect 256141 337784 256437 337786
rect 256141 337728 256146 337784
rect 256202 337728 256376 337784
rect 256432 337728 256437 337784
rect 256141 337726 256437 337728
rect 257294 337784 257403 337789
rect 257294 337728 257342 337784
rect 257398 337728 257403 337784
rect 257294 337726 257403 337728
rect 256141 337723 256207 337726
rect 256371 337723 256437 337726
rect 257337 337723 257403 337726
rect 257429 337650 257495 337653
rect 257662 337650 257722 337893
rect 261894 337789 261954 337893
rect 263363 337864 263368 337920
rect 263424 337864 263429 337920
rect 263363 337859 263429 337864
rect 263726 337860 263732 337924
rect 263796 337896 263854 337924
rect 264467 337920 264533 337925
rect 263796 337860 263802 337896
rect 264467 337864 264472 337920
rect 264528 337864 264533 337920
rect 270815 337898 270820 337954
rect 270876 337898 270924 337954
rect 276427 337954 276493 337959
rect 270815 337893 270924 337898
rect 264467 337859 264533 337864
rect 268331 337886 268397 337891
rect 263366 337789 263426 337859
rect 261894 337784 262003 337789
rect 261894 337728 261942 337784
rect 261998 337728 262003 337784
rect 261894 337726 262003 337728
rect 263366 337784 263475 337789
rect 263366 337728 263414 337784
rect 263470 337728 263475 337784
rect 263366 337726 263475 337728
rect 261937 337723 262003 337726
rect 263409 337723 263475 337726
rect 257429 337648 257722 337650
rect 257429 337592 257434 337648
rect 257490 337592 257722 337648
rect 257429 337590 257722 337592
rect 264329 337650 264395 337653
rect 264470 337650 264530 337859
rect 268331 337830 268336 337886
rect 268392 337830 268397 337886
rect 268331 337825 268397 337830
rect 264329 337648 264530 337650
rect 264329 337592 264334 337648
rect 264390 337592 264530 337648
rect 264329 337590 264530 337592
rect 268334 337650 268394 337825
rect 268469 337650 268535 337653
rect 268334 337648 268535 337650
rect 268334 337592 268474 337648
rect 268530 337592 268535 337648
rect 268334 337590 268535 337592
rect 270864 337650 270924 337893
rect 272747 337920 272813 337925
rect 272747 337864 272752 337920
rect 272808 337864 272813 337920
rect 276427 337898 276432 337954
rect 276488 337922 276493 337954
rect 279555 337954 279621 337959
rect 277623 337922 277689 337925
rect 276488 337898 276674 337922
rect 276427 337893 276674 337898
rect 272747 337859 272813 337864
rect 276430 337862 276674 337893
rect 272750 337786 272810 337859
rect 276473 337786 276539 337789
rect 272750 337784 276539 337786
rect 272750 337728 276478 337784
rect 276534 337728 276539 337784
rect 272750 337726 276539 337728
rect 276473 337723 276539 337726
rect 275277 337650 275343 337653
rect 270864 337648 275343 337650
rect 270864 337592 275282 337648
rect 275338 337592 275343 337648
rect 270864 337590 275343 337592
rect 276614 337650 276674 337862
rect 277623 337920 277962 337922
rect 277623 337864 277628 337920
rect 277684 337864 277962 337920
rect 279555 337898 279560 337954
rect 279616 337898 279621 337954
rect 280751 337956 280817 337959
rect 280751 337954 280860 337956
rect 279555 337893 279621 337898
rect 280475 337920 280541 337925
rect 277623 337862 277962 337864
rect 277623 337859 277689 337862
rect 277902 337789 277962 337862
rect 279558 337789 279618 337893
rect 280475 337864 280480 337920
rect 280536 337864 280541 337920
rect 280751 337898 280756 337954
rect 280812 337922 280860 337954
rect 283971 337922 284037 337925
rect 285765 337922 285831 337925
rect 280812 337898 280906 337922
rect 280751 337893 280906 337898
rect 280475 337859 280541 337864
rect 280800 337862 280906 337893
rect 277902 337784 278011 337789
rect 277902 337728 277950 337784
rect 278006 337728 278011 337784
rect 277902 337726 278011 337728
rect 277945 337723 278011 337726
rect 279509 337784 279618 337789
rect 279509 337728 279514 337784
rect 279570 337728 279618 337784
rect 279509 337726 279618 337728
rect 279509 337723 279575 337726
rect 279601 337650 279667 337653
rect 276614 337648 279667 337650
rect 276614 337592 279606 337648
rect 279662 337592 279667 337648
rect 276614 337590 279667 337592
rect 280478 337650 280538 337859
rect 280705 337786 280771 337789
rect 280846 337786 280906 337862
rect 283971 337920 285831 337922
rect 283971 337864 283976 337920
rect 284032 337864 285770 337920
rect 285826 337864 285831 337920
rect 283971 337862 285831 337864
rect 283971 337859 284037 337862
rect 285765 337859 285831 337862
rect 280705 337784 280906 337786
rect 280705 337728 280710 337784
rect 280766 337728 280906 337784
rect 280705 337726 280906 337728
rect 283879 337786 283945 337789
rect 284109 337786 284175 337789
rect 283879 337784 284175 337786
rect 283879 337728 283884 337784
rect 283940 337728 284114 337784
rect 284170 337728 284175 337784
rect 283879 337726 284175 337728
rect 280705 337723 280771 337726
rect 283879 337723 283945 337726
rect 284109 337723 284175 337726
rect 285581 337650 285647 337653
rect 280478 337648 285647 337650
rect 280478 337592 285586 337648
rect 285642 337592 285647 337648
rect 280478 337590 285647 337592
rect 257429 337587 257495 337590
rect 264329 337587 264395 337590
rect 268469 337587 268535 337590
rect 275277 337587 275343 337590
rect 279601 337587 279667 337590
rect 285581 337587 285647 337590
rect 253473 337512 255698 337514
rect 253473 337456 253478 337512
rect 253534 337456 255698 337512
rect 253473 337454 255698 337456
rect 253473 337451 253539 337454
rect 68921 336698 68987 336701
rect 237005 336698 237071 336701
rect 68921 336696 237071 336698
rect 68921 336640 68926 336696
rect 68982 336640 237010 336696
rect 237066 336640 237071 336696
rect 68921 336638 237071 336640
rect 68921 336635 68987 336638
rect 237005 336635 237071 336638
rect 62021 336562 62087 336565
rect 240041 336562 240107 336565
rect 62021 336560 240107 336562
rect 62021 336504 62026 336560
rect 62082 336504 240046 336560
rect 240102 336504 240107 336560
rect 62021 336502 240107 336504
rect 62021 336499 62087 336502
rect 240041 336499 240107 336502
rect 274449 336562 274515 336565
rect 290549 336562 290615 336565
rect 274449 336560 290615 336562
rect 274449 336504 274454 336560
rect 274510 336504 290554 336560
rect 290610 336504 290615 336560
rect 274449 336502 290615 336504
rect 274449 336499 274515 336502
rect 290549 336499 290615 336502
rect 53741 336426 53807 336429
rect 239489 336426 239555 336429
rect 53741 336424 239555 336426
rect 53741 336368 53746 336424
rect 53802 336368 239494 336424
rect 239550 336368 239555 336424
rect 53741 336366 239555 336368
rect 53741 336363 53807 336366
rect 239489 336363 239555 336366
rect 275461 336426 275527 336429
rect 293217 336426 293283 336429
rect 275461 336424 293283 336426
rect 275461 336368 275466 336424
rect 275522 336368 293222 336424
rect 293278 336368 293283 336424
rect 275461 336366 293283 336368
rect 275461 336363 275527 336366
rect 293217 336363 293283 336366
rect 37181 336290 37247 336293
rect 237925 336290 237991 336293
rect 37181 336288 237991 336290
rect 37181 336232 37186 336288
rect 37242 336232 237930 336288
rect 237986 336232 237991 336288
rect 37181 336230 237991 336232
rect 37181 336227 37247 336230
rect 237925 336227 237991 336230
rect 278497 336290 278563 336293
rect 286409 336290 286475 336293
rect 309777 336290 309843 336293
rect 278497 336288 278698 336290
rect 278497 336232 278502 336288
rect 278558 336232 278698 336288
rect 278497 336230 278698 336232
rect 278497 336227 278563 336230
rect 278638 336157 278698 336230
rect 286409 336288 309843 336290
rect 286409 336232 286414 336288
rect 286470 336232 309782 336288
rect 309838 336232 309843 336288
rect 286409 336230 309843 336232
rect 286409 336227 286475 336230
rect 309777 336227 309843 336230
rect 35801 336154 35867 336157
rect 237833 336154 237899 336157
rect 35801 336152 237899 336154
rect 35801 336096 35806 336152
rect 35862 336096 237838 336152
rect 237894 336096 237899 336152
rect 35801 336094 237899 336096
rect 35801 336091 35867 336094
rect 237833 336091 237899 336094
rect 276197 336154 276263 336157
rect 276933 336154 276999 336157
rect 276197 336152 276999 336154
rect 276197 336096 276202 336152
rect 276258 336096 276938 336152
rect 276994 336096 276999 336152
rect 276197 336094 276999 336096
rect 278638 336152 278747 336157
rect 278638 336096 278686 336152
rect 278742 336096 278747 336152
rect 278638 336094 278747 336096
rect 276197 336091 276263 336094
rect 276933 336091 276999 336094
rect 278681 336091 278747 336094
rect 279141 336154 279207 336157
rect 283373 336154 283439 336157
rect 279141 336152 283439 336154
rect 279141 336096 279146 336152
rect 279202 336096 283378 336152
rect 283434 336096 283439 336152
rect 279141 336094 283439 336096
rect 279141 336091 279207 336094
rect 283373 336091 283439 336094
rect 283741 336154 283807 336157
rect 319437 336154 319503 336157
rect 283741 336152 319503 336154
rect 283741 336096 283746 336152
rect 283802 336096 319442 336152
rect 319498 336096 319503 336152
rect 283741 336094 319503 336096
rect 283741 336091 283807 336094
rect 319437 336091 319503 336094
rect 28809 336018 28875 336021
rect 237373 336018 237439 336021
rect 28809 336016 237439 336018
rect 28809 335960 28814 336016
rect 28870 335960 237378 336016
rect 237434 335960 237439 336016
rect 28809 335958 237439 335960
rect 28809 335955 28875 335958
rect 237373 335955 237439 335958
rect 271781 336018 271847 336021
rect 308397 336018 308463 336021
rect 271781 336016 308463 336018
rect 271781 335960 271786 336016
rect 271842 335960 308402 336016
rect 308458 335960 308463 336016
rect 271781 335958 308463 335960
rect 271781 335955 271847 335958
rect 308397 335955 308463 335958
rect 237281 335882 237347 335885
rect 237649 335882 237715 335885
rect 243353 335882 243419 335885
rect 237281 335880 243419 335882
rect 237281 335824 237286 335880
rect 237342 335824 237654 335880
rect 237710 335824 243358 335880
rect 243414 335824 243419 335880
rect 237281 335822 243419 335824
rect 237281 335819 237347 335822
rect 237649 335819 237715 335822
rect 243353 335819 243419 335822
rect 272425 335882 272491 335885
rect 276197 335882 276263 335885
rect 272425 335880 276263 335882
rect 272425 335824 272430 335880
rect 272486 335824 276202 335880
rect 276258 335824 276263 335880
rect 272425 335822 276263 335824
rect 272425 335819 272491 335822
rect 276197 335819 276263 335822
rect 276933 335882 276999 335885
rect 283741 335882 283807 335885
rect 276933 335880 283807 335882
rect 276933 335824 276938 335880
rect 276994 335824 283746 335880
rect 283802 335824 283807 335880
rect 276933 335822 283807 335824
rect 276933 335819 276999 335822
rect 283741 335819 283807 335822
rect 236269 335746 236335 335749
rect 269113 335746 269179 335749
rect 275553 335746 275619 335749
rect 283281 335746 283347 335749
rect 284661 335746 284727 335749
rect 236269 335744 244290 335746
rect 236269 335688 236274 335744
rect 236330 335688 244290 335744
rect 236269 335686 244290 335688
rect 236269 335683 236335 335686
rect 19333 335610 19399 335613
rect 236729 335610 236795 335613
rect 19333 335608 236795 335610
rect 19333 335552 19338 335608
rect 19394 335552 236734 335608
rect 236790 335552 236795 335608
rect 19333 335550 236795 335552
rect 19333 335547 19399 335550
rect 236729 335547 236795 335550
rect 238017 335610 238083 335613
rect 239029 335610 239095 335613
rect 238017 335608 239095 335610
rect 238017 335552 238022 335608
rect 238078 335552 239034 335608
rect 239090 335552 239095 335608
rect 238017 335550 239095 335552
rect 238017 335547 238083 335550
rect 239029 335547 239095 335550
rect 11053 335474 11119 335477
rect 235533 335474 235599 335477
rect 235901 335474 235967 335477
rect 11053 335472 235967 335474
rect 11053 335416 11058 335472
rect 11114 335416 235538 335472
rect 235594 335416 235906 335472
rect 235962 335416 235967 335472
rect 11053 335414 235967 335416
rect 244230 335474 244290 335686
rect 269113 335744 270510 335746
rect 269113 335688 269118 335744
rect 269174 335688 270510 335744
rect 269113 335686 270510 335688
rect 269113 335683 269179 335686
rect 255313 335474 255379 335477
rect 244230 335472 255379 335474
rect 244230 335416 255318 335472
rect 255374 335416 255379 335472
rect 244230 335414 255379 335416
rect 270450 335474 270510 335686
rect 275553 335744 283347 335746
rect 275553 335688 275558 335744
rect 275614 335688 283286 335744
rect 283342 335688 283347 335744
rect 275553 335686 283347 335688
rect 275553 335683 275619 335686
rect 283281 335683 283347 335686
rect 283422 335744 284727 335746
rect 283422 335688 284666 335744
rect 284722 335688 284727 335744
rect 283422 335686 284727 335688
rect 283422 335613 283482 335686
rect 284661 335683 284727 335686
rect 272241 335610 272307 335613
rect 279141 335610 279207 335613
rect 272241 335608 279207 335610
rect 272241 335552 272246 335608
rect 272302 335552 279146 335608
rect 279202 335552 279207 335608
rect 272241 335550 279207 335552
rect 272241 335547 272307 335550
rect 279141 335547 279207 335550
rect 279877 335610 279943 335613
rect 282637 335610 282703 335613
rect 283005 335610 283071 335613
rect 279877 335608 281458 335610
rect 279877 335552 279882 335608
rect 279938 335552 281458 335608
rect 279877 335550 281458 335552
rect 279877 335547 279943 335550
rect 273713 335474 273779 335477
rect 270450 335472 273779 335474
rect 270450 335416 273718 335472
rect 273774 335416 273779 335472
rect 270450 335414 273779 335416
rect 11053 335411 11119 335414
rect 235533 335411 235599 335414
rect 235901 335411 235967 335414
rect 255313 335411 255379 335414
rect 273713 335411 273779 335414
rect 273989 335474 274055 335477
rect 277945 335474 278011 335477
rect 280429 335474 280495 335477
rect 273989 335472 274098 335474
rect 273989 335416 273994 335472
rect 274050 335416 274098 335472
rect 273989 335411 274098 335416
rect 277945 335472 280495 335474
rect 277945 335416 277950 335472
rect 278006 335416 280434 335472
rect 280490 335416 280495 335472
rect 277945 335414 280495 335416
rect 281398 335474 281458 335550
rect 282637 335608 283071 335610
rect 282637 335552 282642 335608
rect 282698 335552 283010 335608
rect 283066 335552 283071 335608
rect 282637 335550 283071 335552
rect 282637 335547 282703 335550
rect 283005 335547 283071 335550
rect 283373 335608 283482 335613
rect 283373 335552 283378 335608
rect 283434 335552 283482 335608
rect 283373 335550 283482 335552
rect 283373 335547 283439 335550
rect 284569 335474 284635 335477
rect 281398 335472 284635 335474
rect 281398 335416 284574 335472
rect 284630 335416 284635 335472
rect 281398 335414 284635 335416
rect 277945 335411 278011 335414
rect 280429 335411 280495 335414
rect 284569 335411 284635 335414
rect 136541 335338 136607 335341
rect 246573 335338 246639 335341
rect 136541 335336 246639 335338
rect 136541 335280 136546 335336
rect 136602 335280 246578 335336
rect 246634 335280 246639 335336
rect 136541 335278 246639 335280
rect 136541 335275 136607 335278
rect 246573 335275 246639 335278
rect 133781 335202 133847 335205
rect 246205 335202 246271 335205
rect 133781 335200 246271 335202
rect 133781 335144 133786 335200
rect 133842 335144 246210 335200
rect 246266 335144 246271 335200
rect 133781 335142 246271 335144
rect 274038 335202 274098 335411
rect 280889 335338 280955 335341
rect 543733 335338 543799 335341
rect 280889 335336 543799 335338
rect 280889 335280 280894 335336
rect 280950 335280 543738 335336
rect 543794 335280 543799 335336
rect 280889 335278 543799 335280
rect 280889 335275 280955 335278
rect 543733 335275 543799 335278
rect 274265 335202 274331 335205
rect 274038 335200 274331 335202
rect 274038 335144 274270 335200
rect 274326 335144 274331 335200
rect 274038 335142 274331 335144
rect 133781 335139 133847 335142
rect 246205 335139 246271 335142
rect 274265 335139 274331 335142
rect 281441 335202 281507 335205
rect 547873 335202 547939 335205
rect 281441 335200 547939 335202
rect 281441 335144 281446 335200
rect 281502 335144 547878 335200
rect 547934 335144 547939 335200
rect 281441 335142 547939 335144
rect 281441 335139 281507 335142
rect 547873 335139 547939 335142
rect 129641 335066 129707 335069
rect 245878 335066 245884 335068
rect 129641 335064 245884 335066
rect 129641 335008 129646 335064
rect 129702 335008 245884 335064
rect 129641 335006 245884 335008
rect 129641 335003 129707 335006
rect 245878 335004 245884 335006
rect 245948 335004 245954 335068
rect 281625 335066 281691 335069
rect 557533 335066 557599 335069
rect 281625 335064 557599 335066
rect 281625 335008 281630 335064
rect 281686 335008 557538 335064
rect 557594 335008 557599 335064
rect 281625 335006 557599 335008
rect 281625 335003 281691 335006
rect 557533 335003 557599 335006
rect 92381 334930 92447 334933
rect 238569 334930 238635 334933
rect 92381 334928 238635 334930
rect 92381 334872 92386 334928
rect 92442 334872 238574 334928
rect 238630 334872 238635 334928
rect 92381 334870 238635 334872
rect 92381 334867 92447 334870
rect 238569 334867 238635 334870
rect 282913 334930 282979 334933
rect 561673 334930 561739 334933
rect 282913 334928 561739 334930
rect 282913 334872 282918 334928
rect 282974 334872 561678 334928
rect 561734 334872 561739 334928
rect 282913 334870 561739 334872
rect 282913 334867 282979 334870
rect 561673 334867 561739 334870
rect 26233 334794 26299 334797
rect 236637 334794 236703 334797
rect 26233 334792 236703 334794
rect 26233 334736 26238 334792
rect 26294 334736 236642 334792
rect 236698 334736 236703 334792
rect 26233 334734 236703 334736
rect 26233 334731 26299 334734
rect 236637 334731 236703 334734
rect 280061 334794 280127 334797
rect 282177 334794 282243 334797
rect 280061 334792 282243 334794
rect 280061 334736 280066 334792
rect 280122 334736 282182 334792
rect 282238 334736 282243 334792
rect 280061 334734 282243 334736
rect 280061 334731 280127 334734
rect 282177 334731 282243 334734
rect 282821 334794 282887 334797
rect 564433 334794 564499 334797
rect 282821 334792 564499 334794
rect 282821 334736 282826 334792
rect 282882 334736 564438 334792
rect 564494 334736 564499 334792
rect 282821 334734 564499 334736
rect 282821 334731 282887 334734
rect 564433 334731 564499 334734
rect 16573 334658 16639 334661
rect 235901 334658 235967 334661
rect 16573 334656 235967 334658
rect 16573 334600 16578 334656
rect 16634 334600 235906 334656
rect 235962 334600 235967 334656
rect 16573 334598 235967 334600
rect 16573 334595 16639 334598
rect 235901 334595 235967 334598
rect 279417 334658 279483 334661
rect 282637 334658 282703 334661
rect 279417 334656 282703 334658
rect 279417 334600 279422 334656
rect 279478 334600 282642 334656
rect 282698 334600 282703 334656
rect 279417 334598 282703 334600
rect 279417 334595 279483 334598
rect 282637 334595 282703 334598
rect 283649 334658 283715 334661
rect 575473 334658 575539 334661
rect 283649 334656 575539 334658
rect 283649 334600 283654 334656
rect 283710 334600 575478 334656
rect 575534 334600 575539 334656
rect 283649 334598 575539 334600
rect 283649 334595 283715 334598
rect 575473 334595 575539 334598
rect 144821 334522 144887 334525
rect 247033 334522 247099 334525
rect 144821 334520 247099 334522
rect 144821 334464 144826 334520
rect 144882 334464 247038 334520
rect 247094 334464 247099 334520
rect 144821 334462 247099 334464
rect 144821 334459 144887 334462
rect 247033 334459 247099 334462
rect 279233 334522 279299 334525
rect 407757 334522 407823 334525
rect 279233 334520 407823 334522
rect 279233 334464 279238 334520
rect 279294 334464 407762 334520
rect 407818 334464 407823 334520
rect 279233 334462 407823 334464
rect 279233 334459 279299 334462
rect 407757 334459 407823 334462
rect 237925 334114 237991 334117
rect 249149 334114 249215 334117
rect 237925 334112 249215 334114
rect 237925 334056 237930 334112
rect 237986 334056 249154 334112
rect 249210 334056 249215 334112
rect 237925 334054 249215 334056
rect 237925 334051 237991 334054
rect 249149 334051 249215 334054
rect 55121 333842 55187 333845
rect 239581 333842 239647 333845
rect 55121 333840 239647 333842
rect 55121 333784 55126 333840
rect 55182 333784 239586 333840
rect 239642 333784 239647 333840
rect 55121 333782 239647 333784
rect 55121 333779 55187 333782
rect 239581 333779 239647 333782
rect 273437 333842 273503 333845
rect 409137 333842 409203 333845
rect 273437 333840 409203 333842
rect 273437 333784 273442 333840
rect 273498 333784 409142 333840
rect 409198 333784 409203 333840
rect 273437 333782 409203 333784
rect 273437 333779 273503 333782
rect 409137 333779 409203 333782
rect 52361 333706 52427 333709
rect 239213 333706 239279 333709
rect 52361 333704 239279 333706
rect 52361 333648 52366 333704
rect 52422 333648 239218 333704
rect 239274 333648 239279 333704
rect 52361 333646 239279 333648
rect 52361 333643 52427 333646
rect 239213 333643 239279 333646
rect 273345 333706 273411 333709
rect 414657 333706 414723 333709
rect 273345 333704 414723 333706
rect 273345 333648 273350 333704
rect 273406 333648 414662 333704
rect 414718 333648 414723 333704
rect 273345 333646 414723 333648
rect 273345 333643 273411 333646
rect 414657 333643 414723 333646
rect 48221 333570 48287 333573
rect 238937 333570 239003 333573
rect 48221 333568 239003 333570
rect 48221 333512 48226 333568
rect 48282 333512 238942 333568
rect 238998 333512 239003 333568
rect 48221 333510 239003 333512
rect 48221 333507 48287 333510
rect 238937 333507 239003 333510
rect 263726 333508 263732 333572
rect 263796 333570 263802 333572
rect 269113 333570 269179 333573
rect 263796 333568 269179 333570
rect 263796 333512 269118 333568
rect 269174 333512 269179 333568
rect 263796 333510 269179 333512
rect 263796 333508 263802 333510
rect 269113 333507 269179 333510
rect 274633 333570 274699 333573
rect 417417 333570 417483 333573
rect 274633 333568 417483 333570
rect 274633 333512 274638 333568
rect 274694 333512 417422 333568
rect 417478 333512 417483 333568
rect 274633 333510 417483 333512
rect 274633 333507 274699 333510
rect 417417 333507 417483 333510
rect 2681 333434 2747 333437
rect 235073 333434 235139 333437
rect 2681 333432 235139 333434
rect 2681 333376 2686 333432
rect 2742 333376 235078 333432
rect 235134 333376 235139 333432
rect 2681 333374 235139 333376
rect 2681 333371 2747 333374
rect 235073 333371 235139 333374
rect 272885 333434 272951 333437
rect 439589 333434 439655 333437
rect 272885 333432 439655 333434
rect 272885 333376 272890 333432
rect 272946 333376 439594 333432
rect 439650 333376 439655 333432
rect 272885 333374 439655 333376
rect 272885 333371 272951 333374
rect 439589 333371 439655 333374
rect 13 333298 79 333301
rect 234705 333298 234771 333301
rect 268377 333298 268443 333301
rect 13 333296 268443 333298
rect 13 333240 18 333296
rect 74 333240 234710 333296
rect 234766 333240 268382 333296
rect 268438 333240 268443 333296
rect 13 333238 268443 333240
rect 13 333235 79 333238
rect 234705 333235 234771 333238
rect 268377 333235 268443 333238
rect 283833 333298 283899 333301
rect 576853 333298 576919 333301
rect 283833 333296 576919 333298
rect 283833 333240 283838 333296
rect 283894 333240 576858 333296
rect 576914 333240 576919 333296
rect 283833 333238 576919 333240
rect 283833 333235 283899 333238
rect 576853 333235 576919 333238
rect -960 332196 480 332436
rect 277301 332210 277367 332213
rect 400857 332210 400923 332213
rect 277301 332208 400923 332210
rect 277301 332152 277306 332208
rect 277362 332152 400862 332208
rect 400918 332152 400923 332208
rect 277301 332150 400923 332152
rect 277301 332147 277367 332150
rect 400857 332147 400923 332150
rect 281533 332074 281599 332077
rect 552013 332074 552079 332077
rect 281533 332072 552079 332074
rect 281533 332016 281538 332072
rect 281594 332016 552018 332072
rect 552074 332016 552079 332072
rect 281533 332014 552079 332016
rect 281533 332011 281599 332014
rect 552013 332011 552079 332014
rect 283097 331938 283163 331941
rect 567193 331938 567259 331941
rect 283097 331936 567259 331938
rect 283097 331880 283102 331936
rect 283158 331880 567198 331936
rect 567254 331880 567259 331936
rect 283097 331878 567259 331880
rect 283097 331875 283163 331878
rect 567193 331875 567259 331878
rect 283189 331802 283255 331805
rect 571333 331802 571399 331805
rect 283189 331800 571399 331802
rect 283189 331744 283194 331800
rect 283250 331744 571338 331800
rect 571394 331744 571399 331800
rect 283189 331742 571399 331744
rect 283189 331739 283255 331742
rect 571333 331739 571399 331742
rect 284569 331394 284635 331397
rect 285029 331394 285095 331397
rect 284569 331392 285095 331394
rect 284569 331336 284574 331392
rect 284630 331336 285034 331392
rect 285090 331336 285095 331392
rect 284569 331334 285095 331336
rect 284569 331331 284635 331334
rect 285029 331331 285095 331334
rect 284661 331258 284727 331261
rect 285213 331258 285279 331261
rect 284661 331256 285279 331258
rect 284661 331200 284666 331256
rect 284722 331200 285218 331256
rect 285274 331200 285279 331256
rect 284661 331198 285279 331200
rect 284661 331195 284727 331198
rect 285213 331195 285279 331198
rect 254393 326498 254459 326501
rect 254350 326496 254459 326498
rect 254350 326440 254398 326496
rect 254454 326440 254459 326496
rect 254350 326435 254459 326440
rect 254209 326226 254275 326229
rect 254350 326226 254410 326435
rect 254209 326224 254410 326226
rect 254209 326168 254214 326224
rect 254270 326168 254410 326224
rect 254209 326166 254410 326168
rect 254209 326163 254275 326166
rect 580901 325274 580967 325277
rect 583520 325274 584960 325364
rect 580901 325272 584960 325274
rect 580901 325216 580906 325272
rect 580962 325216 584960 325272
rect 580901 325214 584960 325216
rect 580901 325211 580967 325214
rect 583520 325124 584960 325214
rect 470593 322826 470659 322829
rect 470550 322824 470659 322826
rect 470550 322768 470598 322824
rect 470654 322768 470659 322824
rect 470550 322763 470659 322768
rect 470550 322693 470610 322763
rect 470501 322688 470610 322693
rect 470501 322632 470506 322688
rect 470562 322632 470610 322688
rect 470501 322630 470610 322632
rect 470501 322627 470567 322630
rect 467833 322554 467899 322557
rect 468150 322554 468156 322556
rect 467833 322552 468156 322554
rect 467833 322496 467838 322552
rect 467894 322496 468156 322552
rect 467833 322494 468156 322496
rect 467833 322491 467899 322494
rect 468150 322492 468156 322494
rect 468220 322492 468226 322556
rect 472065 322554 472131 322557
rect 473118 322554 473124 322556
rect 472065 322552 473124 322554
rect 472065 322496 472070 322552
rect 472126 322496 473124 322552
rect 472065 322494 473124 322496
rect 472065 322491 472131 322494
rect 473118 322492 473124 322494
rect 473188 322492 473194 322556
rect 474733 322554 474799 322557
rect 475694 322554 475700 322556
rect 474733 322552 475700 322554
rect 474733 322496 474738 322552
rect 474794 322496 475700 322552
rect 474733 322494 475700 322496
rect 474733 322491 474799 322494
rect 475694 322492 475700 322494
rect 475764 322492 475770 322556
rect 478873 322554 478939 322557
rect 479190 322554 479196 322556
rect 478873 322552 479196 322554
rect 478873 322496 478878 322552
rect 478934 322496 479196 322552
rect 478873 322494 479196 322496
rect 478873 322491 478939 322494
rect 479190 322492 479196 322494
rect 479260 322492 479266 322556
rect 480253 322554 480319 322557
rect 480662 322554 480668 322556
rect 480253 322552 480668 322554
rect 480253 322496 480258 322552
rect 480314 322496 480668 322552
rect 480253 322494 480668 322496
rect 480253 322491 480319 322494
rect 480662 322492 480668 322494
rect 480732 322492 480738 322556
rect 481633 322554 481699 322557
rect 481950 322554 481956 322556
rect 481633 322552 481956 322554
rect 481633 322496 481638 322552
rect 481694 322496 481956 322552
rect 481633 322494 481956 322496
rect 481633 322491 481699 322494
rect 481950 322492 481956 322494
rect 482020 322492 482026 322556
rect 483013 322554 483079 322557
rect 483238 322554 483244 322556
rect 483013 322552 483244 322554
rect 483013 322496 483018 322552
rect 483074 322496 483244 322552
rect 483013 322494 483244 322496
rect 483013 322491 483079 322494
rect 483238 322492 483244 322494
rect 483308 322492 483314 322556
rect 486325 322554 486391 322557
rect 486918 322554 486924 322556
rect 486325 322552 486924 322554
rect 486325 322496 486330 322552
rect 486386 322496 486924 322552
rect 486325 322494 486924 322496
rect 486325 322491 486391 322494
rect 486918 322492 486924 322494
rect 486988 322492 486994 322556
rect 488533 322554 488599 322557
rect 489494 322554 489500 322556
rect 488533 322552 489500 322554
rect 488533 322496 488538 322552
rect 488594 322496 489500 322552
rect 488533 322494 489500 322496
rect 488533 322491 488599 322494
rect 489494 322492 489500 322494
rect 489564 322492 489570 322556
rect 489913 322554 489979 322557
rect 490598 322554 490604 322556
rect 489913 322552 490604 322554
rect 489913 322496 489918 322552
rect 489974 322496 490604 322552
rect 489913 322494 490604 322496
rect 489913 322491 489979 322494
rect 490598 322492 490604 322494
rect 490668 322492 490674 322556
rect 491293 322554 491359 322557
rect 496813 322556 496879 322557
rect 492254 322554 492260 322556
rect 491293 322552 492260 322554
rect 491293 322496 491298 322552
rect 491354 322496 492260 322552
rect 491293 322494 492260 322496
rect 491293 322491 491359 322494
rect 492254 322492 492260 322494
rect 492324 322492 492330 322556
rect 496813 322552 496860 322556
rect 496924 322554 496930 322556
rect 496813 322496 496818 322552
rect 496813 322492 496860 322496
rect 496924 322494 496970 322554
rect 496924 322492 496930 322494
rect 496813 322491 496879 322492
rect 519537 322420 519603 322421
rect 519486 322356 519492 322420
rect 519556 322418 519603 322420
rect 519556 322416 519648 322418
rect 519598 322360 519648 322416
rect 519556 322358 519648 322360
rect 519556 322356 519603 322358
rect 519537 322355 519603 322356
rect 469397 321604 469463 321605
rect 471973 321604 472039 321605
rect 474549 321604 474615 321605
rect 476757 321604 476823 321605
rect 478229 321604 478295 321605
rect 484393 321604 484459 321605
rect 469397 321600 469444 321604
rect 469508 321602 469514 321604
rect 469397 321544 469402 321600
rect 469397 321540 469444 321544
rect 469508 321542 469554 321602
rect 471973 321600 472020 321604
rect 472084 321602 472090 321604
rect 471973 321544 471978 321600
rect 469508 321540 469514 321542
rect 471973 321540 472020 321544
rect 472084 321542 472130 321602
rect 474549 321600 474596 321604
rect 474660 321602 474666 321604
rect 474549 321544 474554 321600
rect 472084 321540 472090 321542
rect 474549 321540 474596 321544
rect 474660 321542 474706 321602
rect 476757 321600 476804 321604
rect 476868 321602 476874 321604
rect 476757 321544 476762 321600
rect 474660 321540 474666 321542
rect 476757 321540 476804 321544
rect 476868 321542 476914 321602
rect 478229 321600 478276 321604
rect 478340 321602 478346 321604
rect 484342 321602 484348 321604
rect 478229 321544 478234 321600
rect 476868 321540 476874 321542
rect 478229 321540 478276 321544
rect 478340 321542 478386 321602
rect 484302 321542 484348 321602
rect 484412 321600 484459 321604
rect 484454 321544 484459 321600
rect 478340 321540 478346 321542
rect 484342 321540 484348 321542
rect 484412 321540 484459 321544
rect 469397 321539 469463 321540
rect 471973 321539 472039 321540
rect 474549 321539 474615 321540
rect 476757 321539 476823 321540
rect 478229 321539 478295 321540
rect 484393 321539 484459 321540
rect 485405 321604 485471 321605
rect 485405 321600 485452 321604
rect 485516 321602 485522 321604
rect 488165 321602 488231 321605
rect 492765 321602 492831 321605
rect 494237 321604 494303 321605
rect 492990 321602 492996 321604
rect 485405 321544 485410 321600
rect 485405 321540 485452 321544
rect 485516 321542 485562 321602
rect 488165 321600 488274 321602
rect 488165 321544 488170 321600
rect 488226 321544 488274 321600
rect 485516 321540 485522 321542
rect 485405 321539 485471 321540
rect 488165 321539 488274 321544
rect 492765 321600 492996 321602
rect 492765 321544 492770 321600
rect 492826 321544 492996 321600
rect 492765 321542 492996 321544
rect 492765 321539 492831 321542
rect 492990 321540 492996 321542
rect 493060 321540 493066 321604
rect 494237 321600 494284 321604
rect 494348 321602 494354 321604
rect 495525 321602 495591 321605
rect 498193 321604 498259 321605
rect 498142 321602 498148 321604
rect 494237 321544 494242 321600
rect 494237 321540 494284 321544
rect 494348 321542 494394 321602
rect 495525 321600 495634 321602
rect 495525 321544 495530 321600
rect 495586 321544 495634 321600
rect 494348 321540 494354 321542
rect 494237 321539 494303 321540
rect 495525 321539 495634 321544
rect 498102 321542 498148 321602
rect 498212 321600 498259 321604
rect 498254 321544 498259 321600
rect 498142 321540 498148 321542
rect 498212 321540 498259 321544
rect 498193 321539 498259 321540
rect 499205 321602 499271 321605
rect 500677 321604 500743 321605
rect 499205 321600 499314 321602
rect 499205 321544 499210 321600
rect 499266 321544 499314 321600
rect 499205 321539 499314 321544
rect 500677 321600 500724 321604
rect 500788 321602 500794 321604
rect 501229 321602 501295 321605
rect 503253 321604 503319 321605
rect 501822 321602 501828 321604
rect 500677 321544 500682 321600
rect 500677 321540 500724 321544
rect 500788 321542 500834 321602
rect 501229 321600 501828 321602
rect 501229 321544 501234 321600
rect 501290 321544 501828 321600
rect 501229 321542 501828 321544
rect 500788 321540 500794 321542
rect 500677 321539 500743 321540
rect 501229 321539 501295 321542
rect 501822 321540 501828 321542
rect 501892 321540 501898 321604
rect 503253 321600 503300 321604
rect 503364 321602 503370 321604
rect 503805 321602 503871 321605
rect 505461 321604 505527 321605
rect 506933 321604 506999 321605
rect 530025 321604 530091 321605
rect 504214 321602 504220 321604
rect 503253 321544 503258 321600
rect 503253 321540 503300 321544
rect 503364 321542 503410 321602
rect 503805 321600 504220 321602
rect 503805 321544 503810 321600
rect 503866 321544 504220 321600
rect 503805 321542 504220 321544
rect 503364 321540 503370 321542
rect 503253 321539 503319 321540
rect 503805 321539 503871 321542
rect 504214 321540 504220 321542
rect 504284 321540 504290 321604
rect 505461 321600 505508 321604
rect 505572 321602 505578 321604
rect 505461 321544 505466 321600
rect 505461 321540 505508 321544
rect 505572 321542 505618 321602
rect 506933 321600 506980 321604
rect 507044 321602 507050 321604
rect 529974 321602 529980 321604
rect 506933 321544 506938 321600
rect 505572 321540 505578 321542
rect 506933 321540 506980 321544
rect 507044 321542 507090 321602
rect 529934 321542 529980 321602
rect 530044 321600 530091 321604
rect 530086 321544 530091 321600
rect 507044 321540 507050 321542
rect 529974 321540 529980 321542
rect 530044 321540 530091 321544
rect 505461 321539 505527 321540
rect 506933 321539 506999 321540
rect 530025 321539 530091 321540
rect 488214 321332 488274 321539
rect 495574 321332 495634 321539
rect 499254 321332 499314 321539
rect 488206 321268 488212 321332
rect 488276 321268 488282 321332
rect 495566 321268 495572 321332
rect 495636 321268 495642 321332
rect 499246 321268 499252 321332
rect 499316 321268 499322 321332
rect 470501 319970 470567 319973
rect 470726 319970 470732 319972
rect 470456 319968 470732 319970
rect 470456 319912 470506 319968
rect 470562 319912 470732 319968
rect 470456 319910 470732 319912
rect 470501 319907 470567 319910
rect 470726 319908 470732 319910
rect 470796 319908 470802 319972
rect -960 319290 480 319380
rect 4061 319290 4127 319293
rect -960 319288 4127 319290
rect -960 319232 4066 319288
rect 4122 319232 4127 319288
rect -960 319230 4127 319232
rect -960 319140 480 319230
rect 4061 319227 4127 319230
rect 537109 316570 537175 316573
rect 536422 316568 537175 316570
rect 536422 316512 537114 316568
rect 537170 316512 537175 316568
rect 536422 316510 537175 316512
rect 536422 316500 536482 316510
rect 537109 316507 537175 316510
rect 535900 316440 536482 316500
rect 580901 312082 580967 312085
rect 583520 312082 584960 312172
rect 580901 312080 584960 312082
rect 580901 312024 580906 312080
rect 580962 312024 584960 312080
rect 580901 312022 584960 312024
rect 580901 312019 580967 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 580809 298754 580875 298757
rect 583520 298754 584960 298844
rect 580809 298752 584960 298754
rect 580809 298696 580814 298752
rect 580870 298696 584960 298752
rect 580809 298694 584960 298696
rect 580809 298691 580875 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3969 293178 4035 293181
rect -960 293176 4035 293178
rect -960 293120 3974 293176
rect 4030 293120 4035 293176
rect -960 293118 4035 293120
rect -960 293028 480 293118
rect 3969 293115 4035 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 439822 274144 440032 274204
rect 437381 274138 437447 274141
rect 439822 274138 439882 274144
rect 437381 274136 439882 274138
rect 437381 274080 437386 274136
rect 437442 274080 439882 274136
rect 437381 274078 439882 274080
rect 437381 274075 437447 274078
rect 437105 273050 437171 273053
rect 438761 273050 438827 273053
rect 437105 273048 439882 273050
rect 437105 272992 437110 273048
rect 437166 272992 438766 273048
rect 438822 272992 439882 273048
rect 437105 272990 439882 272992
rect 437105 272987 437171 272990
rect 438761 272987 438827 272990
rect 439822 272980 439882 272990
rect 439822 272920 440032 272980
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 436921 271282 436987 271285
rect 438669 271282 438735 271285
rect 436921 271280 439882 271282
rect 436921 271224 436926 271280
rect 436982 271224 438674 271280
rect 438730 271224 439882 271280
rect 436921 271222 439882 271224
rect 436921 271219 436987 271222
rect 438669 271219 438735 271222
rect 439822 271212 439882 271222
rect 439822 271152 440032 271212
rect 439822 270064 440032 270124
rect 437013 270058 437079 270061
rect 439822 270058 439882 270064
rect 437013 270056 439882 270058
rect 437013 270000 437018 270056
rect 437074 270000 439882 270056
rect 437013 269998 439882 270000
rect 437013 269995 437079 269998
rect 439822 268432 440032 268492
rect 436921 268426 436987 268429
rect 439822 268426 439882 268432
rect 436921 268424 439882 268426
rect 436921 268368 436926 268424
rect 436982 268368 439882 268424
rect 436921 268366 439882 268368
rect 436921 268363 436987 268366
rect 439822 267480 440032 267540
rect 436829 267474 436895 267477
rect 439822 267474 439882 267480
rect 436829 267472 439882 267474
rect 436829 267416 436834 267472
rect 436890 267416 439882 267472
rect 436829 267414 439882 267416
rect 436829 267411 436895 267414
rect -960 267202 480 267292
rect 3877 267202 3943 267205
rect -960 267200 3943 267202
rect -960 267144 3882 267200
rect 3938 267144 3943 267200
rect -960 267142 3943 267144
rect -960 267052 480 267142
rect 3877 267139 3943 267142
rect 439822 265712 440032 265772
rect 436737 265706 436803 265709
rect 439822 265706 439882 265712
rect 436737 265704 439882 265706
rect 436737 265648 436742 265704
rect 436798 265648 439882 265704
rect 436737 265646 439882 265648
rect 436737 265643 436803 265646
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect 535900 256600 536482 256660
rect 536422 256594 536482 256600
rect 538305 256594 538371 256597
rect 536422 256592 538371 256594
rect 536422 256536 538310 256592
rect 538366 256536 538371 256592
rect 536422 256534 538371 256536
rect 538305 256531 538371 256534
rect 535900 254968 536482 255028
rect 536422 254962 536482 254968
rect 538397 254962 538463 254965
rect 536422 254960 538463 254962
rect 536422 254904 538402 254960
rect 538458 254904 538463 254960
rect 536422 254902 538463 254904
rect 538397 254899 538463 254902
rect -960 254146 480 254236
rect 2773 254146 2839 254149
rect -960 254144 2839 254146
rect -960 254088 2778 254144
rect 2834 254088 2839 254144
rect -960 254086 2839 254088
rect -960 253996 480 254086
rect 2773 254083 2839 254086
rect 535900 253608 536482 253668
rect 536422 253602 536482 253608
rect 538489 253602 538555 253605
rect 536422 253600 538555 253602
rect 536422 253544 538494 253600
rect 538550 253544 538555 253600
rect 536422 253542 538555 253544
rect 538489 253539 538555 253542
rect 436093 247346 436159 247349
rect 436093 247344 439514 247346
rect 436093 247288 436098 247344
rect 436154 247288 439514 247344
rect 436093 247286 439514 247288
rect 436093 247283 436159 247286
rect 439454 247276 439514 247286
rect 439454 247216 440032 247276
rect 439454 245584 440032 245644
rect 436093 245578 436159 245581
rect 439454 245578 439514 245584
rect 436093 245576 439514 245578
rect 436093 245520 436098 245576
rect 436154 245520 439514 245576
rect 436093 245518 439514 245520
rect 580717 245578 580783 245581
rect 583520 245578 584960 245668
rect 580717 245576 584960 245578
rect 580717 245520 580722 245576
rect 580778 245520 584960 245576
rect 580717 245518 584960 245520
rect 436093 245515 436159 245518
rect 580717 245515 580783 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 236085 240138 236151 240141
rect 236821 240138 236887 240141
rect 236085 240136 236887 240138
rect 236085 240080 236090 240136
rect 236146 240080 236826 240136
rect 236882 240080 236887 240136
rect 236085 240078 236887 240080
rect 236085 240075 236151 240078
rect 236821 240075 236887 240078
rect 277945 239866 278011 239869
rect 502333 239866 502399 239869
rect 523125 239868 523191 239869
rect 277945 239864 502399 239866
rect 277945 239808 277950 239864
rect 278006 239808 502338 239864
rect 502394 239808 502399 239864
rect 277945 239806 502399 239808
rect 277945 239803 278011 239806
rect 502333 239803 502399 239806
rect 523096 239804 523102 239868
rect 523166 239866 523191 239868
rect 523166 239864 523258 239866
rect 523186 239808 523258 239864
rect 523166 239806 523258 239808
rect 523166 239804 523191 239806
rect 523125 239803 523191 239804
rect 279877 239730 279943 239733
rect 520273 239730 520339 239733
rect 279877 239728 520339 239730
rect 279877 239672 279882 239728
rect 279938 239672 520278 239728
rect 520334 239672 520339 239728
rect 279877 239670 520339 239672
rect 279877 239667 279943 239670
rect 520273 239667 520339 239670
rect 279417 239594 279483 239597
rect 522665 239596 522731 239597
rect 522849 239596 522915 239597
rect 522665 239594 522694 239596
rect 279417 239592 521026 239594
rect 279417 239536 279422 239592
rect 279478 239536 521026 239592
rect 279417 239534 521026 239536
rect 522602 239592 522694 239594
rect 522602 239536 522670 239592
rect 522602 239534 522694 239536
rect 279417 239531 279483 239534
rect 279509 239458 279575 239461
rect 520966 239458 521026 239534
rect 522665 239532 522694 239534
rect 522758 239532 522764 239596
rect 522824 239532 522830 239596
rect 522894 239594 522915 239596
rect 522894 239592 522986 239594
rect 522910 239536 522986 239592
rect 522894 239534 522986 239536
rect 522894 239532 522915 239534
rect 522665 239531 522731 239532
rect 522849 239531 522915 239532
rect 523217 239458 523283 239461
rect 279509 239456 509250 239458
rect 279509 239400 279514 239456
rect 279570 239400 509250 239456
rect 279509 239398 509250 239400
rect 520966 239456 523283 239458
rect 520966 239400 523222 239456
rect 523278 239400 523283 239456
rect 520966 239398 523283 239400
rect 279509 239395 279575 239398
rect 275461 239322 275527 239325
rect 484577 239322 484643 239325
rect 275461 239320 484643 239322
rect 275461 239264 275466 239320
rect 275522 239264 484582 239320
rect 484638 239264 484643 239320
rect 275461 239262 484643 239264
rect 509190 239322 509250 239398
rect 523217 239395 523283 239398
rect 527173 239322 527239 239325
rect 509190 239320 527239 239322
rect 509190 239264 527178 239320
rect 527234 239264 527239 239320
rect 509190 239262 527239 239264
rect 275461 239259 275527 239262
rect 484577 239259 484643 239262
rect 527173 239259 527239 239262
rect 256233 239186 256299 239189
rect 452101 239186 452167 239189
rect 467833 239188 467899 239189
rect 256233 239184 452026 239186
rect 256233 239128 256238 239184
rect 256294 239128 452026 239184
rect 256233 239126 452026 239128
rect 256233 239123 256299 239126
rect 237005 239050 237071 239053
rect 451966 239050 452026 239126
rect 452101 239184 456994 239186
rect 452101 239128 452106 239184
rect 452162 239128 456994 239184
rect 452101 239126 456994 239128
rect 452101 239123 452167 239126
rect 456793 239050 456859 239053
rect 237005 239048 451842 239050
rect 237005 238992 237010 239048
rect 237066 238992 451842 239048
rect 237005 238990 451842 238992
rect 451966 239048 456859 239050
rect 451966 238992 456798 239048
rect 456854 238992 456859 239048
rect 451966 238990 456859 238992
rect 456934 239050 456994 239126
rect 467782 239124 467788 239188
rect 467852 239186 467899 239188
rect 469213 239188 469279 239189
rect 469213 239186 469260 239188
rect 467852 239184 467944 239186
rect 467894 239128 467944 239184
rect 467852 239126 467944 239128
rect 469168 239184 469260 239186
rect 469168 239128 469218 239184
rect 469168 239126 469260 239128
rect 467852 239124 467899 239126
rect 467833 239123 467899 239124
rect 469213 239124 469260 239126
rect 469324 239124 469330 239188
rect 469213 239123 469279 239124
rect 480437 239052 480503 239053
rect 483013 239052 483079 239053
rect 460054 239050 460060 239052
rect 456934 238990 460060 239050
rect 237005 238987 237071 238990
rect 235441 238914 235507 238917
rect 451641 238914 451707 238917
rect 235441 238912 451707 238914
rect 235441 238856 235446 238912
rect 235502 238856 451646 238912
rect 451702 238856 451707 238912
rect 235441 238854 451707 238856
rect 451782 238914 451842 238990
rect 456793 238987 456859 238990
rect 460054 238988 460060 238990
rect 460124 238988 460130 239052
rect 480437 239050 480484 239052
rect 480392 239048 480484 239050
rect 480392 238992 480442 239048
rect 480392 238990 480484 238992
rect 480437 238988 480484 238990
rect 480548 238988 480554 239052
rect 483013 239050 483060 239052
rect 482968 239048 483060 239050
rect 482968 238992 483018 239048
rect 482968 238990 483060 238992
rect 483013 238988 483060 238990
rect 483124 238988 483130 239052
rect 480437 238987 480503 238988
rect 483013 238987 483079 238988
rect 457069 238914 457135 238917
rect 479149 238916 479215 238917
rect 494237 238916 494303 238917
rect 457846 238914 457852 238916
rect 451782 238854 456994 238914
rect 235441 238851 235507 238854
rect 451641 238851 451707 238854
rect 236821 238778 236887 238781
rect 452101 238778 452167 238781
rect 236821 238776 452167 238778
rect 236821 238720 236826 238776
rect 236882 238720 452106 238776
rect 452162 238720 452167 238776
rect 236821 238718 452167 238720
rect 236821 238715 236887 238718
rect 452101 238715 452167 238718
rect 452285 238778 452351 238781
rect 456742 238778 456748 238780
rect 452285 238776 456748 238778
rect 452285 238720 452290 238776
rect 452346 238720 456748 238776
rect 452285 238718 456748 238720
rect 452285 238715 452351 238718
rect 456742 238716 456748 238718
rect 456812 238716 456818 238780
rect 456934 238778 456994 238854
rect 457069 238912 457852 238914
rect 457069 238856 457074 238912
rect 457130 238856 457852 238912
rect 457069 238854 457852 238856
rect 457069 238851 457135 238854
rect 457846 238852 457852 238854
rect 457916 238852 457922 238916
rect 479149 238914 479196 238916
rect 479104 238912 479196 238914
rect 479104 238856 479154 238912
rect 479104 238854 479196 238856
rect 479149 238852 479196 238854
rect 479260 238852 479266 238916
rect 494237 238914 494284 238916
rect 494192 238912 494284 238914
rect 494192 238856 494242 238912
rect 494192 238854 494284 238856
rect 494237 238852 494284 238854
rect 494348 238852 494354 238916
rect 479149 238851 479215 238852
rect 494237 238851 494303 238852
rect 476757 238780 476823 238781
rect 477585 238780 477651 238781
rect 459134 238778 459140 238780
rect 456934 238718 459140 238778
rect 459134 238716 459140 238718
rect 459204 238716 459210 238780
rect 476757 238778 476804 238780
rect 476712 238776 476804 238778
rect 476712 238720 476762 238776
rect 476712 238718 476804 238720
rect 476757 238716 476804 238718
rect 476868 238716 476874 238780
rect 477534 238716 477540 238780
rect 477604 238778 477651 238780
rect 477604 238776 477696 238778
rect 477646 238720 477696 238776
rect 477604 238718 477696 238720
rect 477604 238716 477651 238718
rect 476757 238715 476823 238716
rect 477585 238715 477651 238716
rect 233049 238642 233115 238645
rect 490557 238644 490623 238645
rect 490557 238642 490604 238644
rect 233049 238640 489930 238642
rect 233049 238584 233054 238640
rect 233110 238584 489930 238640
rect 233049 238582 489930 238584
rect 490512 238640 490604 238642
rect 490512 238584 490562 238640
rect 490512 238582 490604 238584
rect 233049 238579 233115 238582
rect 232957 238506 233023 238509
rect 483657 238506 483723 238509
rect 484853 238508 484919 238509
rect 485405 238508 485471 238509
rect 487797 238508 487863 238509
rect 484853 238506 484900 238508
rect 232957 238504 483723 238506
rect 232957 238448 232962 238504
rect 233018 238448 483662 238504
rect 483718 238448 483723 238504
rect 232957 238446 483723 238448
rect 484808 238504 484900 238506
rect 484808 238448 484858 238504
rect 484808 238446 484900 238448
rect 232957 238443 233023 238446
rect 483657 238443 483723 238446
rect 484853 238444 484900 238446
rect 484964 238444 484970 238508
rect 485405 238506 485452 238508
rect 485360 238504 485452 238506
rect 485360 238448 485410 238504
rect 485360 238446 485452 238448
rect 485405 238444 485452 238446
rect 485516 238444 485522 238508
rect 487797 238506 487844 238508
rect 487752 238504 487844 238506
rect 487752 238448 487802 238504
rect 487752 238446 487844 238448
rect 487797 238444 487844 238446
rect 487908 238444 487914 238508
rect 489870 238506 489930 238582
rect 490557 238580 490604 238582
rect 490668 238580 490674 238644
rect 497590 238642 497596 238644
rect 490790 238582 497596 238642
rect 490557 238579 490623 238580
rect 490790 238506 490850 238582
rect 497590 238580 497596 238582
rect 497660 238580 497666 238644
rect 491661 238508 491727 238509
rect 491661 238506 491708 238508
rect 489870 238446 490850 238506
rect 491616 238504 491708 238506
rect 491616 238448 491666 238504
rect 491616 238446 491708 238448
rect 491661 238444 491708 238446
rect 491772 238444 491778 238508
rect 495198 238506 495204 238508
rect 492446 238446 495204 238506
rect 484853 238443 484919 238444
rect 485405 238443 485471 238444
rect 487797 238443 487863 238444
rect 491661 238443 491727 238444
rect 293401 238370 293467 238373
rect 492446 238370 492506 238446
rect 495198 238444 495204 238446
rect 495268 238444 495274 238508
rect 492765 238372 492831 238373
rect 496813 238372 496879 238373
rect 492765 238370 492812 238372
rect 293401 238368 492506 238370
rect 293401 238312 293406 238368
rect 293462 238312 492506 238368
rect 293401 238310 492506 238312
rect 492720 238368 492812 238370
rect 492720 238312 492770 238368
rect 492720 238310 492812 238312
rect 293401 238307 293467 238310
rect 492765 238308 492812 238310
rect 492876 238308 492882 238372
rect 496813 238370 496860 238372
rect 496768 238368 496860 238370
rect 496768 238312 496818 238368
rect 496768 238310 496860 238312
rect 496813 238308 496860 238310
rect 496924 238308 496930 238372
rect 492765 238307 492831 238308
rect 496813 238307 496879 238308
rect 294689 238234 294755 238237
rect 499205 238236 499271 238237
rect 496486 238234 496492 238236
rect 294689 238232 496492 238234
rect 294689 238176 294694 238232
rect 294750 238176 496492 238232
rect 294689 238174 496492 238176
rect 294689 238171 294755 238174
rect 496486 238172 496492 238174
rect 496556 238172 496562 238236
rect 499205 238234 499252 238236
rect 499160 238232 499252 238234
rect 499160 238176 499210 238232
rect 499160 238174 499252 238176
rect 499205 238172 499252 238174
rect 499316 238172 499322 238236
rect 499205 238171 499271 238172
rect 292021 238098 292087 238101
rect 470685 238100 470751 238101
rect 471789 238100 471855 238101
rect 475653 238100 475719 238101
rect 292021 238096 470610 238098
rect 292021 238040 292026 238096
rect 292082 238040 470610 238096
rect 292021 238038 470610 238040
rect 292021 238035 292087 238038
rect 232865 237962 232931 237965
rect 461577 237962 461643 237965
rect 463693 237964 463759 237965
rect 465073 237964 465139 237965
rect 463693 237962 463740 237964
rect 232865 237960 461643 237962
rect 232865 237904 232870 237960
rect 232926 237904 461582 237960
rect 461638 237904 461643 237960
rect 232865 237902 461643 237904
rect 463648 237960 463740 237962
rect 463648 237904 463698 237960
rect 463648 237902 463740 237904
rect 232865 237899 232931 237902
rect 461577 237899 461643 237902
rect 463693 237900 463740 237902
rect 463804 237900 463810 237964
rect 465022 237900 465028 237964
rect 465092 237962 465139 237964
rect 467189 237964 467255 237965
rect 468293 237964 468359 237965
rect 467189 237962 467236 237964
rect 465092 237960 465184 237962
rect 465134 237904 465184 237960
rect 465092 237902 465184 237904
rect 467144 237960 467236 237962
rect 467144 237904 467194 237960
rect 467144 237902 467236 237904
rect 465092 237900 465139 237902
rect 463693 237899 463759 237900
rect 465073 237899 465139 237900
rect 467189 237900 467236 237902
rect 467300 237900 467306 237964
rect 468293 237962 468340 237964
rect 468248 237960 468340 237962
rect 468248 237904 468298 237960
rect 468248 237902 468340 237904
rect 468293 237900 468340 237902
rect 468404 237900 468410 237964
rect 470550 237962 470610 238038
rect 470685 238096 470732 238100
rect 470796 238098 470802 238100
rect 471789 238098 471836 238100
rect 470685 238040 470690 238096
rect 470685 238036 470732 238040
rect 470796 238038 470842 238098
rect 471744 238096 471836 238098
rect 471744 238040 471794 238096
rect 471744 238038 471836 238040
rect 470796 238036 470802 238038
rect 471789 238036 471836 238038
rect 471900 238036 471906 238100
rect 475653 238098 475700 238100
rect 475608 238096 475700 238098
rect 475608 238040 475658 238096
rect 475608 238038 475700 238040
rect 475653 238036 475700 238038
rect 475764 238036 475770 238100
rect 483657 238098 483723 238101
rect 487102 238098 487108 238100
rect 483657 238096 487108 238098
rect 483657 238040 483662 238096
rect 483718 238040 487108 238096
rect 483657 238038 487108 238040
rect 470685 238035 470751 238036
rect 471789 238035 471855 238036
rect 475653 238035 475719 238036
rect 483657 238035 483723 238038
rect 487102 238036 487108 238038
rect 487172 238036 487178 238100
rect 490782 237962 490788 237964
rect 470550 237902 490788 237962
rect 490782 237900 490788 237902
rect 490852 237900 490858 237964
rect 467189 237899 467255 237900
rect 468293 237899 468359 237900
rect 292205 237826 292271 237829
rect 489310 237826 489316 237828
rect 292205 237824 489316 237826
rect 292205 237768 292210 237824
rect 292266 237768 489316 237824
rect 292205 237766 489316 237768
rect 292205 237763 292271 237766
rect 489310 237764 489316 237766
rect 489380 237764 489386 237828
rect 437197 237690 437263 237693
rect 538397 237690 538463 237693
rect 437197 237688 538463 237690
rect 437197 237632 437202 237688
rect 437258 237632 538402 237688
rect 538458 237632 538463 237688
rect 437197 237630 538463 237632
rect 437197 237627 437263 237630
rect 538397 237627 538463 237630
rect 455270 237492 455276 237556
rect 455340 237554 455346 237556
rect 459553 237554 459619 237557
rect 455340 237552 459619 237554
rect 455340 237496 459558 237552
rect 459614 237496 459619 237552
rect 455340 237494 459619 237496
rect 455340 237492 455346 237494
rect 459553 237491 459619 237494
rect 445886 237220 445892 237284
rect 445956 237282 445962 237284
rect 447041 237282 447107 237285
rect 445956 237280 447107 237282
rect 445956 237224 447046 237280
rect 447102 237224 447107 237280
rect 445956 237222 447107 237224
rect 445956 237220 445962 237222
rect 447041 237219 447107 237222
rect 460933 237282 460999 237285
rect 461342 237282 461348 237284
rect 460933 237280 461348 237282
rect 460933 237224 460938 237280
rect 460994 237224 461348 237280
rect 460933 237222 461348 237224
rect 460933 237219 460999 237222
rect 461342 237220 461348 237222
rect 461412 237220 461418 237284
rect 469213 237282 469279 237285
rect 470542 237282 470548 237284
rect 469213 237280 470548 237282
rect 469213 237224 469218 237280
rect 469274 237224 470548 237280
rect 469213 237222 470548 237224
rect 469213 237219 469279 237222
rect 470542 237220 470548 237222
rect 470612 237220 470618 237284
rect 471973 237282 472039 237285
rect 472934 237282 472940 237284
rect 471973 237280 472940 237282
rect 471973 237224 471978 237280
rect 472034 237224 472940 237280
rect 471973 237222 472940 237224
rect 471973 237219 472039 237222
rect 472934 237220 472940 237222
rect 473004 237220 473010 237284
rect 481633 237282 481699 237285
rect 481766 237282 481772 237284
rect 481633 237280 481772 237282
rect 481633 237224 481638 237280
rect 481694 237224 481772 237280
rect 481633 237222 481772 237224
rect 481633 237219 481699 237222
rect 481766 237220 481772 237222
rect 481836 237220 481842 237284
rect 481909 237282 481975 237285
rect 482318 237282 482324 237284
rect 481909 237280 482324 237282
rect 481909 237224 481914 237280
rect 481970 237224 482324 237280
rect 481909 237222 482324 237224
rect 481909 237219 481975 237222
rect 482318 237220 482324 237222
rect 482388 237220 482394 237284
rect 487153 237282 487219 237285
rect 487470 237282 487476 237284
rect 487153 237280 487476 237282
rect 487153 237224 487158 237280
rect 487214 237224 487476 237280
rect 487153 237222 487476 237224
rect 487153 237219 487219 237222
rect 487470 237220 487476 237222
rect 487540 237220 487546 237284
rect 492673 237282 492739 237285
rect 493174 237282 493180 237284
rect 492673 237280 493180 237282
rect 492673 237224 492678 237280
rect 492734 237224 493180 237280
rect 492673 237222 493180 237224
rect 492673 237219 492739 237222
rect 493174 237220 493180 237222
rect 493244 237220 493250 237284
rect 493317 237282 493383 237285
rect 493910 237282 493916 237284
rect 493317 237280 493916 237282
rect 493317 237224 493322 237280
rect 493378 237224 493916 237280
rect 493317 237222 493916 237224
rect 493317 237219 493383 237222
rect 493910 237220 493916 237222
rect 493980 237220 493986 237284
rect 495433 237282 495499 237285
rect 495934 237282 495940 237284
rect 495433 237280 495940 237282
rect 495433 237224 495438 237280
rect 495494 237224 495940 237280
rect 495433 237222 495940 237224
rect 495433 237219 495499 237222
rect 495934 237220 495940 237222
rect 496004 237220 496010 237284
rect 500953 237282 501019 237285
rect 523033 237284 523099 237285
rect 501822 237282 501828 237284
rect 500953 237280 501828 237282
rect 500953 237224 500958 237280
rect 501014 237224 501828 237280
rect 500953 237222 501828 237224
rect 500953 237219 501019 237222
rect 501822 237220 501828 237222
rect 501892 237220 501898 237284
rect 522982 237220 522988 237284
rect 523052 237282 523099 237284
rect 523052 237280 523144 237282
rect 523094 237224 523144 237280
rect 523052 237222 523144 237224
rect 523052 237220 523099 237222
rect 523033 237219 523099 237220
rect 234429 237146 234495 237149
rect 466126 237146 466132 237148
rect 234429 237144 466132 237146
rect 234429 237088 234434 237144
rect 234490 237088 466132 237144
rect 234429 237086 466132 237088
rect 234429 237083 234495 237086
rect 466126 237084 466132 237086
rect 466196 237084 466202 237148
rect 483013 237146 483079 237149
rect 483422 237146 483428 237148
rect 483013 237144 483428 237146
rect 483013 237088 483018 237144
rect 483074 237088 483428 237144
rect 483013 237086 483428 237088
rect 483013 237083 483079 237086
rect 483422 237084 483428 237086
rect 483492 237084 483498 237148
rect 488533 237146 488599 237149
rect 489126 237146 489132 237148
rect 488533 237144 489132 237146
rect 488533 237088 488538 237144
rect 488594 237088 489132 237144
rect 488533 237086 489132 237088
rect 488533 237083 488599 237086
rect 489126 237084 489132 237086
rect 489196 237084 489202 237148
rect 496813 237146 496879 237149
rect 497774 237146 497780 237148
rect 496813 237144 497780 237146
rect 496813 237088 496818 237144
rect 496874 237088 497780 237144
rect 496813 237086 497780 237088
rect 496813 237083 496879 237086
rect 497774 237084 497780 237086
rect 497844 237084 497850 237148
rect 499849 237146 499915 237149
rect 500534 237146 500540 237148
rect 499849 237144 500540 237146
rect 499849 237088 499854 237144
rect 499910 237088 500540 237144
rect 499849 237086 500540 237088
rect 499849 237083 499915 237086
rect 500534 237084 500540 237086
rect 500604 237084 500610 237148
rect 297449 237010 297515 237013
rect 506790 237010 506796 237012
rect 297449 237008 506796 237010
rect 297449 236952 297454 237008
rect 297510 236952 506796 237008
rect 297449 236950 506796 236952
rect 297449 236947 297515 236950
rect 506790 236948 506796 236950
rect 506860 236948 506866 237012
rect 299013 236874 299079 236877
rect 484393 236876 484459 236877
rect 475326 236874 475332 236876
rect 299013 236872 475332 236874
rect 299013 236816 299018 236872
rect 299074 236816 475332 236872
rect 299013 236814 475332 236816
rect 299013 236811 299079 236814
rect 475326 236812 475332 236814
rect 475396 236812 475402 236876
rect 484342 236812 484348 236876
rect 484412 236874 484459 236876
rect 491293 236876 491359 236877
rect 491293 236874 491340 236876
rect 484412 236872 484504 236874
rect 484454 236816 484504 236872
rect 484412 236814 484504 236816
rect 491248 236872 491340 236874
rect 491248 236816 491298 236872
rect 491248 236814 491340 236816
rect 484412 236812 484459 236814
rect 484393 236811 484459 236812
rect 491293 236812 491340 236814
rect 491404 236812 491410 236876
rect 491293 236811 491359 236812
rect 298829 236738 298895 236741
rect 480253 236740 480319 236741
rect 473302 236738 473308 236740
rect 298829 236736 473308 236738
rect 298829 236680 298834 236736
rect 298890 236680 473308 236736
rect 298829 236678 473308 236680
rect 298829 236675 298895 236678
rect 473302 236676 473308 236678
rect 473372 236676 473378 236740
rect 480253 236736 480300 236740
rect 480364 236738 480370 236740
rect 485773 236738 485839 236741
rect 486550 236738 486556 236740
rect 480253 236680 480258 236736
rect 480253 236676 480300 236680
rect 480364 236678 480410 236738
rect 485773 236736 486556 236738
rect 485773 236680 485778 236736
rect 485834 236680 486556 236736
rect 485773 236678 486556 236680
rect 480364 236676 480370 236678
rect 480253 236675 480319 236676
rect 485773 236675 485839 236678
rect 486550 236676 486556 236678
rect 486620 236676 486626 236740
rect 503713 236738 503779 236741
rect 504214 236738 504220 236740
rect 503713 236736 504220 236738
rect 503713 236680 503718 236736
rect 503774 236680 504220 236736
rect 503713 236678 504220 236680
rect 503713 236675 503779 236678
rect 504214 236676 504220 236678
rect 504284 236676 504290 236740
rect 439405 236602 439471 236605
rect 472065 236602 472131 236605
rect 473118 236602 473124 236604
rect 439405 236600 471898 236602
rect 439405 236544 439410 236600
rect 439466 236544 471898 236600
rect 439405 236542 471898 236544
rect 439405 236539 439471 236542
rect 446397 236466 446463 236469
rect 471838 236466 471898 236542
rect 472065 236600 473124 236602
rect 472065 236544 472070 236600
rect 472126 236544 473124 236600
rect 472065 236542 473124 236544
rect 472065 236539 472131 236542
rect 473118 236540 473124 236542
rect 473188 236540 473194 236604
rect 473445 236602 473511 236605
rect 474406 236602 474412 236604
rect 473445 236600 474412 236602
rect 473445 236544 473450 236600
rect 473506 236544 474412 236600
rect 473445 236542 474412 236544
rect 473445 236539 473511 236542
rect 474406 236540 474412 236542
rect 474476 236540 474482 236604
rect 477493 236602 477559 236605
rect 478086 236602 478092 236604
rect 477493 236600 478092 236602
rect 477493 236544 477498 236600
rect 477554 236544 478092 236600
rect 477493 236542 478092 236544
rect 477493 236539 477559 236542
rect 478086 236540 478092 236542
rect 478156 236540 478162 236604
rect 480529 236602 480595 236605
rect 480662 236602 480668 236604
rect 480529 236600 480668 236602
rect 480529 236544 480534 236600
rect 480590 236544 480668 236600
rect 480529 236542 480668 236544
rect 480529 236539 480595 236542
rect 480662 236540 480668 236542
rect 480732 236540 480738 236604
rect 476614 236466 476620 236468
rect 446397 236464 470610 236466
rect 446397 236408 446402 236464
rect 446458 236408 470610 236464
rect 446397 236406 470610 236408
rect 471838 236406 476620 236466
rect 446397 236403 446463 236406
rect 234521 236330 234587 236333
rect 469622 236330 469628 236332
rect 234521 236328 469628 236330
rect 234521 236272 234526 236328
rect 234582 236272 469628 236328
rect 234521 236270 469628 236272
rect 234521 236267 234587 236270
rect 469622 236268 469628 236270
rect 469692 236268 469698 236332
rect 470550 236194 470610 236406
rect 476614 236404 476620 236406
rect 476684 236404 476690 236468
rect 485773 236466 485839 236469
rect 485998 236466 486004 236468
rect 485773 236464 486004 236466
rect 485773 236408 485778 236464
rect 485834 236408 486004 236464
rect 485773 236406 486004 236408
rect 485773 236403 485839 236406
rect 485998 236404 486004 236406
rect 486068 236404 486074 236468
rect 471973 236332 472039 236333
rect 471973 236330 472020 236332
rect 471928 236328 472020 236330
rect 471928 236272 471978 236328
rect 471928 236270 472020 236272
rect 471973 236268 472020 236270
rect 472084 236268 472090 236332
rect 505093 236330 505159 236333
rect 505502 236330 505508 236332
rect 505093 236328 505508 236330
rect 505093 236272 505098 236328
rect 505154 236272 505508 236328
rect 505093 236270 505508 236272
rect 471973 236267 472039 236268
rect 505093 236267 505159 236270
rect 505502 236268 505508 236270
rect 505572 236268 505578 236332
rect 478822 236194 478828 236196
rect 470550 236134 478828 236194
rect 478822 236132 478828 236134
rect 478892 236132 478898 236196
rect 462405 236058 462471 236061
rect 462630 236058 462636 236060
rect 462405 236056 462636 236058
rect 462405 236000 462410 236056
rect 462466 236000 462636 236056
rect 462405 235998 462636 236000
rect 462405 235995 462471 235998
rect 462630 235996 462636 235998
rect 462700 235996 462706 236060
rect 502425 236058 502491 236061
rect 503110 236058 503116 236060
rect 502425 236056 503116 236058
rect 502425 236000 502430 236056
rect 502486 236000 503116 236056
rect 502425 235998 503116 236000
rect 502425 235995 502491 235998
rect 503110 235996 503116 235998
rect 503180 235996 503186 236060
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 579981 219058 580047 219061
rect 583520 219058 584960 219148
rect 579981 219056 584960 219058
rect 579981 219000 579986 219056
rect 580042 219000 584960 219056
rect 579981 218998 584960 219000
rect 579981 218995 580047 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3785 214978 3851 214981
rect -960 214976 3851 214978
rect -960 214920 3790 214976
rect 3846 214920 3851 214976
rect -960 214918 3851 214920
rect -960 214828 480 214918
rect 3785 214915 3851 214918
rect 580625 205730 580691 205733
rect 583520 205730 584960 205820
rect 580625 205728 584960 205730
rect 580625 205672 580630 205728
rect 580686 205672 584960 205728
rect 580625 205670 584960 205672
rect 580625 205667 580691 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 2957 201922 3023 201925
rect -960 201920 3023 201922
rect -960 201864 2962 201920
rect 3018 201864 3023 201920
rect -960 201862 3023 201864
rect -960 201772 480 201862
rect 2957 201859 3023 201862
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 2773 188866 2839 188869
rect -960 188864 2839 188866
rect -960 188808 2778 188864
rect 2834 188808 2839 188864
rect -960 188806 2839 188808
rect -960 188716 480 188806
rect 2773 188803 2839 188806
rect 579613 179210 579679 179213
rect 583520 179210 584960 179300
rect 579613 179208 584960 179210
rect 579613 179152 579618 179208
rect 579674 179152 584960 179208
rect 579613 179150 584960 179152
rect 579613 179147 579679 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580533 165882 580599 165885
rect 583520 165882 584960 165972
rect 580533 165880 584960 165882
rect 580533 165824 580538 165880
rect 580594 165824 584960 165880
rect 580533 165822 584960 165824
rect 580533 165819 580599 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3693 162890 3759 162893
rect -960 162888 3759 162890
rect -960 162832 3698 162888
rect 3754 162832 3759 162888
rect -960 162830 3759 162832
rect -960 162740 480 162830
rect 3693 162827 3759 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3141 149834 3207 149837
rect -960 149832 3207 149834
rect -960 149776 3146 149832
rect 3202 149776 3207 149832
rect -960 149774 3207 149776
rect -960 149684 480 149774
rect 3141 149771 3207 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 2773 136778 2839 136781
rect -960 136776 2839 136778
rect -960 136720 2778 136776
rect 2834 136720 2839 136776
rect -960 136718 2839 136720
rect -960 136628 480 136718
rect 2773 136715 2839 136718
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 579613 125971 579679 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3601 110666 3667 110669
rect -960 110664 3667 110666
rect -960 110608 3606 110664
rect 3662 110608 3667 110664
rect -960 110606 3667 110608
rect -960 110516 480 110606
rect 3601 110603 3667 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3233 97610 3299 97613
rect -960 97608 3299 97610
rect -960 97552 3238 97608
rect 3294 97552 3299 97608
rect -960 97550 3299 97552
rect -960 97460 480 97550
rect 3233 97547 3299 97550
rect 579613 86186 579679 86189
rect 583520 86186 584960 86276
rect 579613 86184 584960 86186
rect 579613 86128 579618 86184
rect 579674 86128 584960 86184
rect 579613 86126 584960 86128
rect 579613 86123 579679 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 2773 84690 2839 84693
rect -960 84688 2839 84690
rect -960 84632 2778 84688
rect 2834 84632 2839 84688
rect -960 84630 2839 84632
rect -960 84540 480 84630
rect 2773 84627 2839 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 580349 59666 580415 59669
rect 583520 59666 584960 59756
rect 580349 59664 584960 59666
rect 580349 59608 580354 59664
rect 580410 59608 584960 59664
rect 580349 59606 584960 59608
rect 580349 59603 580415 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2957 58578 3023 58581
rect -960 58576 3023 58578
rect -960 58520 2962 58576
rect 3018 58520 3023 58576
rect -960 58518 3023 58520
rect -960 58428 480 58518
rect 2957 58515 3023 58518
rect 580257 46338 580323 46341
rect 583520 46338 584960 46428
rect 580257 46336 584960 46338
rect 580257 46280 580262 46336
rect 580318 46280 584960 46336
rect 580257 46278 584960 46280
rect 580257 46275 580323 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2773 45522 2839 45525
rect -960 45520 2839 45522
rect -960 45464 2778 45520
rect 2834 45464 2839 45520
rect -960 45462 2839 45464
rect -960 45372 480 45462
rect 2773 45459 2839 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 2957 19410 3023 19413
rect -960 19408 3023 19410
rect -960 19352 2962 19408
rect 3018 19352 3023 19408
rect -960 19350 3023 19352
rect -960 19260 480 19350
rect 2957 19347 3023 19350
rect 284109 8938 284175 8941
rect 578601 8938 578667 8941
rect 284109 8936 578667 8938
rect 284109 8880 284114 8936
rect 284170 8880 578606 8936
rect 578662 8880 578667 8936
rect 284109 8878 578667 8880
rect 284109 8875 284175 8878
rect 578601 8875 578667 8878
rect 279969 7850 280035 7853
rect 532509 7850 532575 7853
rect 279969 7848 532575 7850
rect 279969 7792 279974 7848
rect 280030 7792 532514 7848
rect 532570 7792 532575 7848
rect 279969 7790 532575 7792
rect 279969 7787 280035 7790
rect 532509 7787 532575 7790
rect 281257 7714 281323 7717
rect 536097 7714 536163 7717
rect 281257 7712 536163 7714
rect 281257 7656 281262 7712
rect 281318 7656 536102 7712
rect 536158 7656 536163 7712
rect 281257 7654 536163 7656
rect 281257 7651 281323 7654
rect 536097 7651 536163 7654
rect 281165 7578 281231 7581
rect 539593 7578 539659 7581
rect 281165 7576 539659 7578
rect 281165 7520 281170 7576
rect 281226 7520 539598 7576
rect 539654 7520 539659 7576
rect 281165 7518 539659 7520
rect 281165 7515 281231 7518
rect 539593 7515 539659 7518
rect 93945 6626 94011 6629
rect 241697 6626 241763 6629
rect 93945 6624 241763 6626
rect -960 6490 480 6580
rect 93945 6568 93950 6624
rect 94006 6568 241702 6624
rect 241758 6568 241763 6624
rect 93945 6566 241763 6568
rect 93945 6563 94011 6566
rect 241697 6563 241763 6566
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 2773 6490 2839 6493
rect -960 6488 2839 6490
rect -960 6432 2778 6488
rect 2834 6432 2839 6488
rect -960 6430 2839 6432
rect -960 6340 480 6430
rect 2773 6427 2839 6430
rect 90357 6490 90423 6493
rect 241789 6490 241855 6493
rect 90357 6488 241855 6490
rect 90357 6432 90362 6488
rect 90418 6432 241794 6488
rect 241850 6432 241855 6488
rect 90357 6430 241855 6432
rect 90357 6427 90423 6430
rect 241789 6427 241855 6430
rect 269389 6490 269455 6493
rect 410793 6490 410859 6493
rect 269389 6488 410859 6490
rect 269389 6432 269394 6488
rect 269450 6432 410798 6488
rect 410854 6432 410859 6488
rect 583520 6476 584960 6566
rect 269389 6430 410859 6432
rect 269389 6427 269455 6430
rect 410793 6427 410859 6430
rect 86861 6354 86927 6357
rect 241881 6354 241947 6357
rect 86861 6352 241947 6354
rect 86861 6296 86866 6352
rect 86922 6296 241886 6352
rect 241942 6296 241947 6352
rect 86861 6294 241947 6296
rect 86861 6291 86927 6294
rect 241881 6291 241947 6294
rect 270217 6354 270283 6357
rect 414289 6354 414355 6357
rect 270217 6352 414355 6354
rect 270217 6296 270222 6352
rect 270278 6296 414294 6352
rect 414350 6296 414355 6352
rect 270217 6294 414355 6296
rect 270217 6291 270283 6294
rect 414289 6291 414355 6294
rect 56041 6218 56107 6221
rect 238937 6218 239003 6221
rect 56041 6216 239003 6218
rect 56041 6160 56046 6216
rect 56102 6160 238942 6216
rect 238998 6160 239003 6216
rect 56041 6158 239003 6160
rect 56041 6155 56107 6158
rect 238937 6155 239003 6158
rect 270953 6218 271019 6221
rect 428457 6218 428523 6221
rect 270953 6216 428523 6218
rect 270953 6160 270958 6216
rect 271014 6160 428462 6216
rect 428518 6160 428523 6216
rect 270953 6158 428523 6160
rect 270953 6155 271019 6158
rect 428457 6155 428523 6158
rect 137645 5266 137711 5269
rect 246481 5266 246547 5269
rect 137645 5264 246547 5266
rect 137645 5208 137650 5264
rect 137706 5208 246486 5264
rect 246542 5208 246547 5264
rect 137645 5206 246547 5208
rect 137645 5203 137711 5206
rect 246481 5203 246547 5206
rect 280429 5266 280495 5269
rect 549069 5266 549135 5269
rect 280429 5264 549135 5266
rect 280429 5208 280434 5264
rect 280490 5208 549074 5264
rect 549130 5208 549135 5264
rect 280429 5206 549135 5208
rect 280429 5203 280495 5206
rect 549069 5203 549135 5206
rect 131757 5130 131823 5133
rect 245837 5130 245903 5133
rect 131757 5128 245903 5130
rect 131757 5072 131762 5128
rect 131818 5072 245842 5128
rect 245898 5072 245903 5128
rect 131757 5070 245903 5072
rect 131757 5067 131823 5070
rect 245837 5067 245903 5070
rect 281717 5130 281783 5133
rect 559741 5130 559807 5133
rect 281717 5128 559807 5130
rect 281717 5072 281722 5128
rect 281778 5072 559746 5128
rect 559802 5072 559807 5128
rect 281717 5070 559807 5072
rect 281717 5067 281783 5070
rect 559741 5067 559807 5070
rect 128169 4994 128235 4997
rect 246573 4994 246639 4997
rect 128169 4992 246639 4994
rect 128169 4936 128174 4992
rect 128230 4936 246578 4992
rect 246634 4936 246639 4992
rect 128169 4934 246639 4936
rect 128169 4931 128235 4934
rect 246573 4931 246639 4934
rect 282545 4994 282611 4997
rect 563237 4994 563303 4997
rect 282545 4992 563303 4994
rect 282545 4936 282550 4992
rect 282606 4936 563242 4992
rect 563298 4936 563303 4992
rect 282545 4934 563303 4936
rect 282545 4931 282611 4934
rect 563237 4931 563303 4934
rect 2865 4858 2931 4861
rect 234797 4858 234863 4861
rect 2865 4856 234863 4858
rect 2865 4800 2870 4856
rect 2926 4800 234802 4856
rect 234858 4800 234863 4856
rect 2865 4798 234863 4800
rect 2865 4795 2931 4798
rect 234797 4795 234863 4798
rect 282637 4858 282703 4861
rect 566825 4858 566891 4861
rect 282637 4856 566891 4858
rect 282637 4800 282642 4856
rect 282698 4800 566830 4856
rect 566886 4800 566891 4856
rect 282637 4798 566891 4800
rect 282637 4795 282703 4798
rect 566825 4795 566891 4798
rect 234429 4722 234495 4725
rect 235717 4722 235783 4725
rect 234429 4720 235783 4722
rect 234429 4664 234434 4720
rect 234490 4664 235722 4720
rect 235778 4664 235783 4720
rect 234429 4662 235783 4664
rect 234429 4659 234495 4662
rect 235717 4659 235783 4662
rect 226241 4178 226307 4181
rect 227713 4178 227779 4181
rect 226241 4176 227779 4178
rect 226241 4120 226246 4176
rect 226302 4120 227718 4176
rect 227774 4120 227779 4176
rect 226241 4118 227779 4120
rect 226241 4115 226307 4118
rect 227713 4115 227779 4118
rect 232037 4042 232103 4045
rect 234061 4042 234127 4045
rect 232037 4040 234127 4042
rect 232037 3984 232042 4040
rect 232098 3984 234066 4040
rect 234122 3984 234127 4040
rect 232037 3982 234127 3984
rect 232037 3979 232103 3982
rect 234061 3979 234127 3982
rect 290733 3770 290799 3773
rect 472249 3770 472315 3773
rect 290733 3768 472315 3770
rect 290733 3712 290738 3768
rect 290794 3712 472254 3768
rect 472310 3712 472315 3768
rect 290733 3710 472315 3712
rect 290733 3707 290799 3710
rect 472249 3707 472315 3710
rect 290917 3634 290983 3637
rect 479333 3634 479399 3637
rect 290917 3632 479399 3634
rect 290917 3576 290922 3632
rect 290978 3576 479338 3632
rect 479394 3576 479399 3632
rect 290917 3574 479399 3576
rect 290917 3571 290983 3574
rect 479333 3571 479399 3574
rect 25313 3498 25379 3501
rect 236821 3498 236887 3501
rect 25313 3496 236887 3498
rect 25313 3440 25318 3496
rect 25374 3440 236826 3496
rect 236882 3440 236887 3496
rect 25313 3438 236887 3440
rect 25313 3435 25379 3438
rect 236821 3435 236887 3438
rect 282269 3498 282335 3501
rect 484025 3498 484091 3501
rect 282269 3496 484091 3498
rect 282269 3440 282274 3496
rect 282330 3440 484030 3496
rect 484086 3440 484091 3496
rect 282269 3438 484091 3440
rect 282269 3435 282335 3438
rect 484025 3435 484091 3438
rect 15929 3362 15995 3365
rect 236637 3362 236703 3365
rect 15929 3360 236703 3362
rect 15929 3304 15934 3360
rect 15990 3304 236642 3360
rect 236698 3304 236703 3360
rect 15929 3302 236703 3304
rect 15929 3299 15995 3302
rect 236637 3299 236703 3302
rect 309869 3362 309935 3365
rect 582189 3362 582255 3365
rect 309869 3360 582255 3362
rect 309869 3304 309874 3360
rect 309930 3304 582194 3360
rect 582250 3304 582255 3360
rect 309869 3302 582255 3304
rect 309869 3299 309935 3302
rect 582189 3299 582255 3302
<< via3 >>
rect 245884 337898 245888 337924
rect 245888 337898 245944 337924
rect 245944 337898 245948 337924
rect 245884 337860 245948 337898
rect 263732 337898 263736 337924
rect 263736 337898 263792 337924
rect 263792 337898 263796 337924
rect 263732 337860 263796 337898
rect 245884 335004 245948 335068
rect 263732 333508 263796 333572
rect 468156 322492 468220 322556
rect 473124 322492 473188 322556
rect 475700 322492 475764 322556
rect 479196 322492 479260 322556
rect 480668 322492 480732 322556
rect 481956 322492 482020 322556
rect 483244 322492 483308 322556
rect 486924 322492 486988 322556
rect 489500 322492 489564 322556
rect 490604 322492 490668 322556
rect 492260 322492 492324 322556
rect 496860 322552 496924 322556
rect 496860 322496 496874 322552
rect 496874 322496 496924 322552
rect 496860 322492 496924 322496
rect 519492 322416 519556 322420
rect 519492 322360 519542 322416
rect 519542 322360 519556 322416
rect 519492 322356 519556 322360
rect 469444 321600 469508 321604
rect 469444 321544 469458 321600
rect 469458 321544 469508 321600
rect 469444 321540 469508 321544
rect 472020 321600 472084 321604
rect 472020 321544 472034 321600
rect 472034 321544 472084 321600
rect 472020 321540 472084 321544
rect 474596 321600 474660 321604
rect 474596 321544 474610 321600
rect 474610 321544 474660 321600
rect 474596 321540 474660 321544
rect 476804 321600 476868 321604
rect 476804 321544 476818 321600
rect 476818 321544 476868 321600
rect 476804 321540 476868 321544
rect 478276 321600 478340 321604
rect 478276 321544 478290 321600
rect 478290 321544 478340 321600
rect 478276 321540 478340 321544
rect 484348 321600 484412 321604
rect 484348 321544 484398 321600
rect 484398 321544 484412 321600
rect 484348 321540 484412 321544
rect 485452 321600 485516 321604
rect 485452 321544 485466 321600
rect 485466 321544 485516 321600
rect 485452 321540 485516 321544
rect 492996 321540 493060 321604
rect 494284 321600 494348 321604
rect 494284 321544 494298 321600
rect 494298 321544 494348 321600
rect 494284 321540 494348 321544
rect 498148 321600 498212 321604
rect 498148 321544 498198 321600
rect 498198 321544 498212 321600
rect 498148 321540 498212 321544
rect 500724 321600 500788 321604
rect 500724 321544 500738 321600
rect 500738 321544 500788 321600
rect 500724 321540 500788 321544
rect 501828 321540 501892 321604
rect 503300 321600 503364 321604
rect 503300 321544 503314 321600
rect 503314 321544 503364 321600
rect 503300 321540 503364 321544
rect 504220 321540 504284 321604
rect 505508 321600 505572 321604
rect 505508 321544 505522 321600
rect 505522 321544 505572 321600
rect 505508 321540 505572 321544
rect 506980 321600 507044 321604
rect 506980 321544 506994 321600
rect 506994 321544 507044 321600
rect 506980 321540 507044 321544
rect 529980 321600 530044 321604
rect 529980 321544 530030 321600
rect 530030 321544 530044 321600
rect 529980 321540 530044 321544
rect 488212 321268 488276 321332
rect 495572 321268 495636 321332
rect 499252 321268 499316 321332
rect 470732 319908 470796 319972
rect 523102 239864 523166 239868
rect 523102 239808 523130 239864
rect 523130 239808 523166 239864
rect 523102 239804 523166 239808
rect 522694 239592 522758 239596
rect 522694 239536 522726 239592
rect 522726 239536 522758 239592
rect 522694 239532 522758 239536
rect 522830 239592 522894 239596
rect 522830 239536 522854 239592
rect 522854 239536 522894 239592
rect 522830 239532 522894 239536
rect 467788 239184 467852 239188
rect 467788 239128 467838 239184
rect 467838 239128 467852 239184
rect 467788 239124 467852 239128
rect 469260 239184 469324 239188
rect 469260 239128 469274 239184
rect 469274 239128 469324 239184
rect 469260 239124 469324 239128
rect 460060 238988 460124 239052
rect 480484 239048 480548 239052
rect 480484 238992 480498 239048
rect 480498 238992 480548 239048
rect 480484 238988 480548 238992
rect 483060 239048 483124 239052
rect 483060 238992 483074 239048
rect 483074 238992 483124 239048
rect 483060 238988 483124 238992
rect 456748 238716 456812 238780
rect 457852 238852 457916 238916
rect 479196 238912 479260 238916
rect 479196 238856 479210 238912
rect 479210 238856 479260 238912
rect 479196 238852 479260 238856
rect 494284 238912 494348 238916
rect 494284 238856 494298 238912
rect 494298 238856 494348 238912
rect 494284 238852 494348 238856
rect 459140 238716 459204 238780
rect 476804 238776 476868 238780
rect 476804 238720 476818 238776
rect 476818 238720 476868 238776
rect 476804 238716 476868 238720
rect 477540 238776 477604 238780
rect 477540 238720 477590 238776
rect 477590 238720 477604 238776
rect 477540 238716 477604 238720
rect 490604 238640 490668 238644
rect 490604 238584 490618 238640
rect 490618 238584 490668 238640
rect 484900 238504 484964 238508
rect 484900 238448 484914 238504
rect 484914 238448 484964 238504
rect 484900 238444 484964 238448
rect 485452 238504 485516 238508
rect 485452 238448 485466 238504
rect 485466 238448 485516 238504
rect 485452 238444 485516 238448
rect 487844 238504 487908 238508
rect 487844 238448 487858 238504
rect 487858 238448 487908 238504
rect 487844 238444 487908 238448
rect 490604 238580 490668 238584
rect 497596 238580 497660 238644
rect 491708 238504 491772 238508
rect 491708 238448 491722 238504
rect 491722 238448 491772 238504
rect 491708 238444 491772 238448
rect 495204 238444 495268 238508
rect 492812 238368 492876 238372
rect 492812 238312 492826 238368
rect 492826 238312 492876 238368
rect 492812 238308 492876 238312
rect 496860 238368 496924 238372
rect 496860 238312 496874 238368
rect 496874 238312 496924 238368
rect 496860 238308 496924 238312
rect 496492 238172 496556 238236
rect 499252 238232 499316 238236
rect 499252 238176 499266 238232
rect 499266 238176 499316 238232
rect 499252 238172 499316 238176
rect 463740 237960 463804 237964
rect 463740 237904 463754 237960
rect 463754 237904 463804 237960
rect 463740 237900 463804 237904
rect 465028 237960 465092 237964
rect 465028 237904 465078 237960
rect 465078 237904 465092 237960
rect 465028 237900 465092 237904
rect 467236 237960 467300 237964
rect 467236 237904 467250 237960
rect 467250 237904 467300 237960
rect 467236 237900 467300 237904
rect 468340 237960 468404 237964
rect 468340 237904 468354 237960
rect 468354 237904 468404 237960
rect 468340 237900 468404 237904
rect 470732 238096 470796 238100
rect 470732 238040 470746 238096
rect 470746 238040 470796 238096
rect 470732 238036 470796 238040
rect 471836 238096 471900 238100
rect 471836 238040 471850 238096
rect 471850 238040 471900 238096
rect 471836 238036 471900 238040
rect 475700 238096 475764 238100
rect 475700 238040 475714 238096
rect 475714 238040 475764 238096
rect 475700 238036 475764 238040
rect 487108 238036 487172 238100
rect 490788 237900 490852 237964
rect 489316 237764 489380 237828
rect 455276 237492 455340 237556
rect 445892 237220 445956 237284
rect 461348 237220 461412 237284
rect 470548 237220 470612 237284
rect 472940 237220 473004 237284
rect 481772 237220 481836 237284
rect 482324 237220 482388 237284
rect 487476 237220 487540 237284
rect 493180 237220 493244 237284
rect 493916 237220 493980 237284
rect 495940 237220 496004 237284
rect 501828 237220 501892 237284
rect 522988 237280 523052 237284
rect 522988 237224 523038 237280
rect 523038 237224 523052 237280
rect 522988 237220 523052 237224
rect 466132 237084 466196 237148
rect 483428 237084 483492 237148
rect 489132 237084 489196 237148
rect 497780 237084 497844 237148
rect 500540 237084 500604 237148
rect 506796 236948 506860 237012
rect 475332 236812 475396 236876
rect 484348 236872 484412 236876
rect 484348 236816 484398 236872
rect 484398 236816 484412 236872
rect 484348 236812 484412 236816
rect 491340 236872 491404 236876
rect 491340 236816 491354 236872
rect 491354 236816 491404 236872
rect 491340 236812 491404 236816
rect 473308 236676 473372 236740
rect 480300 236736 480364 236740
rect 480300 236680 480314 236736
rect 480314 236680 480364 236736
rect 480300 236676 480364 236680
rect 486556 236676 486620 236740
rect 504220 236676 504284 236740
rect 473124 236540 473188 236604
rect 474412 236540 474476 236604
rect 478092 236540 478156 236604
rect 480668 236540 480732 236604
rect 469628 236268 469692 236332
rect 476620 236404 476684 236468
rect 486004 236404 486068 236468
rect 472020 236328 472084 236332
rect 472020 236272 472034 236328
rect 472034 236272 472084 236328
rect 472020 236268 472084 236272
rect 505508 236268 505572 236332
rect 478828 236132 478892 236196
rect 462636 235996 462700 236060
rect 503116 235996 503180 236060
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 390000 236414 416898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 390000 240134 420618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 390000 243854 424338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 390000 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 390000 254414 398898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 390000 258134 402618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 390000 261854 406338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 390000 265574 410058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 390000 272414 416898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 390000 276134 420618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 390000 279854 424338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 390000 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 254568 381454 254888 381486
rect 254568 381218 254610 381454
rect 254846 381218 254888 381454
rect 254568 381134 254888 381218
rect 254568 380898 254610 381134
rect 254846 380898 254888 381134
rect 254568 380866 254888 380898
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 239208 363454 239528 363486
rect 239208 363218 239250 363454
rect 239486 363218 239528 363454
rect 239208 363134 239528 363218
rect 239208 362898 239250 363134
rect 239486 362898 239528 363134
rect 239208 362866 239528 362898
rect 269928 363454 270248 363486
rect 269928 363218 269970 363454
rect 270206 363218 270248 363454
rect 269928 363134 270248 363218
rect 269928 362898 269970 363134
rect 270206 362898 270248 363134
rect 269928 362866 270248 362898
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 254568 345454 254888 345486
rect 254568 345218 254610 345454
rect 254846 345218 254888 345454
rect 254568 345134 254888 345218
rect 254568 344898 254610 345134
rect 254846 344898 254888 345134
rect 254568 344866 254888 344898
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 245883 337924 245949 337925
rect 245883 337860 245884 337924
rect 245948 337860 245949 337924
rect 245883 337859 245949 337860
rect 263731 337924 263797 337925
rect 263731 337860 263732 337924
rect 263796 337860 263797 337924
rect 263731 337859 263797 337860
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 309454 236414 336000
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 313174 240134 336000
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 277174 240134 312618
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 316894 243854 336000
rect 245886 335069 245946 337859
rect 245883 335068 245949 335069
rect 245883 335004 245884 335068
rect 245948 335004 245949 335068
rect 245883 335003 245949 335004
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 320614 247574 336000
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 327454 254414 336000
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 331174 258134 336000
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 334894 261854 336000
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 263734 333573 263794 337859
rect 263731 333572 263797 333573
rect 263731 333508 263732 333572
rect 263796 333508 263797 333572
rect 263731 333507 263797 333508
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 302614 265574 336000
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 309454 272414 336000
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 313174 276134 336000
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 316894 279854 336000
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 320614 283574 336000
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 321500 438134 330618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 321500 441854 334338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 321500 445574 338058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 321500 452414 344898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 321500 456134 348618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 321500 459854 352338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 321500 463574 356058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 468155 322556 468221 322557
rect 468155 322492 468156 322556
rect 468220 322492 468221 322556
rect 468155 322491 468221 322492
rect 468158 319970 468218 322491
rect 469443 321604 469509 321605
rect 469443 321540 469444 321604
rect 469508 321540 469509 321604
rect 469443 321539 469509 321540
rect 469446 319970 469506 321539
rect 469794 321500 470414 326898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473123 322556 473189 322557
rect 473123 322492 473124 322556
rect 473188 322492 473189 322556
rect 473123 322491 473189 322492
rect 472019 321604 472085 321605
rect 472019 321540 472020 321604
rect 472084 321540 472085 321604
rect 472019 321539 472085 321540
rect 470731 319972 470797 319973
rect 470731 319970 470732 319972
rect 468158 319910 468220 319970
rect 469446 319910 469580 319970
rect 468160 319394 468220 319910
rect 469520 319394 469580 319910
rect 470608 319910 470732 319970
rect 470608 319394 470668 319910
rect 470731 319908 470732 319910
rect 470796 319908 470797 319972
rect 472022 319970 472082 321539
rect 470731 319907 470797 319908
rect 471968 319910 472082 319970
rect 473126 319970 473186 322491
rect 473514 321500 474134 330618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 475699 322556 475765 322557
rect 475699 322492 475700 322556
rect 475764 322492 475765 322556
rect 475699 322491 475765 322492
rect 474595 321604 474661 321605
rect 474595 321540 474596 321604
rect 474660 321540 474661 321604
rect 474595 321539 474661 321540
rect 474598 319970 474658 321539
rect 473126 319910 473252 319970
rect 471968 319394 472028 319910
rect 473192 319394 473252 319910
rect 474552 319910 474658 319970
rect 475702 319970 475762 322491
rect 476803 321604 476869 321605
rect 476803 321540 476804 321604
rect 476868 321540 476869 321604
rect 476803 321539 476869 321540
rect 476806 319970 476866 321539
rect 477234 321500 477854 334338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 479195 322556 479261 322557
rect 479195 322492 479196 322556
rect 479260 322492 479261 322556
rect 479195 322491 479261 322492
rect 480667 322556 480733 322557
rect 480667 322492 480668 322556
rect 480732 322492 480733 322556
rect 480667 322491 480733 322492
rect 478275 321604 478341 321605
rect 478275 321540 478276 321604
rect 478340 321540 478341 321604
rect 478275 321539 478341 321540
rect 478278 319970 478338 321539
rect 475702 319910 475836 319970
rect 476806 319910 476924 319970
rect 474552 319394 474612 319910
rect 475776 319394 475836 319910
rect 476864 319394 476924 319910
rect 478224 319910 478338 319970
rect 479198 319970 479258 322491
rect 480670 319970 480730 322491
rect 480954 321500 481574 338058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 481955 322556 482021 322557
rect 481955 322492 481956 322556
rect 482020 322492 482021 322556
rect 481955 322491 482021 322492
rect 483243 322556 483309 322557
rect 483243 322492 483244 322556
rect 483308 322492 483309 322556
rect 483243 322491 483309 322492
rect 486923 322556 486989 322557
rect 486923 322492 486924 322556
rect 486988 322492 486989 322556
rect 486923 322491 486989 322492
rect 481958 319970 482018 322491
rect 479198 319910 479372 319970
rect 480670 319910 480732 319970
rect 478224 319394 478284 319910
rect 479312 319394 479372 319910
rect 480672 319394 480732 319910
rect 481896 319910 482018 319970
rect 483246 319970 483306 322491
rect 484347 321604 484413 321605
rect 484347 321540 484348 321604
rect 484412 321540 484413 321604
rect 484347 321539 484413 321540
rect 485451 321604 485517 321605
rect 485451 321540 485452 321604
rect 485516 321540 485517 321604
rect 485451 321539 485517 321540
rect 484350 319970 484410 321539
rect 483246 319910 483316 319970
rect 481896 319394 481956 319910
rect 483256 319394 483316 319910
rect 484344 319910 484410 319970
rect 485454 319970 485514 321539
rect 486926 319970 486986 322491
rect 487794 321500 488414 344898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 489499 322556 489565 322557
rect 489499 322492 489500 322556
rect 489564 322492 489565 322556
rect 489499 322491 489565 322492
rect 490603 322556 490669 322557
rect 490603 322492 490604 322556
rect 490668 322492 490669 322556
rect 490603 322491 490669 322492
rect 488211 321332 488277 321333
rect 488211 321268 488212 321332
rect 488276 321268 488277 321332
rect 488211 321267 488277 321268
rect 488214 319970 488274 321267
rect 485454 319910 485628 319970
rect 486926 319910 486988 319970
rect 484344 319394 484404 319910
rect 485568 319394 485628 319910
rect 486928 319394 486988 319910
rect 488152 319910 488274 319970
rect 489502 319970 489562 322491
rect 490606 319970 490666 322491
rect 491514 321500 492134 348618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 492259 322556 492325 322557
rect 492259 322492 492260 322556
rect 492324 322492 492325 322556
rect 492259 322491 492325 322492
rect 492262 319970 492322 322491
rect 492995 321604 493061 321605
rect 492995 321540 492996 321604
rect 493060 321540 493061 321604
rect 492995 321539 493061 321540
rect 494283 321604 494349 321605
rect 494283 321540 494284 321604
rect 494348 321540 494349 321604
rect 494283 321539 494349 321540
rect 489502 319910 489572 319970
rect 488152 319394 488212 319910
rect 489512 319394 489572 319910
rect 490600 319910 490666 319970
rect 491960 319910 492322 319970
rect 492998 319970 493058 321539
rect 494286 319970 494346 321539
rect 495234 321500 495854 352338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 496859 322556 496925 322557
rect 496859 322492 496860 322556
rect 496924 322492 496925 322556
rect 496859 322491 496925 322492
rect 495571 321332 495637 321333
rect 495571 321268 495572 321332
rect 495636 321268 495637 321332
rect 495571 321267 495637 321268
rect 492998 319910 493108 319970
rect 490600 319394 490660 319910
rect 491960 319394 492020 319910
rect 493048 319394 493108 319910
rect 494272 319910 494346 319970
rect 495574 319970 495634 321267
rect 496862 319970 496922 322491
rect 498147 321604 498213 321605
rect 498147 321540 498148 321604
rect 498212 321540 498213 321604
rect 498147 321539 498213 321540
rect 495574 319910 495692 319970
rect 494272 319394 494332 319910
rect 495632 319394 495692 319910
rect 496856 319910 496922 319970
rect 498150 319970 498210 321539
rect 498954 321500 499574 356058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 500723 321604 500789 321605
rect 500723 321540 500724 321604
rect 500788 321540 500789 321604
rect 500723 321539 500789 321540
rect 501827 321604 501893 321605
rect 501827 321540 501828 321604
rect 501892 321540 501893 321604
rect 501827 321539 501893 321540
rect 503299 321604 503365 321605
rect 503299 321540 503300 321604
rect 503364 321540 503365 321604
rect 503299 321539 503365 321540
rect 504219 321604 504285 321605
rect 504219 321540 504220 321604
rect 504284 321540 504285 321604
rect 504219 321539 504285 321540
rect 505507 321604 505573 321605
rect 505507 321540 505508 321604
rect 505572 321540 505573 321604
rect 505507 321539 505573 321540
rect 499251 321332 499317 321333
rect 499251 321268 499252 321332
rect 499316 321268 499317 321332
rect 499251 321267 499317 321268
rect 499254 319970 499314 321267
rect 500726 319970 500786 321539
rect 498150 319910 498276 319970
rect 499254 319910 499364 319970
rect 496856 319394 496916 319910
rect 498216 319394 498276 319910
rect 499304 319394 499364 319910
rect 500664 319910 500786 319970
rect 501830 319970 501890 321539
rect 503302 319970 503362 321539
rect 501830 319910 501948 319970
rect 500664 319394 500724 319910
rect 501888 319394 501948 319910
rect 503248 319910 503362 319970
rect 504222 319970 504282 321539
rect 505510 319970 505570 321539
rect 505794 321500 506414 326898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 506979 321604 507045 321605
rect 506979 321540 506980 321604
rect 507044 321540 507045 321604
rect 506979 321539 507045 321540
rect 506982 319970 507042 321539
rect 509514 321500 510134 330618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 321500 513854 334338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 321500 517574 338058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 519491 322420 519557 322421
rect 519491 322356 519492 322420
rect 519556 322356 519557 322420
rect 519491 322355 519557 322356
rect 519494 319970 519554 322355
rect 523794 321500 524414 344898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 321500 528134 348618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 529979 321604 530045 321605
rect 529979 321540 529980 321604
rect 530044 321540 530045 321604
rect 529979 321539 530045 321540
rect 504222 319910 504396 319970
rect 505510 319910 505620 319970
rect 503248 319394 503308 319910
rect 504336 319394 504396 319910
rect 505560 319394 505620 319910
rect 506920 319910 507042 319970
rect 519432 319910 519554 319970
rect 529982 319970 530042 321539
rect 531234 321500 531854 352338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 321500 535574 356058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 529982 319910 530100 319970
rect 506920 319394 506980 319910
rect 519432 319394 519492 319910
rect 530040 319394 530100 319910
rect 440272 309454 440620 309486
rect 440272 309218 440328 309454
rect 440564 309218 440620 309454
rect 440272 309134 440620 309218
rect 440272 308898 440328 309134
rect 440564 308898 440620 309134
rect 440272 308866 440620 308898
rect 535336 309454 535684 309486
rect 535336 309218 535392 309454
rect 535628 309218 535684 309454
rect 535336 309134 535684 309218
rect 535336 308898 535392 309134
rect 535628 308898 535684 309134
rect 535336 308866 535684 308898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 440952 291454 441300 291486
rect 440952 291218 441008 291454
rect 441244 291218 441300 291454
rect 440952 291134 441300 291218
rect 440952 290898 441008 291134
rect 441244 290898 441300 291134
rect 440952 290866 441300 290898
rect 534656 291454 535004 291486
rect 534656 291218 534712 291454
rect 534948 291218 535004 291454
rect 534656 291134 535004 291218
rect 534656 290898 534712 291134
rect 534948 290898 535004 291134
rect 534656 290866 535004 290898
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 440272 273454 440620 273486
rect 440272 273218 440328 273454
rect 440564 273218 440620 273454
rect 440272 273134 440620 273218
rect 440272 272898 440328 273134
rect 440564 272898 440620 273134
rect 440272 272866 440620 272898
rect 535336 273454 535684 273486
rect 535336 273218 535392 273454
rect 535628 273218 535684 273454
rect 535336 273134 535684 273218
rect 535336 272898 535392 273134
rect 535628 272898 535684 273134
rect 535336 272866 535684 272898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 440952 255454 441300 255486
rect 440952 255218 441008 255454
rect 441244 255218 441300 255454
rect 440952 255134 441300 255218
rect 440952 254898 441008 255134
rect 441244 254898 441300 255134
rect 440952 254866 441300 254898
rect 534656 255454 535004 255486
rect 534656 255218 534712 255454
rect 534948 255218 535004 255454
rect 534656 255134 535004 255218
rect 534656 254898 534712 255134
rect 534948 254898 535004 255134
rect 534656 254866 535004 254898
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 445856 239730 445916 240040
rect 455512 239730 455572 240040
rect 445856 239670 445954 239730
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 223174 438134 238000
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 226894 441854 238000
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 230614 445574 238000
rect 445894 237285 445954 239670
rect 455278 239670 455572 239730
rect 456736 239730 456796 240040
rect 457824 239730 457884 240040
rect 459184 239730 459244 240040
rect 460136 239730 460196 240040
rect 461360 239730 461420 240040
rect 456736 239670 456810 239730
rect 457824 239670 457914 239730
rect 451794 237454 452414 238000
rect 455278 237557 455338 239670
rect 456750 238781 456810 239670
rect 457854 238917 457914 239670
rect 459142 239670 459244 239730
rect 460062 239670 460196 239730
rect 461350 239670 461420 239730
rect 462584 239730 462644 240040
rect 463672 239730 463732 240040
rect 465032 239730 465092 240040
rect 462584 239670 462698 239730
rect 463672 239670 463802 239730
rect 457851 238916 457917 238917
rect 457851 238852 457852 238916
rect 457916 238852 457917 238916
rect 457851 238851 457917 238852
rect 459142 238781 459202 239670
rect 460062 239053 460122 239670
rect 460059 239052 460125 239053
rect 460059 238988 460060 239052
rect 460124 238988 460125 239052
rect 460059 238987 460125 238988
rect 456747 238780 456813 238781
rect 456747 238716 456748 238780
rect 456812 238716 456813 238780
rect 456747 238715 456813 238716
rect 459139 238780 459205 238781
rect 459139 238716 459140 238780
rect 459204 238716 459205 238780
rect 459139 238715 459205 238716
rect 455275 237556 455341 237557
rect 455275 237492 455276 237556
rect 455340 237492 455341 237556
rect 455275 237491 455341 237492
rect 445891 237284 445957 237285
rect 445891 237220 445892 237284
rect 445956 237220 445957 237284
rect 445891 237219 445957 237220
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 205174 456134 238000
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 208894 459854 238000
rect 461350 237285 461410 239670
rect 461347 237284 461413 237285
rect 461347 237220 461348 237284
rect 461412 237220 461413 237284
rect 461347 237219 461413 237220
rect 462638 236061 462698 239670
rect 462635 236060 462701 236061
rect 462635 235996 462636 236060
rect 462700 235996 462701 236060
rect 462635 235995 462701 235996
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 212614 463574 238000
rect 463742 237965 463802 239670
rect 465030 239670 465092 239730
rect 466120 239730 466180 240040
rect 467208 239730 467268 240040
rect 467888 239730 467948 240040
rect 466120 239670 466194 239730
rect 467208 239670 467298 239730
rect 465030 237965 465090 239670
rect 463739 237964 463805 237965
rect 463739 237900 463740 237964
rect 463804 237900 463805 237964
rect 463739 237899 463805 237900
rect 465027 237964 465093 237965
rect 465027 237900 465028 237964
rect 465092 237900 465093 237964
rect 465027 237899 465093 237900
rect 466134 237149 466194 239670
rect 467238 237965 467298 239670
rect 467790 239670 467948 239730
rect 468296 239730 468356 240040
rect 469248 239730 469308 240040
rect 469656 239730 469716 240040
rect 468296 239670 468402 239730
rect 469248 239670 469322 239730
rect 467790 239189 467850 239670
rect 467787 239188 467853 239189
rect 467787 239124 467788 239188
rect 467852 239124 467853 239188
rect 467787 239123 467853 239124
rect 468342 237965 468402 239670
rect 469262 239189 469322 239670
rect 469630 239670 469716 239730
rect 470336 239730 470396 240040
rect 470744 239730 470804 240040
rect 470336 239670 470426 239730
rect 469259 239188 469325 239189
rect 469259 239124 469260 239188
rect 469324 239124 469325 239188
rect 469259 239123 469325 239124
rect 467235 237964 467301 237965
rect 467235 237900 467236 237964
rect 467300 237900 467301 237964
rect 467235 237899 467301 237900
rect 468339 237964 468405 237965
rect 468339 237900 468340 237964
rect 468404 237900 468405 237964
rect 468339 237899 468405 237900
rect 466131 237148 466197 237149
rect 466131 237084 466132 237148
rect 466196 237084 466197 237148
rect 466131 237083 466197 237084
rect 469630 236333 469690 239670
rect 470366 238770 470426 239670
rect 470734 239670 470804 239730
rect 471832 239730 471892 240040
rect 471968 239730 472028 240040
rect 473056 239730 473116 240040
rect 471832 239670 471898 239730
rect 471968 239670 472082 239730
rect 470366 238710 470610 238770
rect 469627 236332 469693 236333
rect 469627 236268 469628 236332
rect 469692 236268 469693 236332
rect 469627 236267 469693 236268
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 219454 470414 238000
rect 470550 237285 470610 238710
rect 470734 238101 470794 239670
rect 471838 238101 471898 239670
rect 470731 238100 470797 238101
rect 470731 238036 470732 238100
rect 470796 238036 470797 238100
rect 470731 238035 470797 238036
rect 471835 238100 471901 238101
rect 471835 238036 471836 238100
rect 471900 238036 471901 238100
rect 471835 238035 471901 238036
rect 470547 237284 470613 237285
rect 470547 237220 470548 237284
rect 470612 237220 470613 237284
rect 470547 237219 470613 237220
rect 472022 236333 472082 239670
rect 472942 239670 473116 239730
rect 473192 239730 473252 240040
rect 474144 239730 474204 240040
rect 474416 239730 474476 240040
rect 475504 239730 475564 240040
rect 473192 239670 473370 239730
rect 472942 237285 473002 239670
rect 473310 239050 473370 239670
rect 473126 238990 473370 239050
rect 473494 239670 474204 239730
rect 474414 239670 474476 239730
rect 475334 239670 475564 239730
rect 475640 239730 475700 240040
rect 476592 239730 476652 240040
rect 476864 239730 476924 240040
rect 477680 239730 477740 240040
rect 475640 239670 475762 239730
rect 476592 239670 476682 239730
rect 472939 237284 473005 237285
rect 472939 237220 472940 237284
rect 473004 237220 473005 237284
rect 472939 237219 473005 237220
rect 473126 236605 473186 238990
rect 473494 238770 473554 239670
rect 473310 238710 473554 238770
rect 473310 236741 473370 238710
rect 473307 236740 473373 236741
rect 473307 236676 473308 236740
rect 473372 236676 473373 236740
rect 473307 236675 473373 236676
rect 473123 236604 473189 236605
rect 473123 236540 473124 236604
rect 473188 236540 473189 236604
rect 473123 236539 473189 236540
rect 472019 236332 472085 236333
rect 472019 236268 472020 236332
rect 472084 236268 472085 236332
rect 472019 236267 472085 236268
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 223174 474134 238000
rect 474414 236605 474474 239670
rect 475334 236877 475394 239670
rect 475702 238101 475762 239670
rect 475699 238100 475765 238101
rect 475699 238036 475700 238100
rect 475764 238036 475765 238100
rect 475699 238035 475765 238036
rect 475331 236876 475397 236877
rect 475331 236812 475332 236876
rect 475396 236812 475397 236876
rect 475331 236811 475397 236812
rect 474411 236604 474477 236605
rect 474411 236540 474412 236604
rect 474476 236540 474477 236604
rect 474411 236539 474477 236540
rect 476622 236469 476682 239670
rect 476806 239670 476924 239730
rect 477542 239670 477740 239730
rect 477816 239730 477876 240040
rect 478904 239730 478964 240040
rect 479312 239730 479372 240040
rect 477816 239670 478154 239730
rect 476806 238781 476866 239670
rect 477542 238781 477602 239670
rect 476803 238780 476869 238781
rect 476803 238716 476804 238780
rect 476868 238716 476869 238780
rect 476803 238715 476869 238716
rect 477539 238780 477605 238781
rect 477539 238716 477540 238780
rect 477604 238716 477605 238780
rect 477539 238715 477605 238716
rect 476619 236468 476685 236469
rect 476619 236404 476620 236468
rect 476684 236404 476685 236468
rect 476619 236403 476685 236404
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 226894 477854 238000
rect 478094 236605 478154 239670
rect 478830 239670 478964 239730
rect 479198 239670 479372 239730
rect 480264 239730 480324 240040
rect 480672 239730 480732 240040
rect 481352 239730 481412 240040
rect 481896 239730 481956 240040
rect 482440 239730 482500 240040
rect 483120 239730 483180 240040
rect 483528 239730 483588 240040
rect 480264 239670 480362 239730
rect 478091 236604 478157 236605
rect 478091 236540 478092 236604
rect 478156 236540 478157 236604
rect 478091 236539 478157 236540
rect 478830 236197 478890 239670
rect 479198 238917 479258 239670
rect 479195 238916 479261 238917
rect 479195 238852 479196 238916
rect 479260 238852 479261 238916
rect 479195 238851 479261 238852
rect 480302 236741 480362 239670
rect 480486 239670 480732 239730
rect 481222 239670 481412 239730
rect 481774 239670 481956 239730
rect 482326 239670 482500 239730
rect 483062 239670 483180 239730
rect 483430 239670 483588 239730
rect 484344 239730 484404 240040
rect 484888 239730 484948 240040
rect 485568 239730 485628 240040
rect 484344 239670 484410 239730
rect 484888 239670 484962 239730
rect 480486 239053 480546 239670
rect 480483 239052 480549 239053
rect 480483 238988 480484 239052
rect 480548 238988 480549 239052
rect 480483 238987 480549 238988
rect 481222 238770 481282 239670
rect 480670 238710 481282 238770
rect 480299 236740 480365 236741
rect 480299 236676 480300 236740
rect 480364 236676 480365 236740
rect 480299 236675 480365 236676
rect 480670 236605 480730 238710
rect 480667 236604 480733 236605
rect 480667 236540 480668 236604
rect 480732 236540 480733 236604
rect 480667 236539 480733 236540
rect 478827 236196 478893 236197
rect 478827 236132 478828 236196
rect 478892 236132 478893 236196
rect 478827 236131 478893 236132
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 230614 481574 238000
rect 481774 237285 481834 239670
rect 482326 237285 482386 239670
rect 483062 239053 483122 239670
rect 483059 239052 483125 239053
rect 483059 238988 483060 239052
rect 483124 238988 483125 239052
rect 483059 238987 483125 238988
rect 481771 237284 481837 237285
rect 481771 237220 481772 237284
rect 481836 237220 481837 237284
rect 481771 237219 481837 237220
rect 482323 237284 482389 237285
rect 482323 237220 482324 237284
rect 482388 237220 482389 237284
rect 482323 237219 482389 237220
rect 483430 237149 483490 239670
rect 483427 237148 483493 237149
rect 483427 237084 483428 237148
rect 483492 237084 483493 237148
rect 483427 237083 483493 237084
rect 484350 236877 484410 239670
rect 484902 238509 484962 239670
rect 485454 239670 485628 239730
rect 485976 239730 486036 240040
rect 486656 239730 486716 240040
rect 485976 239670 486066 239730
rect 485454 238509 485514 239670
rect 484899 238508 484965 238509
rect 484899 238444 484900 238508
rect 484964 238444 484965 238508
rect 484899 238443 484965 238444
rect 485451 238508 485517 238509
rect 485451 238444 485452 238508
rect 485516 238444 485517 238508
rect 485451 238443 485517 238444
rect 484347 236876 484413 236877
rect 484347 236812 484348 236876
rect 484412 236812 484413 236876
rect 484347 236811 484413 236812
rect 486006 236469 486066 239670
rect 486558 239670 486716 239730
rect 487064 239730 487124 240040
rect 487880 239730 487940 240040
rect 488288 239730 488348 240040
rect 487064 239670 487170 239730
rect 486558 236741 486618 239670
rect 487110 238101 487170 239670
rect 487846 239670 487940 239730
rect 488030 239670 488348 239730
rect 489104 239730 489164 240040
rect 489376 239730 489436 240040
rect 489104 239670 489194 239730
rect 487846 238509 487906 239670
rect 487843 238508 487909 238509
rect 487843 238444 487844 238508
rect 487908 238444 487909 238508
rect 487843 238443 487909 238444
rect 488030 238370 488090 239670
rect 487478 238310 488090 238370
rect 487107 238100 487173 238101
rect 487107 238036 487108 238100
rect 487172 238036 487173 238100
rect 487107 238035 487173 238036
rect 487478 237285 487538 238310
rect 487794 237454 488414 238000
rect 487475 237284 487541 237285
rect 487475 237220 487476 237284
rect 487540 237220 487541 237284
rect 487475 237219 487541 237220
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 489134 237149 489194 239670
rect 489318 239670 489436 239730
rect 490600 239730 490660 240040
rect 490736 239730 490796 240040
rect 491416 239730 491476 240040
rect 491824 239730 491884 240040
rect 492912 239730 492972 240040
rect 493184 239730 493244 240040
rect 494000 239730 494060 240040
rect 494408 239730 494468 240040
rect 495224 239730 495284 240040
rect 490600 239670 490666 239730
rect 490736 239670 490850 239730
rect 489318 237829 489378 239670
rect 490606 238645 490666 239670
rect 490603 238644 490669 238645
rect 490603 238580 490604 238644
rect 490668 238580 490669 238644
rect 490603 238579 490669 238580
rect 490790 237965 490850 239670
rect 491342 239670 491476 239730
rect 491710 239670 491884 239730
rect 492814 239670 492972 239730
rect 493182 239670 493244 239730
rect 493918 239670 494060 239730
rect 494286 239670 494468 239730
rect 495206 239670 495284 239730
rect 495632 239730 495692 240040
rect 496584 239730 496644 240040
rect 495632 239670 496002 239730
rect 490787 237964 490853 237965
rect 490787 237900 490788 237964
rect 490852 237900 490853 237964
rect 490787 237899 490853 237900
rect 489315 237828 489381 237829
rect 489315 237764 489316 237828
rect 489380 237764 489381 237828
rect 489315 237763 489381 237764
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 489131 237148 489197 237149
rect 489131 237084 489132 237148
rect 489196 237084 489197 237148
rect 489131 237083 489197 237084
rect 486555 236740 486621 236741
rect 486555 236676 486556 236740
rect 486620 236676 486621 236740
rect 486555 236675 486621 236676
rect 486003 236468 486069 236469
rect 486003 236404 486004 236468
rect 486068 236404 486069 236468
rect 486003 236403 486069 236404
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 201454 488414 236898
rect 491342 236877 491402 239670
rect 491710 238509 491770 239670
rect 491707 238508 491773 238509
rect 491707 238444 491708 238508
rect 491772 238444 491773 238508
rect 491707 238443 491773 238444
rect 492814 238373 492874 239670
rect 492811 238372 492877 238373
rect 492811 238308 492812 238372
rect 492876 238308 492877 238372
rect 492811 238307 492877 238308
rect 491339 236876 491405 236877
rect 491339 236812 491340 236876
rect 491404 236812 491405 236876
rect 491339 236811 491405 236812
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 205174 492134 238000
rect 493182 237285 493242 239670
rect 493918 237285 493978 239670
rect 494286 238917 494346 239670
rect 494283 238916 494349 238917
rect 494283 238852 494284 238916
rect 494348 238852 494349 238916
rect 494283 238851 494349 238852
rect 495206 238509 495266 239670
rect 495203 238508 495269 238509
rect 495203 238444 495204 238508
rect 495268 238444 495269 238508
rect 495203 238443 495269 238444
rect 493179 237284 493245 237285
rect 493179 237220 493180 237284
rect 493244 237220 493245 237284
rect 493179 237219 493245 237220
rect 493915 237284 493981 237285
rect 493915 237220 493916 237284
rect 493980 237220 493981 237284
rect 493915 237219 493981 237220
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 208894 495854 238000
rect 495942 237285 496002 239670
rect 496494 239670 496644 239730
rect 496856 239730 496916 240040
rect 497672 239730 497732 240040
rect 496856 239670 496922 239730
rect 496494 238237 496554 239670
rect 496862 238373 496922 239670
rect 497598 239670 497732 239730
rect 497598 238645 497658 239670
rect 497808 239050 497868 240040
rect 499304 239730 499364 240040
rect 497782 238990 497868 239050
rect 499254 239670 499364 239730
rect 500528 239730 500588 240040
rect 501888 239730 501948 240040
rect 500528 239670 500602 239730
rect 497595 238644 497661 238645
rect 497595 238580 497596 238644
rect 497660 238580 497661 238644
rect 497595 238579 497661 238580
rect 496859 238372 496925 238373
rect 496859 238308 496860 238372
rect 496924 238308 496925 238372
rect 496859 238307 496925 238308
rect 496491 238236 496557 238237
rect 496491 238172 496492 238236
rect 496556 238172 496557 238236
rect 496491 238171 496557 238172
rect 495939 237284 496005 237285
rect 495939 237220 495940 237284
rect 496004 237220 496005 237284
rect 495939 237219 496005 237220
rect 497782 237149 497842 238990
rect 499254 238237 499314 239670
rect 499251 238236 499317 238237
rect 499251 238172 499252 238236
rect 499316 238172 499317 238236
rect 499251 238171 499317 238172
rect 497779 237148 497845 237149
rect 497779 237084 497780 237148
rect 497844 237084 497845 237148
rect 497779 237083 497845 237084
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 212614 499574 238000
rect 500542 237149 500602 239670
rect 501830 239670 501948 239730
rect 503112 239730 503172 240040
rect 504336 239730 504396 240040
rect 505560 239730 505620 240040
rect 503112 239670 503178 239730
rect 501830 237285 501890 239670
rect 501827 237284 501893 237285
rect 501827 237220 501828 237284
rect 501892 237220 501893 237284
rect 501827 237219 501893 237220
rect 500539 237148 500605 237149
rect 500539 237084 500540 237148
rect 500604 237084 500605 237148
rect 500539 237083 500605 237084
rect 503118 236061 503178 239670
rect 504222 239670 504396 239730
rect 505510 239670 505620 239730
rect 506784 239730 506844 240040
rect 506784 239670 506858 239730
rect 504222 236741 504282 239670
rect 504219 236740 504285 236741
rect 504219 236676 504220 236740
rect 504284 236676 504285 236740
rect 504219 236675 504285 236676
rect 505510 236333 505570 239670
rect 505507 236332 505573 236333
rect 505507 236268 505508 236332
rect 505572 236268 505573 236332
rect 505507 236267 505573 236268
rect 503115 236060 503181 236061
rect 503115 235996 503116 236060
rect 503180 235996 503181 236060
rect 503115 235995 503181 235996
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 219454 506414 238000
rect 506798 237013 506858 239670
rect 522696 239597 522756 240040
rect 522832 239597 522892 240040
rect 522968 239730 523028 240040
rect 523104 239869 523164 240040
rect 523101 239868 523167 239869
rect 523101 239804 523102 239868
rect 523166 239804 523167 239868
rect 523101 239803 523167 239804
rect 522968 239670 523050 239730
rect 522693 239596 522759 239597
rect 522693 239532 522694 239596
rect 522758 239532 522759 239596
rect 522693 239531 522759 239532
rect 522829 239596 522895 239597
rect 522829 239532 522830 239596
rect 522894 239532 522895 239596
rect 522829 239531 522895 239532
rect 506795 237012 506861 237013
rect 506795 236948 506796 237012
rect 506860 236948 506861 237012
rect 506795 236947 506861 236948
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 223174 510134 238000
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 226894 513854 238000
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 230614 517574 238000
rect 522990 237285 523050 239670
rect 523794 237454 524414 238000
rect 522987 237284 523053 237285
rect 522987 237220 522988 237284
rect 523052 237220 523053 237284
rect 522987 237219 523053 237220
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 205174 528134 238000
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 208894 531854 238000
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 212614 535574 238000
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 254610 381218 254846 381454
rect 254610 380898 254846 381134
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 239250 363218 239486 363454
rect 239250 362898 239486 363134
rect 269970 363218 270206 363454
rect 269970 362898 270206 363134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 254610 345218 254846 345454
rect 254610 344898 254846 345134
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 440328 309218 440564 309454
rect 440328 308898 440564 309134
rect 535392 309218 535628 309454
rect 535392 308898 535628 309134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 441008 291218 441244 291454
rect 441008 290898 441244 291134
rect 534712 291218 534948 291454
rect 534712 290898 534948 291134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 440328 273218 440564 273454
rect 440328 272898 440564 273134
rect 535392 273218 535628 273454
rect 535392 272898 535628 273134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 441008 255218 441244 255454
rect 441008 254898 441244 255134
rect 534712 255218 534948 255454
rect 534712 254898 534948 255134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 254610 381454
rect 254846 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 254610 381134
rect 254846 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 239250 363454
rect 239486 363218 269970 363454
rect 270206 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 239250 363134
rect 239486 362898 269970 363134
rect 270206 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 254610 345454
rect 254846 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 254610 345134
rect 254846 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 440328 309454
rect 440564 309218 535392 309454
rect 535628 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 440328 309134
rect 440564 308898 535392 309134
rect 535628 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 441008 291454
rect 441244 291218 534712 291454
rect 534948 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 441008 291134
rect 441244 290898 534712 291134
rect 534948 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 440328 273454
rect 440564 273218 535392 273454
rect 535628 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 440328 273134
rect 440564 272898 535392 273134
rect 535628 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 441008 255454
rect 441244 255218 534712 255454
rect 534948 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 441008 255134
rect 441244 254898 534712 255134
rect 534948 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 1636725598
transform 1 0 235000 0 1 338000
box 0 0 50000 50000
use sky130_sram_1kbyte_1rw1r_32x256_8  SRAM0
timestamp 1636725598
transform 1 0 440000 0 1 240000
box 0 0 95956 79500
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 336000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 390000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 321500 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 321500 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 336000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 390000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 321500 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 321500 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 321500 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 336000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 390000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 321500 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 321500 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 321500 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 336000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 390000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 321500 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 321500 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 321500 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 336000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 336000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 390000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 390000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 321500 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 321500 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 321500 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 336000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 336000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 390000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 390000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 321500 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 321500 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 321500 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 336000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 336000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 390000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 390000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 321500 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 321500 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 321500 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 336000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 336000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 390000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 390000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 321500 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 321500 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 321500 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
