magic
tech sky130A
magscale 1 2
timestamp 1636725486
<< locali >>
rect 32137 46427 32171 46597
rect 28457 45815 28491 45917
rect 30205 45339 30239 45509
rect 30297 44863 30331 44965
rect 9965 44319 9999 44489
rect 17969 44183 18003 44489
rect 12725 43639 12759 43945
rect 24133 42075 24167 42245
rect 48973 12223 49007 31841
rect 49065 9503 49099 30005
rect 673 3315 707 7361
rect 765 4675 799 6069
rect 857 2975 891 7225
rect 949 3995 983 7293
rect 46121 5695 46155 5797
rect 9873 5083 9907 5185
rect 48973 4131 49007 6613
rect 41889 3519 41923 3689
rect 949 2635 983 3417
rect 6319 3009 6411 3043
rect 6377 2839 6411 3009
rect 8769 2431 8803 2533
rect 7389 1343 7423 1649
rect 8861 935 8895 1853
<< viali >>
rect 1501 47209 1535 47243
rect 2329 47209 2363 47243
rect 3985 47209 4019 47243
rect 4629 47209 4663 47243
rect 5365 47209 5399 47243
rect 6561 47209 6595 47243
rect 7205 47209 7239 47243
rect 8309 47209 8343 47243
rect 9505 47209 9539 47243
rect 10885 47209 10919 47243
rect 11989 47209 12023 47243
rect 13369 47209 13403 47243
rect 14565 47209 14599 47243
rect 15853 47209 15887 47243
rect 17049 47209 17083 47243
rect 18245 47209 18279 47243
rect 19533 47209 19567 47243
rect 20821 47209 20855 47243
rect 22109 47209 22143 47243
rect 23305 47209 23339 47243
rect 24593 47209 24627 47243
rect 25881 47209 25915 47243
rect 27169 47209 27203 47243
rect 28365 47209 28399 47243
rect 29745 47209 29779 47243
rect 30849 47209 30883 47243
rect 32229 47209 32263 47243
rect 33241 47209 33275 47243
rect 34069 47209 34103 47243
rect 34897 47209 34931 47243
rect 35817 47209 35851 47243
rect 38209 47209 38243 47243
rect 39037 47209 39071 47243
rect 40049 47209 40083 47243
rect 40693 47209 40727 47243
rect 42625 47209 42659 47243
rect 43361 47209 43395 47243
rect 44373 47209 44407 47243
rect 45477 47209 45511 47243
rect 46213 47209 46247 47243
rect 48053 47209 48087 47243
rect 46949 47141 46983 47175
rect 1685 47005 1719 47039
rect 2145 47005 2179 47039
rect 2881 47005 2915 47039
rect 3801 47005 3835 47039
rect 4813 47005 4847 47039
rect 5549 47005 5583 47039
rect 6377 47005 6411 47039
rect 7389 47005 7423 47039
rect 8125 47005 8159 47039
rect 9689 47005 9723 47039
rect 10701 47005 10735 47039
rect 12173 47005 12207 47039
rect 13185 47005 13219 47039
rect 14381 47005 14415 47039
rect 15669 47005 15703 47039
rect 17233 47005 17267 47039
rect 18429 47005 18463 47039
rect 19717 47005 19751 47039
rect 20637 47005 20671 47039
rect 21925 47005 21959 47039
rect 23121 47005 23155 47039
rect 24409 47005 24443 47039
rect 25697 47005 25731 47039
rect 26985 47005 27019 47039
rect 28181 47005 28215 47039
rect 29561 47005 29595 47039
rect 30665 47005 30699 47039
rect 32413 47005 32447 47039
rect 33425 47005 33459 47039
rect 33885 47005 33919 47039
rect 34713 47005 34747 47039
rect 35633 47005 35667 47039
rect 36369 47005 36403 47039
rect 37565 47005 37599 47039
rect 38393 47005 38427 47039
rect 38853 47005 38887 47039
rect 39865 47005 39899 47039
rect 40877 47005 40911 47039
rect 41337 47005 41371 47039
rect 42441 47005 42475 47039
rect 43177 47005 43211 47039
rect 44189 47005 44223 47039
rect 45293 47005 45327 47039
rect 46029 47005 46063 47039
rect 46765 47005 46799 47039
rect 47869 47005 47903 47039
rect 10241 46937 10275 46971
rect 12633 46937 12667 46971
rect 15209 46937 15243 46971
rect 3065 46869 3099 46903
rect 28917 46869 28951 46903
rect 31401 46869 31435 46903
rect 36553 46869 36587 46903
rect 37381 46869 37415 46903
rect 41521 46869 41555 46903
rect 1501 46665 1535 46699
rect 2421 46665 2455 46699
rect 4353 46665 4387 46699
rect 4905 46665 4939 46699
rect 5733 46665 5767 46699
rect 7389 46665 7423 46699
rect 8769 46665 8803 46699
rect 9965 46665 9999 46699
rect 10793 46665 10827 46699
rect 12265 46665 12299 46699
rect 13001 46665 13035 46699
rect 13645 46665 13679 46699
rect 14933 46665 14967 46699
rect 15945 46665 15979 46699
rect 18153 46665 18187 46699
rect 18889 46665 18923 46699
rect 19993 46665 20027 46699
rect 20545 46665 20579 46699
rect 22017 46665 22051 46699
rect 22753 46665 22787 46699
rect 24317 46665 24351 46699
rect 25053 46665 25087 46699
rect 26157 46665 26191 46699
rect 28273 46665 28307 46699
rect 30021 46665 30055 46699
rect 33057 46665 33091 46699
rect 33701 46665 33735 46699
rect 34529 46665 34563 46699
rect 36185 46665 36219 46699
rect 37473 46665 37507 46699
rect 38025 46665 38059 46699
rect 38669 46665 38703 46699
rect 39957 46665 39991 46699
rect 42625 46665 42659 46699
rect 43729 46665 43763 46699
rect 44741 46665 44775 46699
rect 45477 46665 45511 46699
rect 46213 46665 46247 46699
rect 46949 46665 46983 46699
rect 32137 46597 32171 46631
rect 1685 46529 1719 46563
rect 2605 46529 2639 46563
rect 3433 46529 3467 46563
rect 4169 46529 4203 46563
rect 5089 46529 5123 46563
rect 5549 46529 5583 46563
rect 6377 46529 6411 46563
rect 7573 46529 7607 46563
rect 8585 46529 8619 46563
rect 10149 46529 10183 46563
rect 10977 46529 11011 46563
rect 12081 46529 12115 46563
rect 12817 46529 12851 46563
rect 13829 46529 13863 46563
rect 15117 46529 15151 46563
rect 16129 46529 16163 46563
rect 17325 46529 17359 46563
rect 17969 46529 18003 46563
rect 18705 46529 18739 46563
rect 19809 46529 19843 46563
rect 20729 46529 20763 46563
rect 21833 46529 21867 46563
rect 22569 46529 22603 46563
rect 23489 46529 23523 46563
rect 24133 46529 24167 46563
rect 24869 46529 24903 46563
rect 26341 46529 26375 46563
rect 27445 46529 27479 46563
rect 28089 46529 28123 46563
rect 28917 46529 28951 46563
rect 29837 46529 29871 46563
rect 31125 46529 31159 46563
rect 21281 46461 21315 46495
rect 27629 46461 27663 46495
rect 32321 46529 32355 46563
rect 33241 46529 33275 46563
rect 33885 46529 33919 46563
rect 34345 46529 34379 46563
rect 35081 46529 35115 46563
rect 36369 46529 36403 46563
rect 37289 46529 37323 46563
rect 38209 46529 38243 46563
rect 38853 46529 38887 46563
rect 39773 46529 39807 46563
rect 40509 46529 40543 46563
rect 41337 46529 41371 46563
rect 41797 46529 41831 46563
rect 42441 46529 42475 46563
rect 43545 46529 43579 46563
rect 44557 46529 44591 46563
rect 45293 46529 45327 46563
rect 46029 46529 46063 46563
rect 46765 46529 46799 46563
rect 47869 46529 47903 46563
rect 6561 46393 6595 46427
rect 17509 46393 17543 46427
rect 32137 46393 32171 46427
rect 32505 46393 32539 46427
rect 35265 46393 35299 46427
rect 41153 46393 41187 46427
rect 48053 46393 48087 46427
rect 3617 46325 3651 46359
rect 8125 46325 8159 46359
rect 9413 46325 9447 46359
rect 11529 46325 11563 46359
rect 14289 46325 14323 46359
rect 16681 46325 16715 46359
rect 23581 46325 23615 46359
rect 29009 46325 29043 46359
rect 31217 46325 31251 46359
rect 40693 46325 40727 46359
rect 1961 46121 1995 46155
rect 2605 46121 2639 46155
rect 3801 46121 3835 46155
rect 8217 46121 8251 46155
rect 12449 46121 12483 46155
rect 12909 46121 12943 46155
rect 17785 46121 17819 46155
rect 18429 46121 18463 46155
rect 20545 46121 20579 46155
rect 21741 46121 21775 46155
rect 26893 46121 26927 46155
rect 27997 46121 28031 46155
rect 28733 46121 28767 46155
rect 29561 46121 29595 46155
rect 30573 46121 30607 46155
rect 31217 46121 31251 46155
rect 35541 46121 35575 46155
rect 39313 46121 39347 46155
rect 40969 46121 41003 46155
rect 41889 46121 41923 46155
rect 43085 46121 43119 46155
rect 44281 46121 44315 46155
rect 45845 46121 45879 46155
rect 46581 46121 46615 46155
rect 47317 46121 47351 46155
rect 19901 46053 19935 46087
rect 40049 46053 40083 46087
rect 45201 46053 45235 46087
rect 1501 45985 1535 46019
rect 8953 45985 8987 46019
rect 2145 45917 2179 45951
rect 2789 45917 2823 45951
rect 3985 45917 4019 45951
rect 4445 45917 4479 45951
rect 6377 45917 6411 45951
rect 8401 45917 8435 45951
rect 11069 45917 11103 45951
rect 13093 45917 13127 45951
rect 14105 45917 14139 45951
rect 17325 45917 17359 45951
rect 17969 45917 18003 45951
rect 18613 45917 18647 45951
rect 20361 45917 20395 45951
rect 21097 45917 21131 45951
rect 21557 45917 21591 45951
rect 22385 45917 22419 45951
rect 24869 45917 24903 45951
rect 26709 45917 26743 45951
rect 27813 45917 27847 45951
rect 28457 45917 28491 45951
rect 28549 45917 28583 45951
rect 29745 45917 29779 45951
rect 30389 45917 30423 45951
rect 31033 45917 31067 45951
rect 31861 45917 31895 45951
rect 33793 45917 33827 45951
rect 35357 45917 35391 45951
rect 36001 45917 36035 45951
rect 37933 45917 37967 45951
rect 38485 45917 38519 45951
rect 39129 45917 39163 45951
rect 39865 45917 39899 45951
rect 40785 45917 40819 45951
rect 41705 45917 41739 45951
rect 42441 45917 42475 45951
rect 42901 45917 42935 45951
rect 43637 45917 43671 45951
rect 44097 45917 44131 45951
rect 45661 45917 45695 45951
rect 46397 45917 46431 45951
rect 47133 45917 47167 45951
rect 47869 45917 47903 45951
rect 4712 45849 4746 45883
rect 6622 45849 6656 45883
rect 9220 45849 9254 45883
rect 11336 45849 11370 45883
rect 14372 45849 14406 45883
rect 17058 45849 17092 45883
rect 19717 45849 19751 45883
rect 22652 45849 22686 45883
rect 25136 45849 25170 45883
rect 32106 45849 32140 45883
rect 36268 45849 36302 45883
rect 5825 45781 5859 45815
rect 7757 45781 7791 45815
rect 10333 45781 10367 45815
rect 15485 45781 15519 45815
rect 15945 45781 15979 45815
rect 23765 45781 23799 45815
rect 26249 45781 26283 45815
rect 28457 45781 28491 45815
rect 33241 45781 33275 45815
rect 34805 45781 34839 45815
rect 37381 45781 37415 45815
rect 48053 45781 48087 45815
rect 5273 45577 5307 45611
rect 6469 45577 6503 45611
rect 9321 45577 9355 45611
rect 11529 45577 11563 45611
rect 14289 45577 14323 45611
rect 22753 45577 22787 45611
rect 25053 45577 25087 45611
rect 29561 45577 29595 45611
rect 41061 45577 41095 45611
rect 42441 45577 42475 45611
rect 43453 45577 43487 45611
rect 43913 45577 43947 45611
rect 44649 45577 44683 45611
rect 48053 45577 48087 45611
rect 15577 45509 15611 45543
rect 17509 45509 17543 45543
rect 30205 45509 30239 45543
rect 31585 45509 31619 45543
rect 32229 45509 32263 45543
rect 32781 45509 32815 45543
rect 36645 45509 36679 45543
rect 37534 45509 37568 45543
rect 39221 45509 39255 45543
rect 1777 45441 1811 45475
rect 3534 45441 3568 45475
rect 4537 45441 4571 45475
rect 4721 45441 4755 45475
rect 5089 45441 5123 45475
rect 6653 45441 6687 45475
rect 7021 45441 7055 45475
rect 7205 45441 7239 45475
rect 7849 45441 7883 45475
rect 8585 45441 8619 45475
rect 8769 45441 8803 45475
rect 8861 45441 8895 45475
rect 9137 45441 9171 45475
rect 9965 45441 9999 45475
rect 10425 45441 10459 45475
rect 11713 45441 11747 45475
rect 12081 45441 12115 45475
rect 12265 45441 12299 45475
rect 12909 45441 12943 45475
rect 13553 45441 13587 45475
rect 13737 45441 13771 45475
rect 14105 45441 14139 45475
rect 14841 45441 14875 45475
rect 15025 45441 15059 45475
rect 15393 45441 15427 45475
rect 17325 45441 17359 45475
rect 18604 45441 18638 45475
rect 22937 45441 22971 45475
rect 23305 45441 23339 45475
rect 23489 45441 23523 45475
rect 24317 45441 24351 45475
rect 24501 45441 24535 45475
rect 24869 45441 24903 45475
rect 25513 45441 25547 45475
rect 28437 45441 28471 45475
rect 3801 45373 3835 45407
rect 4813 45373 4847 45407
rect 4905 45373 4939 45407
rect 5733 45373 5767 45407
rect 6837 45373 6871 45407
rect 6929 45373 6963 45407
rect 8953 45373 8987 45407
rect 11897 45373 11931 45407
rect 11989 45373 12023 45407
rect 13829 45373 13863 45407
rect 13921 45373 13955 45407
rect 15117 45373 15151 45407
rect 15209 45373 15243 45407
rect 18337 45373 18371 45407
rect 22293 45373 22327 45407
rect 23121 45373 23155 45407
rect 23213 45373 23247 45407
rect 24593 45373 24627 45407
rect 24685 45373 24719 45407
rect 27169 45373 27203 45407
rect 28181 45373 28215 45407
rect 30849 45441 30883 45475
rect 31033 45441 31067 45475
rect 31401 45441 31435 45475
rect 33241 45441 33275 45475
rect 33508 45441 33542 45475
rect 35909 45441 35943 45475
rect 36093 45441 36127 45475
rect 36277 45441 36311 45475
rect 36461 45441 36495 45475
rect 42625 45441 42659 45475
rect 43269 45441 43303 45475
rect 44465 45441 44499 45475
rect 45109 45441 45143 45475
rect 46029 45441 46063 45475
rect 46765 45441 46799 45475
rect 47869 45441 47903 45475
rect 30389 45373 30423 45407
rect 31125 45373 31159 45407
rect 31217 45373 31251 45407
rect 36185 45373 36219 45407
rect 37289 45373 37323 45407
rect 1961 45305 1995 45339
rect 8033 45305 8067 45339
rect 9781 45305 9815 45339
rect 10609 45305 10643 45339
rect 13093 45305 13127 45339
rect 16681 45305 16715 45339
rect 20177 45305 20211 45339
rect 20821 45305 20855 45339
rect 25697 45305 25731 45339
rect 30205 45305 30239 45339
rect 46213 45305 46247 45339
rect 2421 45237 2455 45271
rect 16129 45237 16163 45271
rect 19717 45237 19751 45271
rect 26249 45237 26283 45271
rect 34621 45237 34655 45271
rect 35357 45237 35391 45271
rect 38669 45237 38703 45271
rect 39681 45237 39715 45271
rect 45293 45237 45327 45271
rect 46949 45237 46983 45271
rect 2513 45033 2547 45067
rect 5549 45033 5583 45067
rect 6929 45033 6963 45067
rect 7849 45033 7883 45067
rect 14381 45033 14415 45067
rect 15669 45033 15703 45067
rect 19809 45033 19843 45067
rect 21741 45033 21775 45067
rect 22937 45033 22971 45067
rect 25145 45033 25179 45067
rect 25697 45033 25731 45067
rect 26985 45033 27019 45067
rect 28273 45033 28307 45067
rect 33517 45033 33551 45067
rect 34069 45033 34103 45067
rect 36461 45033 36495 45067
rect 39037 45033 39071 45067
rect 43913 45033 43947 45067
rect 45109 45033 45143 45067
rect 46029 45033 46063 45067
rect 47869 45033 47903 45067
rect 4997 44965 5031 44999
rect 10149 44965 10183 44999
rect 18705 44965 18739 44999
rect 19349 44965 19383 44999
rect 30297 44965 30331 44999
rect 31769 44965 31803 44999
rect 2973 44897 3007 44931
rect 18245 44897 18279 44931
rect 27721 44897 27755 44931
rect 28641 44897 28675 44931
rect 2697 44829 2731 44863
rect 2881 44829 2915 44863
rect 3065 44829 3099 44863
rect 3249 44829 3283 44863
rect 11805 44829 11839 44863
rect 12633 44829 12667 44863
rect 14197 44829 14231 44863
rect 15485 44829 15519 44863
rect 17969 44829 18003 44863
rect 18153 44831 18187 44865
rect 30389 44897 30423 44931
rect 33149 44897 33183 44931
rect 36001 44897 36035 44931
rect 18337 44829 18371 44863
rect 18521 44829 18555 44863
rect 20361 44829 20395 44863
rect 22293 44829 22327 44863
rect 22753 44829 22787 44863
rect 24593 44829 24627 44863
rect 28457 44829 28491 44863
rect 28733 44829 28767 44863
rect 28825 44829 28859 44863
rect 29009 44829 29043 44863
rect 30297 44829 30331 44863
rect 32781 44829 32815 44863
rect 32965 44829 32999 44863
rect 33057 44829 33091 44863
rect 33333 44829 33367 44863
rect 35725 44829 35759 44863
rect 35909 44829 35943 44863
rect 36093 44829 36127 44863
rect 36277 44829 36311 44863
rect 45845 44829 45879 44863
rect 46949 44829 46983 44863
rect 47685 44829 47719 44863
rect 4445 44761 4479 44795
rect 20628 44761 20662 44795
rect 29653 44761 29687 44795
rect 30634 44761 30668 44795
rect 2053 44693 2087 44727
rect 3893 44693 3927 44727
rect 6377 44693 6411 44727
rect 8309 44693 8343 44727
rect 9505 44693 9539 44727
rect 10793 44693 10827 44727
rect 11253 44693 11287 44727
rect 11989 44693 12023 44727
rect 13461 44693 13495 44727
rect 14933 44693 14967 44727
rect 16221 44693 16255 44727
rect 17417 44693 17451 44727
rect 23857 44693 23891 44727
rect 24409 44693 24443 44727
rect 32229 44693 32263 44727
rect 35173 44693 35207 44727
rect 44373 44693 44407 44727
rect 47133 44693 47167 44727
rect 9965 44489 9999 44523
rect 10149 44489 10183 44523
rect 14473 44489 14507 44523
rect 15025 44489 15059 44523
rect 15853 44489 15887 44523
rect 17969 44489 18003 44523
rect 19625 44489 19659 44523
rect 20913 44489 20947 44523
rect 46397 44489 46431 44523
rect 9045 44421 9079 44455
rect 9229 44421 9263 44455
rect 7941 44353 7975 44387
rect 10241 44353 10275 44387
rect 11713 44353 11747 44387
rect 11989 44353 12023 44387
rect 12081 44353 12115 44387
rect 12265 44353 12299 44387
rect 13829 44353 13863 44387
rect 14381 44353 14415 44387
rect 2145 44285 2179 44319
rect 2605 44285 2639 44319
rect 4353 44285 4387 44319
rect 9965 44285 9999 44319
rect 11897 44285 11931 44319
rect 3709 44217 3743 44251
rect 8125 44217 8159 44251
rect 27721 44421 27755 44455
rect 30481 44421 30515 44455
rect 34253 44421 34287 44455
rect 44741 44421 44775 44455
rect 19533 44353 19567 44387
rect 20177 44353 20211 44387
rect 20361 44353 20395 44387
rect 20453 44353 20487 44387
rect 20729 44353 20763 44387
rect 22293 44353 22327 44387
rect 23029 44353 23063 44387
rect 23581 44353 23615 44387
rect 23765 44353 23799 44387
rect 25053 44353 25087 44387
rect 25309 44353 25343 44387
rect 27537 44353 27571 44387
rect 30682 44353 30716 44387
rect 30941 44353 30975 44387
rect 31045 44355 31079 44389
rect 31217 44353 31251 44387
rect 45293 44353 45327 44387
rect 45845 44353 45879 44387
rect 47869 44353 47903 44387
rect 20545 44285 20579 44319
rect 28365 44285 28399 44319
rect 28641 44285 28675 44319
rect 30849 44285 30883 44319
rect 3157 44149 3191 44183
rect 4905 44149 4939 44183
rect 7389 44149 7423 44183
rect 10885 44149 10919 44183
rect 11529 44149 11563 44183
rect 12817 44149 12851 44183
rect 16773 44149 16807 44183
rect 17969 44149 18003 44183
rect 18153 44149 18187 44183
rect 18981 44149 19015 44183
rect 22385 44149 22419 44183
rect 24317 44149 24351 44183
rect 26433 44149 26467 44183
rect 29653 44149 29687 44183
rect 34897 44149 34931 44183
rect 46949 44149 46983 44183
rect 48053 44149 48087 44183
rect 1869 43945 1903 43979
rect 5917 43945 5951 43979
rect 12725 43945 12759 43979
rect 47501 43945 47535 43979
rect 48053 43945 48087 43979
rect 3893 43877 3927 43911
rect 7573 43877 7607 43911
rect 3249 43809 3283 43843
rect 8309 43809 8343 43843
rect 11897 43809 11931 43843
rect 11630 43741 11664 43775
rect 2982 43673 3016 43707
rect 4905 43673 4939 43707
rect 7757 43673 7791 43707
rect 9413 43673 9447 43707
rect 37749 43877 37783 43911
rect 45661 43877 45695 43911
rect 46213 43877 46247 43911
rect 46765 43877 46799 43911
rect 13093 43809 13127 43843
rect 13185 43809 13219 43843
rect 15577 43809 15611 43843
rect 17049 43809 17083 43843
rect 20085 43809 20119 43843
rect 23489 43809 23523 43843
rect 24777 43809 24811 43843
rect 25145 43809 25179 43843
rect 27353 43809 27387 43843
rect 32956 43809 32990 43843
rect 35449 43809 35483 43843
rect 36369 43809 36403 43843
rect 12817 43741 12851 43775
rect 13001 43741 13035 43775
rect 13369 43741 13403 43775
rect 16865 43741 16899 43775
rect 17141 43741 17175 43775
rect 17233 43741 17267 43775
rect 17417 43741 17451 43775
rect 19809 43741 19843 43775
rect 20637 43741 20671 43775
rect 23305 43741 23339 43775
rect 23581 43741 23615 43775
rect 23673 43741 23707 43775
rect 23857 43741 23891 43775
rect 24409 43741 24443 43775
rect 24593 43741 24627 43775
rect 24685 43741 24719 43775
rect 24961 43741 24995 43775
rect 28457 43741 28491 43775
rect 28641 43741 28675 43775
rect 28730 43741 28764 43775
rect 28825 43743 28859 43777
rect 29009 43741 29043 43775
rect 32689 43741 32723 43775
rect 32873 43741 32907 43775
rect 33057 43741 33091 43775
rect 33241 43741 33275 43775
rect 35173 43741 35207 43775
rect 35357 43741 35391 43775
rect 35541 43741 35575 43775
rect 35725 43741 35759 43775
rect 47317 43741 47351 43775
rect 15761 43673 15795 43707
rect 21373 43673 21407 43707
rect 22661 43673 22695 43707
rect 36614 43673 36648 43707
rect 4445 43605 4479 43639
rect 9505 43605 9539 43639
rect 10517 43605 10551 43639
rect 12725 43605 12759 43639
rect 13553 43605 13587 43639
rect 14197 43605 14231 43639
rect 16681 43605 16715 43639
rect 21281 43605 21315 43639
rect 23121 43605 23155 43639
rect 28273 43605 28307 43639
rect 29561 43605 29595 43639
rect 30389 43605 30423 43639
rect 31953 43605 31987 43639
rect 32505 43605 32539 43639
rect 34989 43605 35023 43639
rect 3065 43401 3099 43435
rect 3709 43401 3743 43435
rect 5825 43401 5859 43435
rect 8125 43401 8159 43435
rect 9965 43401 9999 43435
rect 10609 43401 10643 43435
rect 14473 43401 14507 43435
rect 15025 43401 15059 43435
rect 16037 43401 16071 43435
rect 18061 43401 18095 43435
rect 18521 43401 18555 43435
rect 22017 43401 22051 43435
rect 24317 43401 24351 43435
rect 26341 43401 26375 43435
rect 29561 43401 29595 43435
rect 30205 43401 30239 43435
rect 33609 43401 33643 43435
rect 35081 43401 35115 43435
rect 36369 43401 36403 43435
rect 12173 43333 12207 43367
rect 16948 43333 16982 43367
rect 28426 43333 28460 43367
rect 30113 43333 30147 43367
rect 33517 43333 33551 43367
rect 34161 43333 34195 43367
rect 2329 43265 2363 43299
rect 2513 43265 2547 43299
rect 2697 43265 2731 43299
rect 2881 43265 2915 43299
rect 3525 43265 3559 43299
rect 4445 43265 4479 43299
rect 4712 43265 4746 43299
rect 6745 43265 6779 43299
rect 7012 43265 7046 43299
rect 8953 43265 8987 43299
rect 9873 43265 9907 43299
rect 10701 43265 10735 43299
rect 11989 43265 12023 43299
rect 13093 43265 13127 43299
rect 13360 43265 13394 43299
rect 16681 43265 16715 43299
rect 19634 43265 19668 43299
rect 20361 43265 20395 43299
rect 20545 43265 20579 43299
rect 20729 43265 20763 43299
rect 20913 43265 20947 43299
rect 21833 43265 21867 43299
rect 22937 43265 22971 43299
rect 23204 43265 23238 43299
rect 24961 43265 24995 43299
rect 25228 43265 25262 43299
rect 31585 43265 31619 43299
rect 32413 43265 32447 43299
rect 35633 43265 35667 43299
rect 35817 43265 35851 43299
rect 35909 43265 35943 43299
rect 36185 43265 36219 43299
rect 47869 43265 47903 43299
rect 2605 43197 2639 43231
rect 19901 43197 19935 43231
rect 20637 43197 20671 43231
rect 28181 43197 28215 43231
rect 32137 43197 32171 43231
rect 36001 43197 36035 43231
rect 48053 43129 48087 43163
rect 1777 43061 1811 43095
rect 9229 43061 9263 43095
rect 21097 43061 21131 43095
rect 31493 43061 31527 43095
rect 46949 43061 46983 43095
rect 5549 42857 5583 42891
rect 7113 42857 7147 42891
rect 8309 42857 8343 42891
rect 10517 42857 10551 42891
rect 11989 42857 12023 42891
rect 21005 42857 21039 42891
rect 23305 42857 23339 42891
rect 25145 42857 25179 42891
rect 29929 42857 29963 42891
rect 34069 42857 34103 42891
rect 36277 42789 36311 42823
rect 2697 42721 2731 42755
rect 4353 42721 4387 42755
rect 5181 42721 5215 42755
rect 6745 42721 6779 42755
rect 17877 42721 17911 42755
rect 18337 42721 18371 42755
rect 19625 42721 19659 42755
rect 21925 42721 21959 42755
rect 24777 42721 24811 42755
rect 2513 42653 2547 42687
rect 2780 42653 2814 42687
rect 2881 42647 2915 42681
rect 3065 42653 3099 42687
rect 4813 42653 4847 42687
rect 4997 42653 5031 42687
rect 5089 42653 5123 42687
rect 5365 42653 5399 42687
rect 6377 42653 6411 42687
rect 6561 42653 6595 42687
rect 6653 42653 6687 42687
rect 6929 42653 6963 42687
rect 8217 42653 8251 42687
rect 9413 42653 9447 42687
rect 10517 42653 10551 42687
rect 17601 42653 17635 42687
rect 17785 42653 17819 42687
rect 17969 42653 18003 42687
rect 18153 42653 18187 42687
rect 19892 42653 19926 42687
rect 22201 42653 22235 42687
rect 24409 42653 24443 42687
rect 24593 42653 24627 42687
rect 24685 42653 24719 42687
rect 24961 42653 24995 42687
rect 30573 42653 30607 42687
rect 30757 42653 30791 42687
rect 32689 42653 32723 42687
rect 34897 42653 34931 42687
rect 47869 42653 47903 42687
rect 1869 42585 1903 42619
rect 23397 42585 23431 42619
rect 31217 42585 31251 42619
rect 32934 42585 32968 42619
rect 35142 42585 35176 42619
rect 2329 42517 2363 42551
rect 7757 42517 7791 42551
rect 9689 42517 9723 42551
rect 17141 42517 17175 42551
rect 30665 42517 30699 42551
rect 31953 42517 31987 42551
rect 47317 42517 47351 42551
rect 48053 42517 48087 42551
rect 4261 42313 4295 42347
rect 4813 42313 4847 42347
rect 8309 42313 8343 42347
rect 10241 42313 10275 42347
rect 46949 42313 46983 42347
rect 3442 42245 3476 42279
rect 9137 42245 9171 42279
rect 20269 42245 20303 42279
rect 24133 42245 24167 42279
rect 1685 42177 1719 42211
rect 3709 42177 3743 42211
rect 30205 42177 30239 42211
rect 30472 42177 30506 42211
rect 47869 42177 47903 42211
rect 2329 42041 2363 42075
rect 24133 42041 24167 42075
rect 1501 41973 1535 42007
rect 6469 41973 6503 42007
rect 24225 41973 24259 42007
rect 31585 41973 31619 42007
rect 48053 41973 48087 42007
rect 1961 41769 1995 41803
rect 3893 41769 3927 41803
rect 3249 41701 3283 41735
rect 30573 41701 30607 41735
rect 31125 41701 31159 41735
rect 31585 41633 31619 41667
rect 2145 41565 2179 41599
rect 2697 41565 2731 41599
rect 31309 41565 31343 41599
rect 31401 41565 31435 41599
rect 31677 41565 31711 41599
rect 47409 41565 47443 41599
rect 48053 41565 48087 41599
rect 47869 41497 47903 41531
rect 30757 41225 30791 41259
rect 48053 41089 48087 41123
rect 47869 40953 47903 40987
rect 47593 40681 47627 40715
rect 48053 40341 48087 40375
rect 13829 40069 13863 40103
rect 48053 40069 48087 40103
rect 13645 40001 13679 40035
rect 47961 39797 47995 39831
rect 47409 39321 47443 39355
rect 48053 39321 48087 39355
rect 47961 39253 47995 39287
rect 47041 38913 47075 38947
rect 48053 38913 48087 38947
rect 47869 38777 47903 38811
rect 27997 38437 28031 38471
rect 27813 38233 27847 38267
rect 47409 38233 47443 38267
rect 48053 38233 48087 38267
rect 47961 38165 47995 38199
rect 48053 37825 48087 37859
rect 47869 37689 47903 37723
rect 47593 37417 47627 37451
rect 48053 37077 48087 37111
rect 48053 36737 48087 36771
rect 47869 36601 47903 36635
rect 9965 36329 9999 36363
rect 2145 36261 2179 36295
rect 1685 36125 1719 36159
rect 2329 36125 2363 36159
rect 2881 36125 2915 36159
rect 10057 36057 10091 36091
rect 47409 36057 47443 36091
rect 48053 36057 48087 36091
rect 1501 35989 1535 36023
rect 47961 35989 47995 36023
rect 47041 35649 47075 35683
rect 48053 35649 48087 35683
rect 47869 35513 47903 35547
rect 47409 34969 47443 35003
rect 48053 34969 48087 35003
rect 47961 34901 47995 34935
rect 48053 34561 48087 34595
rect 47869 34493 47903 34527
rect 47593 34153 47627 34187
rect 48053 33813 48087 33847
rect 48053 33473 48087 33507
rect 47869 33337 47903 33371
rect 47409 32793 47443 32827
rect 48053 32793 48087 32827
rect 47961 32725 47995 32759
rect 23397 32453 23431 32487
rect 23213 32385 23247 32419
rect 47041 32385 47075 32419
rect 48053 32385 48087 32419
rect 47869 32249 47903 32283
rect 15945 31909 15979 31943
rect 47869 31841 47903 31875
rect 48973 31841 49007 31875
rect 16129 31773 16163 31807
rect 47409 31773 47443 31807
rect 48053 31773 48087 31807
rect 48053 31297 48087 31331
rect 47869 31161 47903 31195
rect 47593 30889 47627 30923
rect 2145 30821 2179 30855
rect 1685 30685 1719 30719
rect 2329 30685 2363 30719
rect 1501 30549 1535 30583
rect 2881 30549 2915 30583
rect 48053 30549 48087 30583
rect 48053 30209 48087 30243
rect 47961 30005 47995 30039
rect 47409 29529 47443 29563
rect 48053 29529 48087 29563
rect 47961 29461 47995 29495
rect 47041 29121 47075 29155
rect 48053 29121 48087 29155
rect 47869 28985 47903 29019
rect 47409 28441 47443 28475
rect 48053 28441 48087 28475
rect 47961 28373 47995 28407
rect 48053 28033 48087 28067
rect 47961 27829 47995 27863
rect 48145 27557 48179 27591
rect 47593 27285 47627 27319
rect 48053 26945 48087 26979
rect 47869 26809 47903 26843
rect 47961 26537 47995 26571
rect 47409 26265 47443 26299
rect 48053 26265 48087 26299
rect 47041 25857 47075 25891
rect 48053 25857 48087 25891
rect 47869 25721 47903 25755
rect 19993 25313 20027 25347
rect 1685 25245 1719 25279
rect 21649 25177 21683 25211
rect 47409 25177 47443 25211
rect 48053 25177 48087 25211
rect 1501 25109 1535 25143
rect 22201 25109 22235 25143
rect 47961 25109 47995 25143
rect 1961 24905 1995 24939
rect 2145 24769 2179 24803
rect 47041 24769 47075 24803
rect 48053 24769 48087 24803
rect 47869 24633 47903 24667
rect 2697 24565 2731 24599
rect 47409 24089 47443 24123
rect 48053 24089 48087 24123
rect 47961 24021 47995 24055
rect 47409 23001 47443 23035
rect 48053 23001 48087 23035
rect 47961 22933 47995 22967
rect 47041 22593 47075 22627
rect 48053 22593 48087 22627
rect 47869 22457 47903 22491
rect 47409 21981 47443 22015
rect 46857 21913 46891 21947
rect 48053 21913 48087 21947
rect 47961 21845 47995 21879
rect 48053 21505 48087 21539
rect 47041 21369 47075 21403
rect 47961 21301 47995 21335
rect 47317 21029 47351 21063
rect 46305 20893 46339 20927
rect 47501 20893 47535 20927
rect 48145 20893 48179 20927
rect 46857 20757 46891 20791
rect 47961 20757 47995 20791
rect 46397 20553 46431 20587
rect 47041 20553 47075 20587
rect 48145 20417 48179 20451
rect 47961 20213 47995 20247
rect 46949 19873 46983 19907
rect 47869 19873 47903 19907
rect 1685 19805 1719 19839
rect 45753 19805 45787 19839
rect 45937 19805 45971 19839
rect 46305 19805 46339 19839
rect 46397 19805 46431 19839
rect 47409 19805 47443 19839
rect 47593 19805 47627 19839
rect 47961 19805 47995 19839
rect 45293 19737 45327 19771
rect 1501 19669 1535 19703
rect 1961 19465 1995 19499
rect 2697 19465 2731 19499
rect 2145 19329 2179 19363
rect 45845 19329 45879 19363
rect 46305 19329 46339 19363
rect 46489 19329 46523 19363
rect 46857 19329 46891 19363
rect 48145 19329 48179 19363
rect 46765 19261 46799 19295
rect 45385 19193 45419 19227
rect 44833 19125 44867 19159
rect 47961 19125 47995 19159
rect 45845 18853 45879 18887
rect 47409 18785 47443 18819
rect 47869 18785 47903 18819
rect 45293 18717 45327 18751
rect 46305 18717 46339 18751
rect 47593 18717 47627 18751
rect 47961 18717 47995 18751
rect 46489 18581 46523 18615
rect 47041 18581 47075 18615
rect 44833 18309 44867 18343
rect 45385 18241 45419 18275
rect 46489 18241 46523 18275
rect 46857 18241 46891 18275
rect 47041 18241 47075 18275
rect 48145 18241 48179 18275
rect 46397 18173 46431 18207
rect 46121 18037 46155 18071
rect 47961 18037 47995 18071
rect 46489 17765 46523 17799
rect 47409 17697 47443 17731
rect 47869 17697 47903 17731
rect 47593 17629 47627 17663
rect 47961 17629 47995 17663
rect 45937 17493 45971 17527
rect 47041 17493 47075 17527
rect 46489 17153 46523 17187
rect 46857 17153 46891 17187
rect 46949 17153 46983 17187
rect 48145 17153 48179 17187
rect 45845 17085 45879 17119
rect 46305 17085 46339 17119
rect 45385 17017 45419 17051
rect 47961 16949 47995 16983
rect 45845 16745 45879 16779
rect 46489 16745 46523 16779
rect 45293 16609 45327 16643
rect 46305 16541 46339 16575
rect 47409 16541 47443 16575
rect 47593 16541 47627 16575
rect 47961 16541 47995 16575
rect 48053 16541 48087 16575
rect 47041 16405 47075 16439
rect 47777 16201 47811 16235
rect 44925 16065 44959 16099
rect 45937 16065 45971 16099
rect 46581 16065 46615 16099
rect 47593 16065 47627 16099
rect 46121 15929 46155 15963
rect 45477 15861 45511 15895
rect 46765 15861 46799 15895
rect 45293 15657 45327 15691
rect 46949 15521 46983 15555
rect 47409 15521 47443 15555
rect 46305 15453 46339 15487
rect 47593 15453 47627 15487
rect 47961 15453 47995 15487
rect 48053 15453 48087 15487
rect 45845 15385 45879 15419
rect 46489 15317 46523 15351
rect 44741 15045 44775 15079
rect 44189 14977 44223 15011
rect 45201 14977 45235 15011
rect 46489 14977 46523 15011
rect 46857 14977 46891 15011
rect 47041 14977 47075 15011
rect 48145 14977 48179 15011
rect 45845 14909 45879 14943
rect 46397 14909 46431 14943
rect 45385 14773 45419 14807
rect 47961 14773 47995 14807
rect 46397 14569 46431 14603
rect 45661 14501 45695 14535
rect 47409 14433 47443 14467
rect 45477 14365 45511 14399
rect 46213 14365 46247 14399
rect 47593 14365 47627 14399
rect 47961 14365 47995 14399
rect 48053 14365 48087 14399
rect 46949 14297 46983 14331
rect 2145 14025 2179 14059
rect 45385 14025 45419 14059
rect 44833 13957 44867 13991
rect 1685 13889 1719 13923
rect 2329 13889 2363 13923
rect 46489 13889 46523 13923
rect 46857 13889 46891 13923
rect 47041 13889 47075 13923
rect 48145 13889 48179 13923
rect 2789 13821 2823 13855
rect 45845 13821 45879 13855
rect 46581 13821 46615 13855
rect 1501 13753 1535 13787
rect 47961 13685 47995 13719
rect 45293 13481 45327 13515
rect 45845 13345 45879 13379
rect 44465 13277 44499 13311
rect 46305 13277 46339 13311
rect 47409 13277 47443 13311
rect 47593 13277 47627 13311
rect 47961 13277 47995 13311
rect 48053 13277 48087 13311
rect 46489 13141 46523 13175
rect 47041 13141 47075 13175
rect 45385 12801 45419 12835
rect 46489 12801 46523 12835
rect 46857 12801 46891 12835
rect 47041 12801 47075 12835
rect 48145 12801 48179 12835
rect 45845 12733 45879 12767
rect 46581 12733 46615 12767
rect 44833 12665 44867 12699
rect 47961 12597 47995 12631
rect 46489 12393 46523 12427
rect 45845 12325 45879 12359
rect 47869 12257 47903 12291
rect 45293 12189 45327 12223
rect 46305 12189 46339 12223
rect 47409 12189 47443 12223
rect 47593 12189 47627 12223
rect 47961 12189 47995 12223
rect 48973 12189 49007 12223
rect 49065 30005 49099 30039
rect 47041 12053 47075 12087
rect 45385 11781 45419 11815
rect 46489 11713 46523 11747
rect 46857 11713 46891 11747
rect 46949 11713 46983 11747
rect 48145 11713 48179 11747
rect 45845 11645 45879 11679
rect 46581 11645 46615 11679
rect 2053 11509 2087 11543
rect 44833 11509 44867 11543
rect 47961 11509 47995 11543
rect 46397 11305 46431 11339
rect 45753 11169 45787 11203
rect 47409 11169 47443 11203
rect 46213 11101 46247 11135
rect 47593 11101 47627 11135
rect 47961 11101 47995 11135
rect 48053 11101 48087 11135
rect 1777 11033 1811 11067
rect 2605 11033 2639 11067
rect 3157 11033 3191 11067
rect 3893 11033 3927 11067
rect 4445 11033 4479 11067
rect 4997 11033 5031 11067
rect 46949 11033 46983 11067
rect 46765 10761 46799 10795
rect 46581 10625 46615 10659
rect 48145 10625 48179 10659
rect 45569 10557 45603 10591
rect 4261 10489 4295 10523
rect 1501 10421 1535 10455
rect 2053 10421 2087 10455
rect 2513 10421 2547 10455
rect 3249 10421 3283 10455
rect 3801 10421 3835 10455
rect 4813 10421 4847 10455
rect 5365 10421 5399 10455
rect 46121 10421 46155 10455
rect 47961 10421 47995 10455
rect 45753 10217 45787 10251
rect 3801 10013 3835 10047
rect 45293 10013 45327 10047
rect 46305 10013 46339 10047
rect 47409 10013 47443 10047
rect 47593 10013 47627 10047
rect 47961 10013 47995 10047
rect 48053 10013 48087 10047
rect 1961 9945 1995 9979
rect 3065 9945 3099 9979
rect 1409 9877 1443 9911
rect 2513 9877 2547 9911
rect 4353 9877 4387 9911
rect 5181 9877 5215 9911
rect 5825 9877 5859 9911
rect 6469 9877 6503 9911
rect 46489 9877 46523 9911
rect 47041 9877 47075 9911
rect 8125 9605 8159 9639
rect 45385 9605 45419 9639
rect 46489 9537 46523 9571
rect 46857 9537 46891 9571
rect 47041 9537 47075 9571
rect 48145 9537 48179 9571
rect 2513 9469 2547 9503
rect 8677 9469 8711 9503
rect 45845 9469 45879 9503
rect 46581 9469 46615 9503
rect 49065 9469 49099 9503
rect 7573 9401 7607 9435
rect 1501 9333 1535 9367
rect 1961 9333 1995 9367
rect 3065 9333 3099 9367
rect 3709 9333 3743 9367
rect 4445 9333 4479 9367
rect 4905 9333 4939 9367
rect 5549 9333 5583 9367
rect 6377 9333 6411 9367
rect 6929 9333 6963 9367
rect 44833 9333 44867 9367
rect 47961 9333 47995 9367
rect 1593 9129 1627 9163
rect 46397 9129 46431 9163
rect 45753 9061 45787 9095
rect 47409 8993 47443 9027
rect 1409 8925 1443 8959
rect 7113 8925 7147 8959
rect 46213 8925 46247 8959
rect 47593 8925 47627 8959
rect 47961 8925 47995 8959
rect 48053 8925 48087 8959
rect 6653 8857 6687 8891
rect 8953 8857 8987 8891
rect 46949 8857 46983 8891
rect 2421 8789 2455 8823
rect 2973 8789 3007 8823
rect 3801 8789 3835 8823
rect 4353 8789 4387 8823
rect 4905 8789 4939 8823
rect 5549 8789 5583 8823
rect 6101 8789 6135 8823
rect 7665 8789 7699 8823
rect 8309 8789 8343 8823
rect 9505 8789 9539 8823
rect 10057 8789 10091 8823
rect 45201 8789 45235 8823
rect 2145 8585 2179 8619
rect 44649 8585 44683 8619
rect 47777 8585 47811 8619
rect 45845 8517 45879 8551
rect 1685 8449 1719 8483
rect 2329 8449 2363 8483
rect 3433 8449 3467 8483
rect 4077 8449 4111 8483
rect 44189 8449 44223 8483
rect 45201 8449 45235 8483
rect 46489 8449 46523 8483
rect 46857 8449 46891 8483
rect 47041 8449 47075 8483
rect 47593 8449 47627 8483
rect 7205 8381 7239 8415
rect 46397 8381 46431 8415
rect 1501 8313 1535 8347
rect 4721 8313 4755 8347
rect 5181 8313 5215 8347
rect 5825 8313 5859 8347
rect 7665 8313 7699 8347
rect 45385 8313 45419 8347
rect 2881 8245 2915 8279
rect 3617 8245 3651 8279
rect 6561 8245 6595 8279
rect 8217 8245 8251 8279
rect 8769 8245 8803 8279
rect 9321 8245 9355 8279
rect 9873 8245 9907 8279
rect 10425 8245 10459 8279
rect 45845 8041 45879 8075
rect 46489 8041 46523 8075
rect 45201 7973 45235 8007
rect 1409 7837 1443 7871
rect 2237 7837 2271 7871
rect 2881 7837 2915 7871
rect 3985 7837 4019 7871
rect 4629 7837 4663 7871
rect 5089 7837 5123 7871
rect 45661 7837 45695 7871
rect 47409 7837 47443 7871
rect 47593 7837 47627 7871
rect 47961 7837 47995 7871
rect 48053 7837 48087 7871
rect 5733 7769 5767 7803
rect 43821 7769 43855 7803
rect 1593 7701 1627 7735
rect 2421 7701 2455 7735
rect 3065 7701 3099 7735
rect 3801 7701 3835 7735
rect 4445 7701 4479 7735
rect 6653 7701 6687 7735
rect 7481 7701 7515 7735
rect 8033 7701 8067 7735
rect 9045 7701 9079 7735
rect 9781 7701 9815 7735
rect 10241 7701 10275 7735
rect 10793 7701 10827 7735
rect 11345 7701 11379 7735
rect 44281 7701 44315 7735
rect 47041 7701 47075 7735
rect 2697 7497 2731 7531
rect 9137 7497 9171 7531
rect 44557 7429 44591 7463
rect 673 7361 707 7395
rect 1409 7361 1443 7395
rect 2053 7361 2087 7395
rect 2881 7361 2915 7395
rect 3525 7361 3559 7395
rect 4537 7361 4571 7395
rect 5181 7361 5215 7395
rect 5825 7361 5859 7395
rect 6561 7361 6595 7395
rect 7205 7361 7239 7395
rect 7849 7361 7883 7395
rect 8677 7361 8711 7395
rect 9321 7361 9355 7395
rect 10241 7361 10275 7395
rect 43821 7361 43855 7395
rect 43913 7361 43947 7395
rect 44465 7361 44499 7395
rect 45109 7361 45143 7395
rect 46489 7361 46523 7395
rect 46857 7361 46891 7395
rect 949 7293 983 7327
rect 11529 7293 11563 7327
rect 45845 7293 45879 7327
rect 46397 7293 46431 7327
rect 46765 7293 46799 7327
rect 857 7225 891 7259
rect 765 6069 799 6103
rect 765 4641 799 4675
rect 673 3281 707 3315
rect 3341 7225 3375 7259
rect 10425 7225 10459 7259
rect 12725 7225 12759 7259
rect 45293 7225 45327 7259
rect 1593 7157 1627 7191
rect 2237 7157 2271 7191
rect 4353 7157 4387 7191
rect 4997 7157 5031 7191
rect 5641 7157 5675 7191
rect 6377 7157 6411 7191
rect 7021 7157 7055 7191
rect 8033 7157 8067 7191
rect 8493 7157 8527 7191
rect 10885 7157 10919 7191
rect 12081 7157 12115 7191
rect 42809 7157 42843 7191
rect 43269 7157 43303 7191
rect 47777 7157 47811 7191
rect 43821 6953 43855 6987
rect 10885 6885 10919 6919
rect 44465 6885 44499 6919
rect 47409 6817 47443 6851
rect 1409 6749 1443 6783
rect 2053 6749 2087 6783
rect 2697 6749 2731 6783
rect 4077 6749 4111 6783
rect 4813 6749 4847 6783
rect 5641 6749 5675 6783
rect 6285 6749 6319 6783
rect 6929 6749 6963 6783
rect 7573 6749 7607 6783
rect 8217 6749 8251 6783
rect 8953 6749 8987 6783
rect 9781 6749 9815 6783
rect 10425 6749 10459 6783
rect 11069 6749 11103 6783
rect 11713 6749 11747 6783
rect 12725 6749 12759 6783
rect 13277 6749 13311 6783
rect 44281 6749 44315 6783
rect 45017 6749 45051 6783
rect 45661 6749 45695 6783
rect 46489 6749 46523 6783
rect 47593 6749 47627 6783
rect 47961 6749 47995 6783
rect 48053 6749 48087 6783
rect 43269 6681 43303 6715
rect 46949 6681 46983 6715
rect 1593 6613 1627 6647
rect 2145 6613 2179 6647
rect 2881 6613 2915 6647
rect 3893 6613 3927 6647
rect 4629 6613 4663 6647
rect 5457 6613 5491 6647
rect 6101 6613 6135 6647
rect 6745 6613 6779 6647
rect 7389 6613 7423 6647
rect 8033 6613 8067 6647
rect 9045 6613 9079 6647
rect 9597 6613 9631 6647
rect 10241 6613 10275 6647
rect 11529 6613 11563 6647
rect 12173 6613 12207 6647
rect 42717 6613 42751 6647
rect 45201 6613 45235 6647
rect 45845 6613 45879 6647
rect 48973 6613 49007 6647
rect 3341 6409 3375 6443
rect 5733 6409 5767 6443
rect 9689 6409 9723 6443
rect 43269 6409 43303 6443
rect 45937 6409 45971 6443
rect 47777 6409 47811 6443
rect 14013 6341 14047 6375
rect 14565 6341 14599 6375
rect 1961 6273 1995 6307
rect 2789 6273 2823 6307
rect 3525 6273 3559 6307
rect 4261 6273 4295 6307
rect 4997 6273 5031 6307
rect 5641 6273 5675 6307
rect 6653 6273 6687 6307
rect 7389 6273 7423 6307
rect 8125 6273 8159 6307
rect 9229 6273 9263 6307
rect 9873 6273 9907 6307
rect 10517 6273 10551 6307
rect 11989 6273 12023 6307
rect 41889 6273 41923 6307
rect 43729 6273 43763 6307
rect 44373 6273 44407 6307
rect 45201 6273 45235 6307
rect 46489 6273 46523 6307
rect 46857 6273 46891 6307
rect 47041 6273 47075 6307
rect 47593 6273 47627 6307
rect 12265 6205 12299 6239
rect 46581 6205 46615 6239
rect 42717 6137 42751 6171
rect 43913 6137 43947 6171
rect 1777 6069 1811 6103
rect 2605 6069 2639 6103
rect 4077 6069 4111 6103
rect 4813 6069 4847 6103
rect 6469 6069 6503 6103
rect 7205 6069 7239 6103
rect 7941 6069 7975 6103
rect 9045 6069 9079 6103
rect 10333 6069 10367 6103
rect 12909 6069 12943 6103
rect 13461 6069 13495 6103
rect 15209 6069 15243 6103
rect 44557 6069 44591 6103
rect 45109 6069 45143 6103
rect 4077 5865 4111 5899
rect 7389 5865 7423 5899
rect 9045 5865 9079 5899
rect 14749 5865 14783 5899
rect 15853 5865 15887 5899
rect 43821 5865 43855 5899
rect 46397 5865 46431 5899
rect 2237 5797 2271 5831
rect 46121 5797 46155 5831
rect 47225 5797 47259 5831
rect 4169 5729 4203 5763
rect 12449 5729 12483 5763
rect 1685 5661 1719 5695
rect 2421 5661 2455 5695
rect 3157 5661 3191 5695
rect 5089 5661 5123 5695
rect 5825 5661 5859 5695
rect 6573 5661 6607 5695
rect 7297 5661 7331 5695
rect 7481 5661 7515 5695
rect 8401 5661 8435 5695
rect 9229 5661 9263 5695
rect 9689 5661 9723 5695
rect 9965 5661 9999 5695
rect 10885 5661 10919 5695
rect 11713 5661 11747 5695
rect 41521 5661 41555 5695
rect 43637 5661 43671 5695
rect 44281 5661 44315 5695
rect 45385 5661 45419 5695
rect 46121 5661 46155 5695
rect 46213 5661 46247 5695
rect 47409 5661 47443 5695
rect 47593 5661 47627 5695
rect 47961 5661 47995 5695
rect 48053 5661 48087 5695
rect 3985 5593 4019 5627
rect 4353 5593 4387 5627
rect 11069 5593 11103 5627
rect 11253 5593 11287 5627
rect 45605 5593 45639 5627
rect 1501 5525 1535 5559
rect 2973 5525 3007 5559
rect 4261 5525 4295 5559
rect 4905 5525 4939 5559
rect 5641 5525 5675 5559
rect 6377 5525 6411 5559
rect 7665 5525 7699 5559
rect 8217 5525 8251 5559
rect 11897 5525 11931 5559
rect 12909 5525 12943 5559
rect 13461 5525 13495 5559
rect 14105 5525 14139 5559
rect 15209 5525 15243 5559
rect 42073 5525 42107 5559
rect 42625 5525 42659 5559
rect 43177 5525 43211 5559
rect 44465 5525 44499 5559
rect 2881 5321 2915 5355
rect 15853 5321 15887 5355
rect 42809 5321 42843 5355
rect 3709 5253 3743 5287
rect 4629 5253 4663 5287
rect 10241 5253 10275 5287
rect 10977 5253 11011 5287
rect 44557 5253 44591 5287
rect 1685 5185 1719 5219
rect 2789 5185 2823 5219
rect 5733 5185 5767 5219
rect 6745 5185 6779 5219
rect 7757 5185 7791 5219
rect 8861 5185 8895 5219
rect 9873 5185 9907 5219
rect 9965 5185 9999 5219
rect 11805 5185 11839 5219
rect 13093 5185 13127 5219
rect 15301 5185 15335 5219
rect 43269 5185 43303 5219
rect 43913 5185 43947 5219
rect 45201 5185 45235 5219
rect 45569 5185 45603 5219
rect 6837 5117 6871 5151
rect 7941 5117 7975 5151
rect 8953 5117 8987 5151
rect 41889 5117 41923 5151
rect 45109 5117 45143 5151
rect 45477 5117 45511 5151
rect 3893 5049 3927 5083
rect 4905 5049 4939 5083
rect 9229 5049 9263 5083
rect 9873 5049 9907 5083
rect 11621 5049 11655 5083
rect 14657 5049 14691 5083
rect 43453 5049 43487 5083
rect 1501 4981 1535 5015
rect 2145 4981 2179 5015
rect 5549 4981 5583 5015
rect 6837 4981 6871 5015
rect 7113 4981 7147 5015
rect 8861 4981 8895 5015
rect 12265 4981 12299 5015
rect 12909 4981 12943 5015
rect 13553 4981 13587 5015
rect 14105 4981 14139 5015
rect 29101 4981 29135 5015
rect 30021 4981 30055 5015
rect 41337 4981 41371 5015
rect 44097 4981 44131 5015
rect 46213 4981 46247 5015
rect 46857 4981 46891 5015
rect 47593 4981 47627 5015
rect 1593 4777 1627 4811
rect 8953 4777 8987 4811
rect 9413 4777 9447 4811
rect 43361 4777 43395 4811
rect 2421 4709 2455 4743
rect 13093 4709 13127 4743
rect 43913 4709 43947 4743
rect 6561 4641 6595 4675
rect 9137 4641 9171 4675
rect 11069 4641 11103 4675
rect 16957 4641 16991 4675
rect 45477 4641 45511 4675
rect 45937 4641 45971 4675
rect 47409 4641 47443 4675
rect 1409 4573 1443 4607
rect 5181 4573 5215 4607
rect 6285 4573 6319 4607
rect 7205 4573 7239 4607
rect 8401 4573 8435 4607
rect 8953 4573 8987 4607
rect 9229 4573 9263 4607
rect 9873 4573 9907 4607
rect 10793 4573 10827 4607
rect 11989 4573 12023 4607
rect 12449 4573 12483 4607
rect 14105 4573 14139 4607
rect 15669 4573 15703 4607
rect 29009 4573 29043 4607
rect 30113 4573 30147 4607
rect 42533 4573 42567 4607
rect 44092 4573 44126 4607
rect 44465 4573 44499 4607
rect 45017 4573 45051 4607
rect 45661 4573 45695 4607
rect 46029 4573 46063 4607
rect 47593 4573 47627 4607
rect 47961 4573 47995 4607
rect 48053 4573 48087 4607
rect 2697 4505 2731 4539
rect 4261 4505 4295 4539
rect 5549 4505 5583 4539
rect 7481 4505 7515 4539
rect 10149 4505 10183 4539
rect 41981 4505 42015 4539
rect 44189 4505 44223 4539
rect 44281 4505 44315 4539
rect 46949 4505 46983 4539
rect 4353 4437 4387 4471
rect 8217 4437 8251 4471
rect 11805 4437 11839 4471
rect 14749 4437 14783 4471
rect 16313 4437 16347 4471
rect 28825 4437 28859 4471
rect 29561 4437 29595 4471
rect 30297 4437 30331 4471
rect 30757 4437 30791 4471
rect 31401 4437 31435 4471
rect 40417 4437 40451 4471
rect 40877 4437 40911 4471
rect 41521 4437 41555 4471
rect 42717 4437 42751 4471
rect 5641 4233 5675 4267
rect 8585 4233 8619 4267
rect 1961 4165 1995 4199
rect 6837 4165 6871 4199
rect 2329 4097 2363 4131
rect 2789 4097 2823 4131
rect 3065 4097 3099 4131
rect 3801 4097 3835 4131
rect 4528 4097 4562 4131
rect 8217 4097 8251 4131
rect 8769 4097 8803 4131
rect 9229 4097 9263 4131
rect 9505 4097 9539 4131
rect 10425 4097 10459 4131
rect 11805 4097 11839 4131
rect 12541 4097 12575 4131
rect 13277 4097 13311 4131
rect 20085 4097 20119 4131
rect 30757 4097 30791 4131
rect 31401 4097 31435 4131
rect 41245 4097 41279 4131
rect 41705 4097 41739 4131
rect 43453 4097 43487 4131
rect 45201 4097 45235 4131
rect 45569 4097 45603 4131
rect 47869 4097 47903 4131
rect 48973 4097 49007 4131
rect 2881 4029 2915 4063
rect 4261 4029 4295 4063
rect 8309 4029 8343 4063
rect 9689 4029 9723 4063
rect 10701 4029 10735 4063
rect 44557 4029 44591 4063
rect 45109 4029 45143 4063
rect 45477 4029 45511 4063
rect 949 3961 983 3995
rect 9321 3961 9355 3995
rect 13737 3961 13771 3995
rect 15669 3961 15703 3995
rect 22109 3961 22143 3995
rect 40141 3961 40175 3995
rect 46857 3961 46891 3995
rect 2789 3893 2823 3927
rect 3249 3893 3283 3927
rect 7113 3893 7147 3927
rect 11621 3893 11655 3927
rect 12357 3893 12391 3927
rect 13093 3893 13127 3927
rect 14381 3893 14415 3927
rect 15025 3893 15059 3927
rect 16681 3893 16715 3927
rect 17325 3893 17359 3927
rect 18429 3893 18463 3927
rect 27997 3893 28031 3927
rect 28641 3893 28675 3927
rect 29101 3893 29135 3927
rect 30113 3893 30147 3927
rect 30573 3893 30607 3927
rect 31217 3893 31251 3927
rect 40693 3893 40727 3927
rect 41889 3893 41923 3927
rect 42809 3893 42843 3927
rect 44097 3893 44131 3927
rect 46213 3893 46247 3927
rect 48053 3893 48087 3927
rect 1869 3689 1903 3723
rect 3065 3689 3099 3723
rect 3801 3689 3835 3723
rect 6285 3689 6319 3723
rect 6745 3689 6779 3723
rect 41889 3689 41923 3723
rect 45109 3689 45143 3723
rect 4261 3621 4295 3655
rect 7481 3621 7515 3655
rect 12725 3621 12759 3655
rect 16129 3621 16163 3655
rect 23765 3621 23799 3655
rect 30205 3621 30239 3655
rect 6561 3553 6595 3587
rect 7941 3553 7975 3587
rect 9137 3553 9171 3587
rect 11897 3553 11931 3587
rect 13369 3553 13403 3587
rect 16773 3553 16807 3587
rect 46765 3621 46799 3655
rect 47409 3553 47443 3587
rect 2145 3485 2179 3519
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 5181 3485 5215 3519
rect 6469 3485 6503 3519
rect 7389 3485 7423 3519
rect 7665 3485 7699 3519
rect 8953 3485 8987 3519
rect 9873 3485 9907 3519
rect 10149 3485 10183 3519
rect 10793 3485 10827 3519
rect 11713 3485 11747 3519
rect 12909 3485 12943 3519
rect 14381 3485 14415 3519
rect 14841 3485 14875 3519
rect 15485 3485 15519 3519
rect 17417 3485 17451 3519
rect 18061 3485 18095 3519
rect 19257 3485 19291 3519
rect 19901 3485 19935 3519
rect 20545 3485 20579 3519
rect 21189 3485 21223 3519
rect 21833 3485 21867 3519
rect 22477 3485 22511 3519
rect 23305 3485 23339 3519
rect 24409 3485 24443 3519
rect 25053 3485 25087 3519
rect 25973 3485 26007 3519
rect 26433 3485 26467 3519
rect 27353 3485 27387 3519
rect 27997 3485 28031 3519
rect 28457 3485 28491 3519
rect 29561 3485 29595 3519
rect 30849 3485 30883 3519
rect 31493 3485 31527 3519
rect 32137 3485 32171 3519
rect 33057 3485 33091 3519
rect 34713 3485 34747 3519
rect 35357 3485 35391 3519
rect 36001 3485 36035 3519
rect 36645 3485 36679 3519
rect 37289 3485 37323 3519
rect 38209 3485 38243 3519
rect 39129 3485 39163 3519
rect 40325 3485 40359 3519
rect 41245 3485 41279 3519
rect 41889 3485 41923 3519
rect 42165 3485 42199 3519
rect 42993 3485 43027 3519
rect 43821 3485 43855 3519
rect 44465 3485 44499 3519
rect 45288 3485 45322 3519
rect 45385 3485 45419 3519
rect 45661 3485 45695 3519
rect 47869 3485 47903 3519
rect 857 2941 891 2975
rect 949 3417 983 3451
rect 2789 3417 2823 3451
rect 3801 3417 3835 3451
rect 6745 3417 6779 3451
rect 11069 3417 11103 3451
rect 45477 3417 45511 3451
rect 5273 3349 5307 3383
rect 14197 3349 14231 3383
rect 48053 3349 48087 3383
rect 3065 3145 3099 3179
rect 3709 3145 3743 3179
rect 4813 3145 4847 3179
rect 5365 3145 5399 3179
rect 7297 3145 7331 3179
rect 7849 3145 7883 3179
rect 13369 3145 13403 3179
rect 14105 3145 14139 3179
rect 20361 3145 20395 3179
rect 24225 3145 24259 3179
rect 28549 3145 28583 3179
rect 28917 3145 28951 3179
rect 30849 3145 30883 3179
rect 36093 3145 36127 3179
rect 2605 3077 2639 3111
rect 4169 3077 4203 3111
rect 5825 3077 5859 3111
rect 8769 3077 8803 3111
rect 12725 3077 12759 3111
rect 18521 3077 18555 3111
rect 20269 3077 20303 3111
rect 22293 3077 22327 3111
rect 22477 3077 22511 3111
rect 29009 3077 29043 3111
rect 29837 3077 29871 3111
rect 35357 3077 35391 3111
rect 36001 3077 36035 3111
rect 1501 3009 1535 3043
rect 2789 3009 2823 3043
rect 2881 3009 2915 3043
rect 3876 3009 3910 3043
rect 4629 3009 4663 3043
rect 5549 3009 5583 3043
rect 6285 3009 6319 3043
rect 6653 3009 6687 3043
rect 6745 3009 6779 3043
rect 7113 3009 7147 3043
rect 8493 3009 8527 3043
rect 9321 3009 9355 3043
rect 9965 3009 9999 3043
rect 10241 3009 10275 3043
rect 10977 3009 11011 3043
rect 11529 3009 11563 3043
rect 12449 3009 12483 3043
rect 13921 3009 13955 3043
rect 14933 3009 14967 3043
rect 24133 3009 24167 3043
rect 41889 3009 41923 3043
rect 46305 3009 46339 3043
rect 46765 3009 46799 3043
rect 47869 3009 47903 3043
rect 2053 2941 2087 2975
rect 3985 2941 4019 2975
rect 5733 2941 5767 2975
rect 8585 2941 8619 2975
rect 10149 2941 10183 2975
rect 11805 2941 11839 2975
rect 16037 2941 16071 2975
rect 18705 2941 18739 2975
rect 25421 2941 25455 2975
rect 29101 2941 29135 2975
rect 34069 2941 34103 2975
rect 38577 2941 38611 2975
rect 8309 2873 8343 2907
rect 14749 2873 14783 2907
rect 17325 2873 17359 2907
rect 19165 2873 19199 2907
rect 20913 2873 20947 2907
rect 22937 2873 22971 2907
rect 24777 2873 24811 2907
rect 26065 2873 26099 2907
rect 2697 2805 2731 2839
rect 3985 2805 4019 2839
rect 5641 2805 5675 2839
rect 6377 2805 6411 2839
rect 7021 2805 7055 2839
rect 8769 2805 8803 2839
rect 9781 2805 9815 2839
rect 10241 2805 10275 2839
rect 10793 2805 10827 2839
rect 15393 2805 15427 2839
rect 16681 2805 16715 2839
rect 26985 2805 27019 2839
rect 27629 2805 27663 2839
rect 32137 2805 32171 2839
rect 32781 2805 32815 2839
rect 33425 2805 33459 2839
rect 34713 2805 34747 2839
rect 37289 2805 37323 2839
rect 37933 2805 37967 2839
rect 39221 2805 39255 2839
rect 39865 2805 39899 2839
rect 40509 2805 40543 2839
rect 41153 2805 41187 2839
rect 42441 2805 42475 2839
rect 43085 2805 43119 2839
rect 43729 2805 43763 2839
rect 44373 2805 44407 2839
rect 45017 2805 45051 2839
rect 46949 2805 46983 2839
rect 48053 2805 48087 2839
rect 949 2601 983 2635
rect 2789 2601 2823 2635
rect 3157 2601 3191 2635
rect 13461 2601 13495 2635
rect 14933 2601 14967 2635
rect 29009 2601 29043 2635
rect 8769 2533 8803 2567
rect 15577 2533 15611 2567
rect 17325 2533 17359 2567
rect 25053 2533 25087 2567
rect 46949 2533 46983 2567
rect 1961 2465 1995 2499
rect 3065 2465 3099 2499
rect 11713 2465 11747 2499
rect 24409 2465 24443 2499
rect 25697 2465 25731 2499
rect 27629 2465 27663 2499
rect 2237 2397 2271 2431
rect 2973 2397 3007 2431
rect 3249 2397 3283 2431
rect 5181 2397 5215 2431
rect 8769 2397 8803 2431
rect 10885 2397 10919 2431
rect 11989 2397 12023 2431
rect 12449 2397 12483 2431
rect 13369 2399 13403 2433
rect 13553 2397 13587 2431
rect 14381 2397 14415 2431
rect 15117 2397 15151 2431
rect 16681 2397 16715 2431
rect 17969 2397 18003 2431
rect 18613 2397 18647 2431
rect 19257 2397 19291 2431
rect 19901 2397 19935 2431
rect 20545 2397 20579 2431
rect 21833 2397 21867 2431
rect 22477 2397 22511 2431
rect 23213 2397 23247 2431
rect 26985 2397 27019 2431
rect 28273 2397 28307 2431
rect 30665 2397 30699 2431
rect 31309 2397 31343 2431
rect 32137 2397 32171 2431
rect 32781 2397 32815 2431
rect 33793 2397 33827 2431
rect 34713 2397 34747 2431
rect 35357 2397 35391 2431
rect 36001 2397 36035 2431
rect 37289 2397 37323 2431
rect 37933 2397 37967 2431
rect 38853 2397 38887 2431
rect 39865 2397 39899 2431
rect 40969 2397 41003 2431
rect 41429 2397 41463 2431
rect 42441 2397 42475 2431
rect 43453 2397 43487 2431
rect 44097 2397 44131 2431
rect 45017 2397 45051 2431
rect 46029 2397 46063 2431
rect 46765 2397 46799 2431
rect 47869 2397 47903 2431
rect 4261 2329 4295 2363
rect 6837 2329 6871 2363
rect 7757 2329 7791 2363
rect 9413 2329 9447 2363
rect 10333 2329 10367 2363
rect 12725 2329 12759 2363
rect 30021 2329 30055 2363
rect 4537 2261 4571 2295
rect 5457 2261 5491 2295
rect 7113 2261 7147 2295
rect 8033 2261 8067 2295
rect 9689 2261 9723 2295
rect 14197 2261 14231 2295
rect 30113 2261 30147 2295
rect 46213 2261 46247 2295
rect 48053 2261 48087 2295
rect 8861 1853 8895 1887
rect 7389 1649 7423 1683
rect 7389 1309 7423 1343
rect 8861 901 8895 935
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 1486 47240 1492 47252
rect 1447 47212 1492 47240
rect 1486 47200 1492 47212
rect 1544 47200 1550 47252
rect 1854 47200 1860 47252
rect 1912 47240 1918 47252
rect 2317 47243 2375 47249
rect 2317 47240 2329 47243
rect 1912 47212 2329 47240
rect 1912 47200 1918 47212
rect 2317 47209 2329 47212
rect 2363 47209 2375 47243
rect 2317 47203 2375 47209
rect 3050 47200 3056 47252
rect 3108 47240 3114 47252
rect 3973 47243 4031 47249
rect 3973 47240 3985 47243
rect 3108 47212 3985 47240
rect 3108 47200 3114 47212
rect 3973 47209 3985 47212
rect 4019 47209 4031 47243
rect 4614 47240 4620 47252
rect 4575 47212 4620 47240
rect 3973 47203 4031 47209
rect 4614 47200 4620 47212
rect 4672 47200 4678 47252
rect 4706 47200 4712 47252
rect 4764 47240 4770 47252
rect 5353 47243 5411 47249
rect 5353 47240 5365 47243
rect 4764 47212 5365 47240
rect 4764 47200 4770 47212
rect 5353 47209 5365 47212
rect 5399 47209 5411 47243
rect 5353 47203 5411 47209
rect 5534 47200 5540 47252
rect 5592 47240 5598 47252
rect 6549 47243 6607 47249
rect 6549 47240 6561 47243
rect 5592 47212 6561 47240
rect 5592 47200 5598 47212
rect 6549 47209 6561 47212
rect 6595 47209 6607 47243
rect 6549 47203 6607 47209
rect 6914 47200 6920 47252
rect 6972 47240 6978 47252
rect 7193 47243 7251 47249
rect 7193 47240 7205 47243
rect 6972 47212 7205 47240
rect 6972 47200 6978 47212
rect 7193 47209 7205 47212
rect 7239 47209 7251 47243
rect 8294 47240 8300 47252
rect 8255 47212 8300 47240
rect 7193 47203 7251 47209
rect 8294 47200 8300 47212
rect 8352 47200 8358 47252
rect 9306 47200 9312 47252
rect 9364 47240 9370 47252
rect 9493 47243 9551 47249
rect 9493 47240 9505 47243
rect 9364 47212 9505 47240
rect 9364 47200 9370 47212
rect 9493 47209 9505 47212
rect 9539 47209 9551 47243
rect 9493 47203 9551 47209
rect 10594 47200 10600 47252
rect 10652 47240 10658 47252
rect 10873 47243 10931 47249
rect 10873 47240 10885 47243
rect 10652 47212 10885 47240
rect 10652 47200 10658 47212
rect 10873 47209 10885 47212
rect 10919 47209 10931 47243
rect 10873 47203 10931 47209
rect 11790 47200 11796 47252
rect 11848 47240 11854 47252
rect 11977 47243 12035 47249
rect 11977 47240 11989 47243
rect 11848 47212 11989 47240
rect 11848 47200 11854 47212
rect 11977 47209 11989 47212
rect 12023 47209 12035 47243
rect 11977 47203 12035 47209
rect 13078 47200 13084 47252
rect 13136 47240 13142 47252
rect 13357 47243 13415 47249
rect 13357 47240 13369 47243
rect 13136 47212 13369 47240
rect 13136 47200 13142 47212
rect 13357 47209 13369 47212
rect 13403 47209 13415 47243
rect 13357 47203 13415 47209
rect 14274 47200 14280 47252
rect 14332 47240 14338 47252
rect 14553 47243 14611 47249
rect 14553 47240 14565 47243
rect 14332 47212 14565 47240
rect 14332 47200 14338 47212
rect 14553 47209 14565 47212
rect 14599 47209 14611 47243
rect 14553 47203 14611 47209
rect 15562 47200 15568 47252
rect 15620 47240 15626 47252
rect 15841 47243 15899 47249
rect 15841 47240 15853 47243
rect 15620 47212 15853 47240
rect 15620 47200 15626 47212
rect 15841 47209 15853 47212
rect 15887 47209 15899 47243
rect 15841 47203 15899 47209
rect 16850 47200 16856 47252
rect 16908 47240 16914 47252
rect 17037 47243 17095 47249
rect 17037 47240 17049 47243
rect 16908 47212 17049 47240
rect 16908 47200 16914 47212
rect 17037 47209 17049 47212
rect 17083 47209 17095 47243
rect 17037 47203 17095 47209
rect 18046 47200 18052 47252
rect 18104 47240 18110 47252
rect 18233 47243 18291 47249
rect 18233 47240 18245 47243
rect 18104 47212 18245 47240
rect 18104 47200 18110 47212
rect 18233 47209 18245 47212
rect 18279 47209 18291 47243
rect 18233 47203 18291 47209
rect 19334 47200 19340 47252
rect 19392 47240 19398 47252
rect 19521 47243 19579 47249
rect 19521 47240 19533 47243
rect 19392 47212 19533 47240
rect 19392 47200 19398 47212
rect 19521 47209 19533 47212
rect 19567 47209 19579 47243
rect 19521 47203 19579 47209
rect 20714 47200 20720 47252
rect 20772 47240 20778 47252
rect 20809 47243 20867 47249
rect 20809 47240 20821 47243
rect 20772 47212 20821 47240
rect 20772 47200 20778 47212
rect 20809 47209 20821 47212
rect 20855 47209 20867 47243
rect 20809 47203 20867 47209
rect 22094 47200 22100 47252
rect 22152 47240 22158 47252
rect 22152 47212 22197 47240
rect 22152 47200 22158 47212
rect 23014 47200 23020 47252
rect 23072 47240 23078 47252
rect 23293 47243 23351 47249
rect 23293 47240 23305 47243
rect 23072 47212 23305 47240
rect 23072 47200 23078 47212
rect 23293 47209 23305 47212
rect 23339 47209 23351 47243
rect 23293 47203 23351 47209
rect 24302 47200 24308 47252
rect 24360 47240 24366 47252
rect 24581 47243 24639 47249
rect 24581 47240 24593 47243
rect 24360 47212 24593 47240
rect 24360 47200 24366 47212
rect 24581 47209 24593 47212
rect 24627 47209 24639 47243
rect 24581 47203 24639 47209
rect 25590 47200 25596 47252
rect 25648 47240 25654 47252
rect 25869 47243 25927 47249
rect 25869 47240 25881 47243
rect 25648 47212 25881 47240
rect 25648 47200 25654 47212
rect 25869 47209 25881 47212
rect 25915 47209 25927 47243
rect 25869 47203 25927 47209
rect 26786 47200 26792 47252
rect 26844 47240 26850 47252
rect 27157 47243 27215 47249
rect 27157 47240 27169 47243
rect 26844 47212 27169 47240
rect 26844 47200 26850 47212
rect 27157 47209 27169 47212
rect 27203 47209 27215 47243
rect 27157 47203 27215 47209
rect 28074 47200 28080 47252
rect 28132 47240 28138 47252
rect 28353 47243 28411 47249
rect 28353 47240 28365 47243
rect 28132 47212 28365 47240
rect 28132 47200 28138 47212
rect 28353 47209 28365 47212
rect 28399 47209 28411 47243
rect 28353 47203 28411 47209
rect 29270 47200 29276 47252
rect 29328 47240 29334 47252
rect 29733 47243 29791 47249
rect 29733 47240 29745 47243
rect 29328 47212 29745 47240
rect 29328 47200 29334 47212
rect 29733 47209 29745 47212
rect 29779 47209 29791 47243
rect 29733 47203 29791 47209
rect 30558 47200 30564 47252
rect 30616 47240 30622 47252
rect 30837 47243 30895 47249
rect 30837 47240 30849 47243
rect 30616 47212 30849 47240
rect 30616 47200 30622 47212
rect 30837 47209 30849 47212
rect 30883 47209 30895 47243
rect 30837 47203 30895 47209
rect 31754 47200 31760 47252
rect 31812 47240 31818 47252
rect 32217 47243 32275 47249
rect 32217 47240 32229 47243
rect 31812 47212 32229 47240
rect 31812 47200 31818 47212
rect 32217 47209 32229 47212
rect 32263 47209 32275 47243
rect 32217 47203 32275 47209
rect 33134 47200 33140 47252
rect 33192 47240 33198 47252
rect 33229 47243 33287 47249
rect 33229 47240 33241 47243
rect 33192 47212 33241 47240
rect 33192 47200 33198 47212
rect 33229 47209 33241 47212
rect 33275 47209 33287 47243
rect 33229 47203 33287 47209
rect 33502 47200 33508 47252
rect 33560 47240 33566 47252
rect 34057 47243 34115 47249
rect 34057 47240 34069 47243
rect 33560 47212 34069 47240
rect 33560 47200 33566 47212
rect 34057 47209 34069 47212
rect 34103 47209 34115 47243
rect 34057 47203 34115 47209
rect 34514 47200 34520 47252
rect 34572 47240 34578 47252
rect 34885 47243 34943 47249
rect 34885 47240 34897 47243
rect 34572 47212 34897 47240
rect 34572 47200 34578 47212
rect 34885 47209 34897 47212
rect 34931 47209 34943 47243
rect 34885 47203 34943 47209
rect 35526 47200 35532 47252
rect 35584 47240 35590 47252
rect 35805 47243 35863 47249
rect 35805 47240 35817 47243
rect 35584 47212 35817 47240
rect 35584 47200 35590 47212
rect 35805 47209 35817 47212
rect 35851 47209 35863 47243
rect 35805 47203 35863 47209
rect 38010 47200 38016 47252
rect 38068 47240 38074 47252
rect 38197 47243 38255 47249
rect 38197 47240 38209 47243
rect 38068 47212 38209 47240
rect 38068 47200 38074 47212
rect 38197 47209 38209 47212
rect 38243 47209 38255 47243
rect 38197 47203 38255 47209
rect 38654 47200 38660 47252
rect 38712 47240 38718 47252
rect 39025 47243 39083 47249
rect 39025 47240 39037 47243
rect 38712 47212 39037 47240
rect 38712 47200 38718 47212
rect 39025 47209 39037 47212
rect 39071 47209 39083 47243
rect 39025 47203 39083 47209
rect 39298 47200 39304 47252
rect 39356 47240 39362 47252
rect 40037 47243 40095 47249
rect 40037 47240 40049 47243
rect 39356 47212 40049 47240
rect 39356 47200 39362 47212
rect 40037 47209 40049 47212
rect 40083 47209 40095 47243
rect 40037 47203 40095 47209
rect 40494 47200 40500 47252
rect 40552 47240 40558 47252
rect 40681 47243 40739 47249
rect 40681 47240 40693 47243
rect 40552 47212 40693 47240
rect 40552 47200 40558 47212
rect 40681 47209 40693 47212
rect 40727 47209 40739 47243
rect 40681 47203 40739 47209
rect 41782 47200 41788 47252
rect 41840 47240 41846 47252
rect 42613 47243 42671 47249
rect 42613 47240 42625 47243
rect 41840 47212 42625 47240
rect 41840 47200 41846 47212
rect 42613 47209 42625 47212
rect 42659 47209 42671 47243
rect 42613 47203 42671 47209
rect 43070 47200 43076 47252
rect 43128 47240 43134 47252
rect 43349 47243 43407 47249
rect 43349 47240 43361 47243
rect 43128 47212 43361 47240
rect 43128 47200 43134 47212
rect 43349 47209 43361 47212
rect 43395 47209 43407 47243
rect 43349 47203 43407 47209
rect 44266 47200 44272 47252
rect 44324 47240 44330 47252
rect 44361 47243 44419 47249
rect 44361 47240 44373 47243
rect 44324 47212 44373 47240
rect 44324 47200 44330 47212
rect 44361 47209 44373 47212
rect 44407 47209 44419 47243
rect 44361 47203 44419 47209
rect 45465 47243 45523 47249
rect 45465 47209 45477 47243
rect 45511 47240 45523 47243
rect 45646 47240 45652 47252
rect 45511 47212 45652 47240
rect 45511 47209 45523 47212
rect 45465 47203 45523 47209
rect 45646 47200 45652 47212
rect 45704 47200 45710 47252
rect 46201 47243 46259 47249
rect 46201 47209 46213 47243
rect 46247 47240 46259 47243
rect 48041 47243 48099 47249
rect 46247 47212 47716 47240
rect 46247 47209 46259 47212
rect 46201 47203 46259 47209
rect 41046 47132 41052 47184
rect 41104 47172 41110 47184
rect 41104 47144 46796 47172
rect 41104 47132 41110 47144
rect 40218 47064 40224 47116
rect 40276 47104 40282 47116
rect 46768 47104 46796 47144
rect 46842 47132 46848 47184
rect 46900 47172 46906 47184
rect 46937 47175 46995 47181
rect 46937 47172 46949 47175
rect 46900 47144 46949 47172
rect 46900 47132 46906 47144
rect 46937 47141 46949 47144
rect 46983 47141 46995 47175
rect 47688 47172 47716 47212
rect 48041 47209 48053 47243
rect 48087 47240 48099 47243
rect 48406 47240 48412 47252
rect 48087 47212 48412 47240
rect 48087 47209 48099 47212
rect 48041 47203 48099 47209
rect 48406 47200 48412 47212
rect 48464 47200 48470 47252
rect 49234 47172 49240 47184
rect 47688 47144 49240 47172
rect 46937 47135 46995 47141
rect 49234 47132 49240 47144
rect 49292 47132 49298 47184
rect 40276 47076 46060 47104
rect 46768 47076 47900 47104
rect 40276 47064 40282 47076
rect 1670 47036 1676 47048
rect 1631 47008 1676 47036
rect 1670 46996 1676 47008
rect 1728 46996 1734 47048
rect 1946 46996 1952 47048
rect 2004 47036 2010 47048
rect 2133 47039 2191 47045
rect 2133 47036 2145 47039
rect 2004 47008 2145 47036
rect 2004 46996 2010 47008
rect 2133 47005 2145 47008
rect 2179 47005 2191 47039
rect 2866 47036 2872 47048
rect 2827 47008 2872 47036
rect 2133 46999 2191 47005
rect 2866 46996 2872 47008
rect 2924 46996 2930 47048
rect 3786 47036 3792 47048
rect 3747 47008 3792 47036
rect 3786 46996 3792 47008
rect 3844 46996 3850 47048
rect 4798 47036 4804 47048
rect 4759 47008 4804 47036
rect 4798 46996 4804 47008
rect 4856 46996 4862 47048
rect 5537 47039 5595 47045
rect 5537 47005 5549 47039
rect 5583 47036 5595 47039
rect 5810 47036 5816 47048
rect 5583 47008 5816 47036
rect 5583 47005 5595 47008
rect 5537 46999 5595 47005
rect 5810 46996 5816 47008
rect 5868 46996 5874 47048
rect 6362 47036 6368 47048
rect 6323 47008 6368 47036
rect 6362 46996 6368 47008
rect 6420 46996 6426 47048
rect 7374 47036 7380 47048
rect 7335 47008 7380 47036
rect 7374 46996 7380 47008
rect 7432 46996 7438 47048
rect 8018 46996 8024 47048
rect 8076 47036 8082 47048
rect 8113 47039 8171 47045
rect 8113 47036 8125 47039
rect 8076 47008 8125 47036
rect 8076 46996 8082 47008
rect 8113 47005 8125 47008
rect 8159 47005 8171 47039
rect 8113 46999 8171 47005
rect 9677 47039 9735 47045
rect 9677 47005 9689 47039
rect 9723 47036 9735 47039
rect 9766 47036 9772 47048
rect 9723 47008 9772 47036
rect 9723 47005 9735 47008
rect 9677 46999 9735 47005
rect 9766 46996 9772 47008
rect 9824 46996 9830 47048
rect 10594 46996 10600 47048
rect 10652 47036 10658 47048
rect 10689 47039 10747 47045
rect 10689 47036 10701 47039
rect 10652 47008 10701 47036
rect 10652 46996 10658 47008
rect 10689 47005 10701 47008
rect 10735 47005 10747 47039
rect 10689 46999 10747 47005
rect 12161 47039 12219 47045
rect 12161 47005 12173 47039
rect 12207 47036 12219 47039
rect 12894 47036 12900 47048
rect 12207 47008 12900 47036
rect 12207 47005 12219 47008
rect 12161 46999 12219 47005
rect 12894 46996 12900 47008
rect 12952 46996 12958 47048
rect 13078 46996 13084 47048
rect 13136 47036 13142 47048
rect 13173 47039 13231 47045
rect 13173 47036 13185 47039
rect 13136 47008 13185 47036
rect 13136 46996 13142 47008
rect 13173 47005 13185 47008
rect 13219 47005 13231 47039
rect 14366 47036 14372 47048
rect 14327 47008 14372 47036
rect 13173 46999 13231 47005
rect 14366 46996 14372 47008
rect 14424 46996 14430 47048
rect 15654 47036 15660 47048
rect 15615 47008 15660 47036
rect 15654 46996 15660 47008
rect 15712 46996 15718 47048
rect 17221 47039 17279 47045
rect 17221 47005 17233 47039
rect 17267 47036 17279 47039
rect 17770 47036 17776 47048
rect 17267 47008 17776 47036
rect 17267 47005 17279 47008
rect 17221 46999 17279 47005
rect 17770 46996 17776 47008
rect 17828 46996 17834 47048
rect 18414 47036 18420 47048
rect 18375 47008 18420 47036
rect 18414 46996 18420 47008
rect 18472 46996 18478 47048
rect 19705 47039 19763 47045
rect 19705 47005 19717 47039
rect 19751 47036 19763 47039
rect 20438 47036 20444 47048
rect 19751 47008 20444 47036
rect 19751 47005 19763 47008
rect 19705 46999 19763 47005
rect 20438 46996 20444 47008
rect 20496 46996 20502 47048
rect 20622 47036 20628 47048
rect 20583 47008 20628 47036
rect 20622 46996 20628 47008
rect 20680 46996 20686 47048
rect 21910 47036 21916 47048
rect 21871 47008 21916 47036
rect 21910 46996 21916 47008
rect 21968 46996 21974 47048
rect 23106 47036 23112 47048
rect 23067 47008 23112 47036
rect 23106 46996 23112 47008
rect 23164 46996 23170 47048
rect 24394 47036 24400 47048
rect 24355 47008 24400 47036
rect 24394 46996 24400 47008
rect 24452 46996 24458 47048
rect 25682 47036 25688 47048
rect 25643 47008 25688 47036
rect 25682 46996 25688 47008
rect 25740 46996 25746 47048
rect 26970 47036 26976 47048
rect 26931 47008 26976 47036
rect 26970 46996 26976 47008
rect 27028 46996 27034 47048
rect 28166 47036 28172 47048
rect 28127 47008 28172 47036
rect 28166 46996 28172 47008
rect 28224 46996 28230 47048
rect 29546 47036 29552 47048
rect 29507 47008 29552 47036
rect 29546 46996 29552 47008
rect 29604 46996 29610 47048
rect 30650 47036 30656 47048
rect 30611 47008 30656 47036
rect 30650 46996 30656 47008
rect 30708 46996 30714 47048
rect 32398 47036 32404 47048
rect 32359 47008 32404 47036
rect 32398 46996 32404 47008
rect 32456 46996 32462 47048
rect 33410 47036 33416 47048
rect 33371 47008 33416 47036
rect 33410 46996 33416 47008
rect 33468 46996 33474 47048
rect 33873 47039 33931 47045
rect 33873 47005 33885 47039
rect 33919 47005 33931 47039
rect 34698 47036 34704 47048
rect 34659 47008 34704 47036
rect 33873 46999 33931 47005
rect 8938 46928 8944 46980
rect 8996 46968 9002 46980
rect 10229 46971 10287 46977
rect 10229 46968 10241 46971
rect 8996 46940 10241 46968
rect 8996 46928 9002 46940
rect 10229 46937 10241 46940
rect 10275 46968 10287 46971
rect 12621 46971 12679 46977
rect 12621 46968 12633 46971
rect 10275 46940 12633 46968
rect 10275 46937 10287 46940
rect 10229 46931 10287 46937
rect 12621 46937 12633 46940
rect 12667 46937 12679 46971
rect 15194 46968 15200 46980
rect 15155 46940 15200 46968
rect 12621 46931 12679 46937
rect 15194 46928 15200 46940
rect 15252 46928 15258 46980
rect 33134 46928 33140 46980
rect 33192 46968 33198 46980
rect 33888 46968 33916 46999
rect 34698 46996 34704 47008
rect 34756 46996 34762 47048
rect 35618 47036 35624 47048
rect 35579 47008 35624 47036
rect 35618 46996 35624 47008
rect 35676 46996 35682 47048
rect 36357 47039 36415 47045
rect 36357 47005 36369 47039
rect 36403 47005 36415 47039
rect 37550 47036 37556 47048
rect 37511 47008 37556 47036
rect 36357 46999 36415 47005
rect 33192 46940 33916 46968
rect 33192 46928 33198 46940
rect 34606 46928 34612 46980
rect 34664 46968 34670 46980
rect 36372 46968 36400 46999
rect 37550 46996 37556 47008
rect 37608 46996 37614 47048
rect 38381 47039 38439 47045
rect 38381 47005 38393 47039
rect 38427 47036 38439 47039
rect 38654 47036 38660 47048
rect 38427 47008 38660 47036
rect 38427 47005 38439 47008
rect 38381 46999 38439 47005
rect 38654 46996 38660 47008
rect 38712 46996 38718 47048
rect 38746 46996 38752 47048
rect 38804 47036 38810 47048
rect 38841 47039 38899 47045
rect 38841 47036 38853 47039
rect 38804 47008 38853 47036
rect 38804 46996 38810 47008
rect 38841 47005 38853 47008
rect 38887 47005 38899 47039
rect 39850 47036 39856 47048
rect 39811 47008 39856 47036
rect 38841 46999 38899 47005
rect 39850 46996 39856 47008
rect 39908 46996 39914 47048
rect 40865 47039 40923 47045
rect 40865 47005 40877 47039
rect 40911 47036 40923 47039
rect 41138 47036 41144 47048
rect 40911 47008 41144 47036
rect 40911 47005 40923 47008
rect 40865 46999 40923 47005
rect 41138 46996 41144 47008
rect 41196 46996 41202 47048
rect 41322 47036 41328 47048
rect 41283 47008 41328 47036
rect 41322 46996 41328 47008
rect 41380 46996 41386 47048
rect 41874 46996 41880 47048
rect 41932 47036 41938 47048
rect 42429 47039 42487 47045
rect 42429 47036 42441 47039
rect 41932 47008 42441 47036
rect 41932 46996 41938 47008
rect 42429 47005 42441 47008
rect 42475 47005 42487 47039
rect 43162 47036 43168 47048
rect 43123 47008 43168 47036
rect 42429 46999 42487 47005
rect 43162 46996 43168 47008
rect 43220 46996 43226 47048
rect 44174 47036 44180 47048
rect 44135 47008 44180 47036
rect 44174 46996 44180 47008
rect 44232 46996 44238 47048
rect 46032 47045 46060 47076
rect 47872 47045 47900 47076
rect 45281 47039 45339 47045
rect 45281 47005 45293 47039
rect 45327 47005 45339 47039
rect 45281 46999 45339 47005
rect 46017 47039 46075 47045
rect 46017 47005 46029 47039
rect 46063 47005 46075 47039
rect 46017 46999 46075 47005
rect 46753 47039 46811 47045
rect 46753 47005 46765 47039
rect 46799 47005 46811 47039
rect 46753 46999 46811 47005
rect 47857 47039 47915 47045
rect 47857 47005 47869 47039
rect 47903 47036 47915 47039
rect 47946 47036 47952 47048
rect 47903 47008 47952 47036
rect 47903 47005 47915 47008
rect 47857 46999 47915 47005
rect 34664 46940 36400 46968
rect 34664 46928 34670 46940
rect 42702 46928 42708 46980
rect 42760 46968 42766 46980
rect 45296 46968 45324 46999
rect 42760 46940 45324 46968
rect 42760 46928 42766 46940
rect 45738 46928 45744 46980
rect 45796 46968 45802 46980
rect 46768 46968 46796 46999
rect 47946 46996 47952 47008
rect 48004 46996 48010 47048
rect 45796 46940 46796 46968
rect 45796 46928 45802 46940
rect 1026 46860 1032 46912
rect 1084 46900 1090 46912
rect 3053 46903 3111 46909
rect 3053 46900 3065 46903
rect 1084 46872 3065 46900
rect 1084 46860 1090 46872
rect 3053 46869 3065 46872
rect 3099 46869 3111 46903
rect 3053 46863 3111 46869
rect 28810 46860 28816 46912
rect 28868 46900 28874 46912
rect 28905 46903 28963 46909
rect 28905 46900 28917 46903
rect 28868 46872 28917 46900
rect 28868 46860 28874 46872
rect 28905 46869 28917 46872
rect 28951 46869 28963 46903
rect 28905 46863 28963 46869
rect 31294 46860 31300 46912
rect 31352 46900 31358 46912
rect 31389 46903 31447 46909
rect 31389 46900 31401 46903
rect 31352 46872 31401 46900
rect 31352 46860 31358 46872
rect 31389 46869 31401 46872
rect 31435 46869 31447 46903
rect 31389 46863 31447 46869
rect 34790 46860 34796 46912
rect 34848 46900 34854 46912
rect 36541 46903 36599 46909
rect 36541 46900 36553 46903
rect 34848 46872 36553 46900
rect 34848 46860 34854 46872
rect 36541 46869 36553 46872
rect 36587 46869 36599 46903
rect 36541 46863 36599 46869
rect 36814 46860 36820 46912
rect 36872 46900 36878 46912
rect 37369 46903 37427 46909
rect 37369 46900 37381 46903
rect 36872 46872 37381 46900
rect 36872 46860 36878 46872
rect 37369 46869 37381 46872
rect 37415 46869 37427 46903
rect 37369 46863 37427 46869
rect 40954 46860 40960 46912
rect 41012 46900 41018 46912
rect 41509 46903 41567 46909
rect 41509 46900 41521 46903
rect 41012 46872 41521 46900
rect 41012 46860 41018 46872
rect 41509 46869 41521 46872
rect 41555 46869 41567 46903
rect 41509 46863 41567 46869
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 566 46656 572 46708
rect 624 46696 630 46708
rect 1489 46699 1547 46705
rect 1489 46696 1501 46699
rect 624 46668 1501 46696
rect 624 46656 630 46668
rect 1489 46665 1501 46668
rect 1535 46665 1547 46699
rect 1489 46659 1547 46665
rect 2222 46656 2228 46708
rect 2280 46696 2286 46708
rect 2409 46699 2467 46705
rect 2409 46696 2421 46699
rect 2280 46668 2421 46696
rect 2280 46656 2286 46668
rect 2409 46665 2421 46668
rect 2455 46665 2467 46699
rect 2409 46659 2467 46665
rect 3510 46656 3516 46708
rect 3568 46696 3574 46708
rect 4341 46699 4399 46705
rect 4341 46696 4353 46699
rect 3568 46668 4353 46696
rect 3568 46656 3574 46668
rect 4341 46665 4353 46668
rect 4387 46665 4399 46699
rect 4341 46659 4399 46665
rect 4798 46656 4804 46708
rect 4856 46696 4862 46708
rect 4893 46699 4951 46705
rect 4893 46696 4905 46699
rect 4856 46668 4905 46696
rect 4856 46656 4862 46668
rect 4893 46665 4905 46668
rect 4939 46665 4951 46699
rect 4893 46659 4951 46665
rect 5721 46699 5779 46705
rect 5721 46665 5733 46699
rect 5767 46696 5779 46699
rect 6362 46696 6368 46708
rect 5767 46668 6368 46696
rect 5767 46665 5779 46668
rect 5721 46659 5779 46665
rect 6362 46656 6368 46668
rect 6420 46656 6426 46708
rect 7190 46656 7196 46708
rect 7248 46696 7254 46708
rect 7377 46699 7435 46705
rect 7377 46696 7389 46699
rect 7248 46668 7389 46696
rect 7248 46656 7254 46668
rect 7377 46665 7389 46668
rect 7423 46665 7435 46699
rect 7377 46659 7435 46665
rect 8478 46656 8484 46708
rect 8536 46696 8542 46708
rect 8757 46699 8815 46705
rect 8757 46696 8769 46699
rect 8536 46668 8769 46696
rect 8536 46656 8542 46668
rect 8757 46665 8769 46668
rect 8803 46665 8815 46699
rect 8757 46659 8815 46665
rect 9858 46656 9864 46708
rect 9916 46696 9922 46708
rect 9953 46699 10011 46705
rect 9953 46696 9965 46699
rect 9916 46668 9965 46696
rect 9916 46656 9922 46668
rect 9953 46665 9965 46668
rect 9999 46665 10011 46699
rect 9953 46659 10011 46665
rect 10781 46699 10839 46705
rect 10781 46665 10793 46699
rect 10827 46696 10839 46699
rect 10962 46696 10968 46708
rect 10827 46668 10968 46696
rect 10827 46665 10839 46668
rect 10781 46659 10839 46665
rect 10962 46656 10968 46668
rect 11020 46656 11026 46708
rect 12253 46699 12311 46705
rect 12253 46665 12265 46699
rect 12299 46665 12311 46699
rect 12253 46659 12311 46665
rect 12268 46628 12296 46659
rect 12342 46656 12348 46708
rect 12400 46696 12406 46708
rect 12989 46699 13047 46705
rect 12989 46696 13001 46699
rect 12400 46668 13001 46696
rect 12400 46656 12406 46668
rect 12989 46665 13001 46668
rect 13035 46665 13047 46699
rect 12989 46659 13047 46665
rect 13446 46656 13452 46708
rect 13504 46696 13510 46708
rect 13633 46699 13691 46705
rect 13633 46696 13645 46699
rect 13504 46668 13645 46696
rect 13504 46656 13510 46668
rect 13633 46665 13645 46668
rect 13679 46665 13691 46699
rect 13633 46659 13691 46665
rect 14734 46656 14740 46708
rect 14792 46696 14798 46708
rect 14921 46699 14979 46705
rect 14921 46696 14933 46699
rect 14792 46668 14933 46696
rect 14792 46656 14798 46668
rect 14921 46665 14933 46668
rect 14967 46665 14979 46699
rect 15930 46696 15936 46708
rect 15891 46668 15936 46696
rect 14921 46659 14979 46665
rect 15930 46656 15936 46668
rect 15988 46656 15994 46708
rect 17218 46656 17224 46708
rect 17276 46696 17282 46708
rect 18141 46699 18199 46705
rect 18141 46696 18153 46699
rect 17276 46668 18153 46696
rect 17276 46656 17282 46668
rect 18141 46665 18153 46668
rect 18187 46665 18199 46699
rect 18141 46659 18199 46665
rect 18506 46656 18512 46708
rect 18564 46696 18570 46708
rect 18877 46699 18935 46705
rect 18877 46696 18889 46699
rect 18564 46668 18889 46696
rect 18564 46656 18570 46668
rect 18877 46665 18889 46668
rect 18923 46665 18935 46699
rect 19978 46696 19984 46708
rect 19939 46668 19984 46696
rect 18877 46659 18935 46665
rect 19978 46656 19984 46668
rect 20036 46656 20042 46708
rect 20438 46656 20444 46708
rect 20496 46696 20502 46708
rect 20533 46699 20591 46705
rect 20533 46696 20545 46699
rect 20496 46668 20545 46696
rect 20496 46656 20502 46668
rect 20533 46665 20545 46668
rect 20579 46665 20591 46699
rect 20533 46659 20591 46665
rect 20990 46656 20996 46708
rect 21048 46696 21054 46708
rect 22005 46699 22063 46705
rect 22005 46696 22017 46699
rect 21048 46668 22017 46696
rect 21048 46656 21054 46668
rect 22005 46665 22017 46668
rect 22051 46665 22063 46699
rect 22005 46659 22063 46665
rect 22186 46656 22192 46708
rect 22244 46696 22250 46708
rect 22741 46699 22799 46705
rect 22741 46696 22753 46699
rect 22244 46668 22753 46696
rect 22244 46656 22250 46668
rect 22741 46665 22753 46668
rect 22787 46665 22799 46699
rect 22741 46659 22799 46665
rect 23474 46656 23480 46708
rect 23532 46696 23538 46708
rect 24305 46699 24363 46705
rect 24305 46696 24317 46699
rect 23532 46668 24317 46696
rect 23532 46656 23538 46668
rect 24305 46665 24317 46668
rect 24351 46665 24363 46699
rect 24305 46659 24363 46665
rect 24670 46656 24676 46708
rect 24728 46696 24734 46708
rect 25041 46699 25099 46705
rect 25041 46696 25053 46699
rect 24728 46668 25053 46696
rect 24728 46656 24734 46668
rect 25041 46665 25053 46668
rect 25087 46665 25099 46699
rect 25041 46659 25099 46665
rect 25958 46656 25964 46708
rect 26016 46696 26022 46708
rect 26145 46699 26203 46705
rect 26145 46696 26157 46699
rect 26016 46668 26157 46696
rect 26016 46656 26022 46668
rect 26145 46665 26157 46668
rect 26191 46665 26203 46699
rect 26145 46659 26203 46665
rect 27246 46656 27252 46708
rect 27304 46696 27310 46708
rect 28261 46699 28319 46705
rect 28261 46696 28273 46699
rect 27304 46668 28273 46696
rect 27304 46656 27310 46668
rect 28261 46665 28273 46668
rect 28307 46665 28319 46699
rect 28261 46659 28319 46665
rect 29730 46656 29736 46708
rect 29788 46696 29794 46708
rect 30009 46699 30067 46705
rect 30009 46696 30021 46699
rect 29788 46668 30021 46696
rect 29788 46656 29794 46668
rect 30009 46665 30021 46668
rect 30055 46665 30067 46699
rect 30009 46659 30067 46665
rect 32398 46656 32404 46708
rect 32456 46696 32462 46708
rect 33045 46699 33103 46705
rect 33045 46696 33057 46699
rect 32456 46668 33057 46696
rect 32456 46656 32462 46668
rect 33045 46665 33057 46668
rect 33091 46665 33103 46699
rect 33045 46659 33103 46665
rect 33410 46656 33416 46708
rect 33468 46696 33474 46708
rect 33689 46699 33747 46705
rect 33689 46696 33701 46699
rect 33468 46668 33701 46696
rect 33468 46656 33474 46668
rect 33689 46665 33701 46668
rect 33735 46665 33747 46699
rect 33689 46659 33747 46665
rect 34517 46699 34575 46705
rect 34517 46665 34529 46699
rect 34563 46696 34575 46699
rect 34698 46696 34704 46708
rect 34563 46668 34704 46696
rect 34563 46665 34575 46668
rect 34517 46659 34575 46665
rect 34698 46656 34704 46668
rect 34756 46656 34762 46708
rect 35986 46656 35992 46708
rect 36044 46696 36050 46708
rect 36173 46699 36231 46705
rect 36173 46696 36185 46699
rect 36044 46668 36185 46696
rect 36044 46656 36050 46668
rect 36173 46665 36185 46668
rect 36219 46665 36231 46699
rect 36173 46659 36231 46665
rect 37182 46656 37188 46708
rect 37240 46696 37246 46708
rect 37461 46699 37519 46705
rect 37461 46696 37473 46699
rect 37240 46668 37473 46696
rect 37240 46656 37246 46668
rect 37461 46665 37473 46668
rect 37507 46665 37519 46699
rect 37461 46659 37519 46665
rect 37550 46656 37556 46708
rect 37608 46696 37614 46708
rect 38013 46699 38071 46705
rect 38013 46696 38025 46699
rect 37608 46668 38025 46696
rect 37608 46656 37614 46668
rect 38013 46665 38025 46668
rect 38059 46665 38071 46699
rect 38654 46696 38660 46708
rect 38615 46668 38660 46696
rect 38013 46659 38071 46665
rect 38654 46656 38660 46668
rect 38712 46656 38718 46708
rect 39666 46656 39672 46708
rect 39724 46696 39730 46708
rect 39945 46699 40003 46705
rect 39945 46696 39957 46699
rect 39724 46668 39957 46696
rect 39724 46656 39730 46668
rect 39945 46665 39957 46668
rect 39991 46665 40003 46699
rect 39945 46659 40003 46665
rect 42242 46656 42248 46708
rect 42300 46696 42306 46708
rect 42613 46699 42671 46705
rect 42613 46696 42625 46699
rect 42300 46668 42625 46696
rect 42300 46656 42306 46668
rect 42613 46665 42625 46668
rect 42659 46665 42671 46699
rect 42613 46659 42671 46665
rect 43438 46656 43444 46708
rect 43496 46696 43502 46708
rect 43717 46699 43775 46705
rect 43717 46696 43729 46699
rect 43496 46668 43729 46696
rect 43496 46656 43502 46668
rect 43717 46665 43729 46668
rect 43763 46665 43775 46699
rect 44726 46696 44732 46708
rect 44687 46668 44732 46696
rect 43717 46659 43775 46665
rect 44726 46656 44732 46668
rect 44784 46656 44790 46708
rect 45465 46699 45523 46705
rect 45465 46665 45477 46699
rect 45511 46665 45523 46699
rect 46198 46696 46204 46708
rect 46159 46668 46204 46696
rect 45465 46659 45523 46665
rect 32030 46628 32036 46640
rect 12268 46600 32036 46628
rect 32030 46588 32036 46600
rect 32088 46588 32094 46640
rect 32125 46631 32183 46637
rect 32125 46597 32137 46631
rect 32171 46628 32183 46631
rect 41046 46628 41052 46640
rect 32171 46600 41052 46628
rect 32171 46597 32183 46600
rect 32125 46591 32183 46597
rect 41046 46588 41052 46600
rect 41104 46588 41110 46640
rect 41138 46588 41144 46640
rect 41196 46588 41202 46640
rect 45480 46628 45508 46659
rect 46198 46656 46204 46668
rect 46256 46656 46262 46708
rect 46937 46699 46995 46705
rect 46937 46665 46949 46699
rect 46983 46696 46995 46699
rect 48866 46696 48872 46708
rect 46983 46668 48872 46696
rect 46983 46665 46995 46668
rect 46937 46659 46995 46665
rect 48866 46656 48872 46668
rect 48924 46656 48930 46708
rect 48038 46628 48044 46640
rect 45480 46600 48044 46628
rect 48038 46588 48044 46600
rect 48096 46588 48102 46640
rect 1673 46563 1731 46569
rect 1673 46529 1685 46563
rect 1719 46560 1731 46563
rect 2498 46560 2504 46572
rect 1719 46532 2504 46560
rect 1719 46529 1731 46532
rect 1673 46523 1731 46529
rect 2498 46520 2504 46532
rect 2556 46520 2562 46572
rect 2590 46520 2596 46572
rect 2648 46560 2654 46572
rect 2648 46532 2693 46560
rect 2648 46520 2654 46532
rect 3050 46520 3056 46572
rect 3108 46560 3114 46572
rect 3421 46563 3479 46569
rect 3421 46560 3433 46563
rect 3108 46532 3433 46560
rect 3108 46520 3114 46532
rect 3421 46529 3433 46532
rect 3467 46529 3479 46563
rect 4154 46560 4160 46572
rect 4115 46532 4160 46560
rect 3421 46523 3479 46529
rect 4154 46520 4160 46532
rect 4212 46520 4218 46572
rect 5077 46563 5135 46569
rect 5077 46529 5089 46563
rect 5123 46560 5135 46563
rect 5537 46563 5595 46569
rect 5537 46560 5549 46563
rect 5123 46532 5549 46560
rect 5123 46529 5135 46532
rect 5077 46523 5135 46529
rect 5537 46529 5549 46532
rect 5583 46529 5595 46563
rect 6362 46560 6368 46572
rect 6323 46532 6368 46560
rect 5537 46523 5595 46529
rect 5552 46492 5580 46523
rect 6362 46520 6368 46532
rect 6420 46520 6426 46572
rect 7561 46563 7619 46569
rect 7561 46529 7573 46563
rect 7607 46560 7619 46563
rect 7742 46560 7748 46572
rect 7607 46532 7748 46560
rect 7607 46529 7619 46532
rect 7561 46523 7619 46529
rect 7742 46520 7748 46532
rect 7800 46520 7806 46572
rect 8110 46520 8116 46572
rect 8168 46560 8174 46572
rect 8573 46563 8631 46569
rect 8573 46560 8585 46563
rect 8168 46532 8585 46560
rect 8168 46520 8174 46532
rect 8573 46529 8585 46532
rect 8619 46529 8631 46563
rect 8573 46523 8631 46529
rect 9858 46520 9864 46572
rect 9916 46560 9922 46572
rect 10137 46563 10195 46569
rect 10137 46560 10149 46563
rect 9916 46532 10149 46560
rect 9916 46520 9922 46532
rect 10137 46529 10149 46532
rect 10183 46529 10195 46563
rect 10137 46523 10195 46529
rect 10965 46563 11023 46569
rect 10965 46529 10977 46563
rect 11011 46560 11023 46563
rect 11698 46560 11704 46572
rect 11011 46532 11704 46560
rect 11011 46529 11023 46532
rect 10965 46523 11023 46529
rect 11698 46520 11704 46532
rect 11756 46520 11762 46572
rect 12069 46563 12127 46569
rect 12069 46529 12081 46563
rect 12115 46529 12127 46563
rect 12802 46560 12808 46572
rect 12763 46532 12808 46560
rect 12069 46523 12127 46529
rect 12084 46492 12112 46523
rect 12802 46520 12808 46532
rect 12860 46520 12866 46572
rect 13814 46560 13820 46572
rect 13775 46532 13820 46560
rect 13814 46520 13820 46532
rect 13872 46520 13878 46572
rect 15102 46560 15108 46572
rect 15063 46532 15108 46560
rect 15102 46520 15108 46532
rect 15160 46520 15166 46572
rect 15930 46520 15936 46572
rect 15988 46560 15994 46572
rect 16117 46563 16175 46569
rect 16117 46560 16129 46563
rect 15988 46532 16129 46560
rect 15988 46520 15994 46532
rect 16117 46529 16129 46532
rect 16163 46529 16175 46563
rect 16117 46523 16175 46529
rect 16666 46520 16672 46572
rect 16724 46560 16730 46572
rect 17313 46563 17371 46569
rect 17313 46560 17325 46563
rect 16724 46532 17325 46560
rect 16724 46520 16730 46532
rect 17313 46529 17325 46532
rect 17359 46529 17371 46563
rect 17954 46560 17960 46572
rect 17915 46532 17960 46560
rect 17313 46523 17371 46529
rect 17954 46520 17960 46532
rect 18012 46520 18018 46572
rect 18690 46560 18696 46572
rect 18651 46532 18696 46560
rect 18690 46520 18696 46532
rect 18748 46520 18754 46572
rect 19797 46563 19855 46569
rect 19797 46529 19809 46563
rect 19843 46560 19855 46563
rect 19978 46560 19984 46572
rect 19843 46532 19984 46560
rect 19843 46529 19855 46532
rect 19797 46523 19855 46529
rect 19978 46520 19984 46532
rect 20036 46520 20042 46572
rect 20714 46560 20720 46572
rect 20675 46532 20720 46560
rect 20714 46520 20720 46532
rect 20772 46520 20778 46572
rect 21082 46520 21088 46572
rect 21140 46560 21146 46572
rect 21821 46563 21879 46569
rect 21821 46560 21833 46563
rect 21140 46532 21833 46560
rect 21140 46520 21146 46532
rect 21821 46529 21833 46532
rect 21867 46529 21879 46563
rect 22554 46560 22560 46572
rect 22515 46532 22560 46560
rect 21821 46523 21879 46529
rect 22554 46520 22560 46532
rect 22612 46520 22618 46572
rect 23014 46520 23020 46572
rect 23072 46560 23078 46572
rect 23477 46563 23535 46569
rect 23477 46560 23489 46563
rect 23072 46532 23489 46560
rect 23072 46520 23078 46532
rect 23477 46529 23489 46532
rect 23523 46529 23535 46563
rect 23477 46523 23535 46529
rect 23750 46520 23756 46572
rect 23808 46560 23814 46572
rect 24121 46563 24179 46569
rect 24121 46560 24133 46563
rect 23808 46532 24133 46560
rect 23808 46520 23814 46532
rect 24121 46529 24133 46532
rect 24167 46529 24179 46563
rect 24121 46523 24179 46529
rect 24857 46563 24915 46569
rect 24857 46529 24869 46563
rect 24903 46560 24915 46563
rect 24946 46560 24952 46572
rect 24903 46532 24952 46560
rect 24903 46529 24915 46532
rect 24857 46523 24915 46529
rect 24946 46520 24952 46532
rect 25004 46520 25010 46572
rect 26234 46520 26240 46572
rect 26292 46560 26298 46572
rect 26329 46563 26387 46569
rect 26329 46560 26341 46563
rect 26292 46532 26341 46560
rect 26292 46520 26298 46532
rect 26329 46529 26341 46532
rect 26375 46529 26387 46563
rect 27430 46560 27436 46572
rect 27391 46532 27436 46560
rect 26329 46523 26387 46529
rect 27430 46520 27436 46532
rect 27488 46520 27494 46572
rect 27522 46520 27528 46572
rect 27580 46560 27586 46572
rect 28077 46563 28135 46569
rect 28077 46560 28089 46563
rect 27580 46532 28089 46560
rect 27580 46520 27586 46532
rect 28077 46529 28089 46532
rect 28123 46529 28135 46563
rect 28077 46523 28135 46529
rect 28810 46520 28816 46572
rect 28868 46560 28874 46572
rect 28905 46563 28963 46569
rect 28905 46560 28917 46563
rect 28868 46532 28917 46560
rect 28868 46520 28874 46532
rect 28905 46529 28917 46532
rect 28951 46529 28963 46563
rect 29822 46560 29828 46572
rect 29783 46532 29828 46560
rect 28905 46523 28963 46529
rect 29822 46520 29828 46532
rect 29880 46520 29886 46572
rect 31113 46563 31171 46569
rect 31113 46529 31125 46563
rect 31159 46560 31171 46563
rect 31294 46560 31300 46572
rect 31159 46532 31300 46560
rect 31159 46529 31171 46532
rect 31113 46523 31171 46529
rect 31294 46520 31300 46532
rect 31352 46520 31358 46572
rect 31754 46520 31760 46572
rect 31812 46560 31818 46572
rect 32309 46563 32367 46569
rect 32309 46560 32321 46563
rect 31812 46532 32321 46560
rect 31812 46520 31818 46532
rect 32309 46529 32321 46532
rect 32355 46529 32367 46563
rect 32309 46523 32367 46529
rect 33229 46563 33287 46569
rect 33229 46529 33241 46563
rect 33275 46560 33287 46563
rect 33873 46563 33931 46569
rect 33873 46560 33885 46563
rect 33275 46532 33885 46560
rect 33275 46529 33287 46532
rect 33229 46523 33287 46529
rect 33873 46529 33885 46532
rect 33919 46560 33931 46563
rect 34330 46560 34336 46572
rect 33919 46532 34336 46560
rect 33919 46529 33931 46532
rect 33873 46523 33931 46529
rect 34330 46520 34336 46532
rect 34388 46520 34394 46572
rect 34790 46520 34796 46572
rect 34848 46560 34854 46572
rect 35069 46563 35127 46569
rect 35069 46560 35081 46563
rect 34848 46532 35081 46560
rect 34848 46520 34854 46532
rect 35069 46529 35081 46532
rect 35115 46529 35127 46563
rect 35069 46523 35127 46529
rect 36262 46520 36268 46572
rect 36320 46560 36326 46572
rect 36357 46563 36415 46569
rect 36357 46560 36369 46563
rect 36320 46532 36369 46560
rect 36320 46520 36326 46532
rect 36357 46529 36369 46532
rect 36403 46529 36415 46563
rect 36357 46523 36415 46529
rect 37277 46563 37335 46569
rect 37277 46529 37289 46563
rect 37323 46560 37335 46563
rect 37366 46560 37372 46572
rect 37323 46532 37372 46560
rect 37323 46529 37335 46532
rect 37277 46523 37335 46529
rect 37366 46520 37372 46532
rect 37424 46520 37430 46572
rect 38197 46563 38255 46569
rect 38197 46529 38209 46563
rect 38243 46560 38255 46563
rect 38841 46563 38899 46569
rect 38841 46560 38853 46563
rect 38243 46532 38853 46560
rect 38243 46529 38255 46532
rect 38197 46523 38255 46529
rect 38841 46529 38853 46532
rect 38887 46560 38899 46563
rect 39114 46560 39120 46572
rect 38887 46532 39120 46560
rect 38887 46529 38899 46532
rect 38841 46523 38899 46529
rect 39114 46520 39120 46532
rect 39172 46520 39178 46572
rect 39758 46560 39764 46572
rect 39719 46532 39764 46560
rect 39758 46520 39764 46532
rect 39816 46520 39822 46572
rect 40494 46560 40500 46572
rect 40455 46532 40500 46560
rect 40494 46520 40500 46532
rect 40552 46520 40558 46572
rect 5552 46464 8156 46492
rect 5994 46384 6000 46436
rect 6052 46424 6058 46436
rect 6549 46427 6607 46433
rect 6549 46424 6561 46427
rect 6052 46396 6561 46424
rect 6052 46384 6058 46396
rect 6549 46393 6561 46396
rect 6595 46393 6607 46427
rect 6549 46387 6607 46393
rect 3602 46356 3608 46368
rect 3563 46328 3608 46356
rect 3602 46316 3608 46328
rect 3660 46316 3666 46368
rect 8128 46365 8156 46464
rect 11532 46464 12112 46492
rect 21269 46495 21327 46501
rect 8113 46359 8171 46365
rect 8113 46325 8125 46359
rect 8159 46356 8171 46359
rect 9398 46356 9404 46368
rect 8159 46328 9404 46356
rect 8159 46325 8171 46328
rect 8113 46319 8171 46325
rect 9398 46316 9404 46328
rect 9456 46316 9462 46368
rect 11238 46316 11244 46368
rect 11296 46356 11302 46368
rect 11532 46365 11560 46464
rect 21269 46461 21281 46495
rect 21315 46492 21327 46495
rect 23032 46492 23060 46520
rect 21315 46464 23060 46492
rect 27617 46495 27675 46501
rect 21315 46461 21327 46464
rect 21269 46455 21327 46461
rect 27617 46461 27629 46495
rect 27663 46492 27675 46495
rect 40126 46492 40132 46504
rect 27663 46464 40132 46492
rect 27663 46461 27675 46464
rect 27617 46455 27675 46461
rect 40126 46452 40132 46464
rect 40184 46452 40190 46504
rect 17497 46427 17555 46433
rect 17497 46393 17509 46427
rect 17543 46424 17555 46427
rect 32125 46427 32183 46433
rect 32125 46424 32137 46427
rect 17543 46396 32137 46424
rect 17543 46393 17555 46396
rect 17497 46387 17555 46393
rect 32125 46393 32137 46396
rect 32171 46393 32183 46427
rect 32125 46387 32183 46393
rect 32214 46384 32220 46436
rect 32272 46424 32278 46436
rect 32493 46427 32551 46433
rect 32493 46424 32505 46427
rect 32272 46396 32505 46424
rect 32272 46384 32278 46396
rect 32493 46393 32505 46396
rect 32539 46393 32551 46427
rect 32493 46387 32551 46393
rect 35253 46427 35311 46433
rect 35253 46393 35265 46427
rect 35299 46424 35311 46427
rect 41046 46424 41052 46436
rect 35299 46396 41052 46424
rect 35299 46393 35311 46396
rect 35253 46387 35311 46393
rect 41046 46384 41052 46396
rect 41104 46384 41110 46436
rect 41156 46433 41184 46588
rect 41230 46520 41236 46572
rect 41288 46560 41294 46572
rect 41325 46563 41383 46569
rect 41325 46560 41337 46563
rect 41288 46532 41337 46560
rect 41288 46520 41294 46532
rect 41325 46529 41337 46532
rect 41371 46529 41383 46563
rect 41782 46560 41788 46572
rect 41743 46532 41788 46560
rect 41325 46523 41383 46529
rect 41782 46520 41788 46532
rect 41840 46520 41846 46572
rect 42426 46560 42432 46572
rect 42387 46532 42432 46560
rect 42426 46520 42432 46532
rect 42484 46520 42490 46572
rect 43530 46560 43536 46572
rect 43491 46532 43536 46560
rect 43530 46520 43536 46532
rect 43588 46520 43594 46572
rect 44542 46560 44548 46572
rect 44503 46532 44548 46560
rect 44542 46520 44548 46532
rect 44600 46520 44606 46572
rect 45278 46560 45284 46572
rect 45239 46532 45284 46560
rect 45278 46520 45284 46532
rect 45336 46520 45342 46572
rect 46014 46560 46020 46572
rect 45975 46532 46020 46560
rect 46014 46520 46020 46532
rect 46072 46520 46078 46572
rect 46753 46563 46811 46569
rect 46753 46529 46765 46563
rect 46799 46529 46811 46563
rect 47854 46560 47860 46572
rect 47815 46532 47860 46560
rect 46753 46523 46811 46529
rect 41141 46427 41199 46433
rect 41141 46393 41153 46427
rect 41187 46393 41199 46427
rect 41141 46387 41199 46393
rect 11517 46359 11575 46365
rect 11517 46356 11529 46359
rect 11296 46328 11529 46356
rect 11296 46316 11302 46328
rect 11517 46325 11529 46328
rect 11563 46325 11575 46359
rect 11517 46319 11575 46325
rect 14182 46316 14188 46368
rect 14240 46356 14246 46368
rect 14277 46359 14335 46365
rect 14277 46356 14289 46359
rect 14240 46328 14289 46356
rect 14240 46316 14246 46328
rect 14277 46325 14289 46328
rect 14323 46325 14335 46359
rect 16666 46356 16672 46368
rect 16627 46328 16672 46356
rect 14277 46319 14335 46325
rect 16666 46316 16672 46328
rect 16724 46316 16730 46368
rect 23569 46359 23627 46365
rect 23569 46325 23581 46359
rect 23615 46356 23627 46359
rect 24762 46356 24768 46368
rect 23615 46328 24768 46356
rect 23615 46325 23627 46328
rect 23569 46319 23627 46325
rect 24762 46316 24768 46328
rect 24820 46316 24826 46368
rect 28994 46356 29000 46368
rect 28955 46328 29000 46356
rect 28994 46316 29000 46328
rect 29052 46316 29058 46368
rect 31205 46359 31263 46365
rect 31205 46325 31217 46359
rect 31251 46356 31263 46359
rect 40034 46356 40040 46368
rect 31251 46328 40040 46356
rect 31251 46325 31263 46328
rect 31205 46319 31263 46325
rect 40034 46316 40040 46328
rect 40092 46316 40098 46368
rect 40681 46359 40739 46365
rect 40681 46325 40693 46359
rect 40727 46356 40739 46359
rect 42702 46356 42708 46368
rect 40727 46328 42708 46356
rect 40727 46325 40739 46328
rect 40681 46319 40739 46325
rect 42702 46316 42708 46328
rect 42760 46316 42766 46368
rect 45094 46316 45100 46368
rect 45152 46356 45158 46368
rect 46198 46356 46204 46368
rect 45152 46328 46204 46356
rect 45152 46316 45158 46328
rect 46198 46316 46204 46328
rect 46256 46356 46262 46368
rect 46768 46356 46796 46523
rect 47854 46520 47860 46532
rect 47912 46520 47918 46572
rect 48038 46424 48044 46436
rect 47999 46396 48044 46424
rect 48038 46384 48044 46396
rect 48096 46384 48102 46436
rect 46256 46328 46796 46356
rect 46256 46316 46262 46328
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 1670 46112 1676 46164
rect 1728 46152 1734 46164
rect 1949 46155 2007 46161
rect 1949 46152 1961 46155
rect 1728 46124 1961 46152
rect 1728 46112 1734 46124
rect 1949 46121 1961 46124
rect 1995 46121 2007 46155
rect 1949 46115 2007 46121
rect 2498 46112 2504 46164
rect 2556 46152 2562 46164
rect 2593 46155 2651 46161
rect 2593 46152 2605 46155
rect 2556 46124 2605 46152
rect 2556 46112 2562 46124
rect 2593 46121 2605 46124
rect 2639 46121 2651 46155
rect 3786 46152 3792 46164
rect 3747 46124 3792 46152
rect 2593 46115 2651 46121
rect 3786 46112 3792 46124
rect 3844 46112 3850 46164
rect 7374 46112 7380 46164
rect 7432 46152 7438 46164
rect 8205 46155 8263 46161
rect 8205 46152 8217 46155
rect 7432 46124 8217 46152
rect 7432 46112 7438 46124
rect 8205 46121 8217 46124
rect 8251 46121 8263 46155
rect 8205 46115 8263 46121
rect 12437 46155 12495 46161
rect 12437 46121 12449 46155
rect 12483 46152 12495 46155
rect 12802 46152 12808 46164
rect 12483 46124 12808 46152
rect 12483 46121 12495 46124
rect 12437 46115 12495 46121
rect 12802 46112 12808 46124
rect 12860 46112 12866 46164
rect 12894 46112 12900 46164
rect 12952 46152 12958 46164
rect 17770 46152 17776 46164
rect 12952 46124 12997 46152
rect 17731 46124 17776 46152
rect 12952 46112 12958 46124
rect 17770 46112 17776 46124
rect 17828 46112 17834 46164
rect 18414 46152 18420 46164
rect 18375 46124 18420 46152
rect 18414 46112 18420 46124
rect 18472 46112 18478 46164
rect 20533 46155 20591 46161
rect 20533 46121 20545 46155
rect 20579 46152 20591 46155
rect 20622 46152 20628 46164
rect 20579 46124 20628 46152
rect 20579 46121 20591 46124
rect 20533 46115 20591 46121
rect 20622 46112 20628 46124
rect 20680 46112 20686 46164
rect 21729 46155 21787 46161
rect 21729 46121 21741 46155
rect 21775 46152 21787 46155
rect 21910 46152 21916 46164
rect 21775 46124 21916 46152
rect 21775 46121 21787 46124
rect 21729 46115 21787 46121
rect 21910 46112 21916 46124
rect 21968 46112 21974 46164
rect 26881 46155 26939 46161
rect 22066 46124 25820 46152
rect 19889 46087 19947 46093
rect 19889 46053 19901 46087
rect 19935 46084 19947 46087
rect 22066 46084 22094 46124
rect 19935 46056 22094 46084
rect 25792 46084 25820 46124
rect 26881 46121 26893 46155
rect 26927 46152 26939 46155
rect 26970 46152 26976 46164
rect 26927 46124 26976 46152
rect 26927 46121 26939 46124
rect 26881 46115 26939 46121
rect 26970 46112 26976 46124
rect 27028 46112 27034 46164
rect 27985 46155 28043 46161
rect 27985 46121 27997 46155
rect 28031 46152 28043 46155
rect 28166 46152 28172 46164
rect 28031 46124 28172 46152
rect 28031 46121 28043 46124
rect 27985 46115 28043 46121
rect 28166 46112 28172 46124
rect 28224 46112 28230 46164
rect 28442 46112 28448 46164
rect 28500 46152 28506 46164
rect 28721 46155 28779 46161
rect 28721 46152 28733 46155
rect 28500 46124 28733 46152
rect 28500 46112 28506 46124
rect 28721 46121 28733 46124
rect 28767 46121 28779 46155
rect 29546 46152 29552 46164
rect 29507 46124 29552 46152
rect 28721 46115 28779 46121
rect 29546 46112 29552 46124
rect 29604 46112 29610 46164
rect 30561 46155 30619 46161
rect 30561 46121 30573 46155
rect 30607 46152 30619 46155
rect 30650 46152 30656 46164
rect 30607 46124 30656 46152
rect 30607 46121 30619 46124
rect 30561 46115 30619 46121
rect 30650 46112 30656 46124
rect 30708 46112 30714 46164
rect 30926 46112 30932 46164
rect 30984 46152 30990 46164
rect 31205 46155 31263 46161
rect 31205 46152 31217 46155
rect 30984 46124 31217 46152
rect 30984 46112 30990 46124
rect 31205 46121 31217 46124
rect 31251 46121 31263 46155
rect 31205 46115 31263 46121
rect 32030 46112 32036 46164
rect 32088 46152 32094 46164
rect 35434 46152 35440 46164
rect 32088 46124 35440 46152
rect 32088 46112 32094 46124
rect 35434 46112 35440 46124
rect 35492 46112 35498 46164
rect 35529 46155 35587 46161
rect 35529 46121 35541 46155
rect 35575 46152 35587 46155
rect 35618 46152 35624 46164
rect 35575 46124 35624 46152
rect 35575 46121 35587 46124
rect 35529 46115 35587 46121
rect 35618 46112 35624 46124
rect 35676 46112 35682 46164
rect 39114 46152 39120 46164
rect 35820 46124 39120 46152
rect 25792 46056 26924 46084
rect 19935 46053 19947 46056
rect 19889 46047 19947 46053
rect 1489 46019 1547 46025
rect 1489 45985 1501 46019
rect 1535 46016 1547 46019
rect 3050 46016 3056 46028
rect 1535 45988 3056 46016
rect 1535 45985 1547 45988
rect 1489 45979 1547 45985
rect 3050 45976 3056 45988
rect 3108 45976 3114 46028
rect 8938 46016 8944 46028
rect 7392 45988 8944 46016
rect 2038 45908 2044 45960
rect 2096 45948 2102 45960
rect 2133 45951 2191 45957
rect 2133 45948 2145 45951
rect 2096 45920 2145 45948
rect 2096 45908 2102 45920
rect 2133 45917 2145 45920
rect 2179 45917 2191 45951
rect 2133 45911 2191 45917
rect 2774 45908 2780 45960
rect 2832 45948 2838 45960
rect 3973 45951 4031 45957
rect 3973 45948 3985 45951
rect 2832 45920 3985 45948
rect 2832 45908 2838 45920
rect 3973 45917 3985 45920
rect 4019 45917 4031 45951
rect 3973 45911 4031 45917
rect 4433 45951 4491 45957
rect 4433 45917 4445 45951
rect 4479 45948 4491 45951
rect 6365 45951 6423 45957
rect 6365 45948 6377 45951
rect 4479 45920 6377 45948
rect 4479 45917 4491 45920
rect 4433 45911 4491 45917
rect 6365 45917 6377 45920
rect 6411 45948 6423 45951
rect 6914 45948 6920 45960
rect 6411 45920 6920 45948
rect 6411 45917 6423 45920
rect 6365 45911 6423 45917
rect 3988 45812 4016 45911
rect 6914 45908 6920 45920
rect 6972 45948 6978 45960
rect 7392 45948 7420 45988
rect 8938 45976 8944 45988
rect 8996 45976 9002 46028
rect 26896 46016 26924 46056
rect 28994 46044 29000 46096
rect 29052 46084 29058 46096
rect 31846 46084 31852 46096
rect 29052 46056 31852 46084
rect 29052 46044 29058 46056
rect 31846 46044 31852 46056
rect 31904 46044 31910 46096
rect 26896 45988 31754 46016
rect 8386 45948 8392 45960
rect 6972 45920 7420 45948
rect 8299 45920 8392 45948
rect 6972 45908 6978 45920
rect 8386 45908 8392 45920
rect 8444 45948 8450 45960
rect 11057 45951 11115 45957
rect 8444 45920 9444 45948
rect 8444 45908 8450 45920
rect 9416 45892 9444 45920
rect 11057 45917 11069 45951
rect 11103 45948 11115 45951
rect 11146 45948 11152 45960
rect 11103 45920 11152 45948
rect 11103 45917 11115 45920
rect 11057 45911 11115 45917
rect 11146 45908 11152 45920
rect 11204 45908 11210 45960
rect 13081 45951 13139 45957
rect 13081 45917 13093 45951
rect 13127 45917 13139 45951
rect 13081 45911 13139 45917
rect 14093 45951 14151 45957
rect 14093 45917 14105 45951
rect 14139 45948 14151 45951
rect 15194 45948 15200 45960
rect 14139 45920 15200 45948
rect 14139 45917 14151 45920
rect 14093 45911 14151 45917
rect 4700 45883 4758 45889
rect 4700 45849 4712 45883
rect 4746 45880 4758 45883
rect 5258 45880 5264 45892
rect 4746 45852 5264 45880
rect 4746 45849 4758 45852
rect 4700 45843 4758 45849
rect 5258 45840 5264 45852
rect 5316 45840 5322 45892
rect 6454 45840 6460 45892
rect 6512 45880 6518 45892
rect 6610 45883 6668 45889
rect 6610 45880 6622 45883
rect 6512 45852 6622 45880
rect 6512 45840 6518 45852
rect 6610 45849 6622 45852
rect 6656 45849 6668 45883
rect 6610 45843 6668 45849
rect 9208 45883 9266 45889
rect 9208 45849 9220 45883
rect 9254 45880 9266 45883
rect 9306 45880 9312 45892
rect 9254 45852 9312 45880
rect 9254 45849 9266 45852
rect 9208 45843 9266 45849
rect 9306 45840 9312 45852
rect 9364 45840 9370 45892
rect 9398 45840 9404 45892
rect 9456 45840 9462 45892
rect 11324 45883 11382 45889
rect 11324 45849 11336 45883
rect 11370 45880 11382 45883
rect 11514 45880 11520 45892
rect 11370 45852 11520 45880
rect 11370 45849 11382 45852
rect 11324 45843 11382 45849
rect 11514 45840 11520 45852
rect 11572 45840 11578 45892
rect 12894 45840 12900 45892
rect 12952 45880 12958 45892
rect 13096 45880 13124 45911
rect 15194 45908 15200 45920
rect 15252 45948 15258 45960
rect 15838 45948 15844 45960
rect 15252 45920 15844 45948
rect 15252 45908 15258 45920
rect 15838 45908 15844 45920
rect 15896 45948 15902 45960
rect 17313 45951 17371 45957
rect 17313 45948 17325 45951
rect 15896 45920 17325 45948
rect 15896 45908 15902 45920
rect 17313 45917 17325 45920
rect 17359 45948 17371 45951
rect 17402 45948 17408 45960
rect 17359 45920 17408 45948
rect 17359 45917 17371 45920
rect 17313 45911 17371 45917
rect 17402 45908 17408 45920
rect 17460 45908 17466 45960
rect 17957 45951 18015 45957
rect 17957 45917 17969 45951
rect 18003 45948 18015 45951
rect 18601 45951 18659 45957
rect 18601 45948 18613 45951
rect 18003 45920 18613 45948
rect 18003 45917 18015 45920
rect 17957 45911 18015 45917
rect 18601 45917 18613 45920
rect 18647 45948 18659 45951
rect 20349 45951 20407 45957
rect 20349 45948 20361 45951
rect 18647 45920 20361 45948
rect 18647 45917 18659 45920
rect 18601 45911 18659 45917
rect 20349 45917 20361 45920
rect 20395 45948 20407 45951
rect 20714 45948 20720 45960
rect 20395 45920 20720 45948
rect 20395 45917 20407 45920
rect 20349 45911 20407 45917
rect 20714 45908 20720 45920
rect 20772 45948 20778 45960
rect 21085 45951 21143 45957
rect 21085 45948 21097 45951
rect 20772 45920 21097 45948
rect 20772 45908 20778 45920
rect 21085 45917 21097 45920
rect 21131 45948 21143 45951
rect 21542 45948 21548 45960
rect 21131 45920 21548 45948
rect 21131 45917 21143 45920
rect 21085 45911 21143 45917
rect 21542 45908 21548 45920
rect 21600 45908 21606 45960
rect 22373 45951 22431 45957
rect 22373 45917 22385 45951
rect 22419 45948 22431 45951
rect 24854 45948 24860 45960
rect 22419 45920 24860 45948
rect 22419 45917 22431 45920
rect 22373 45911 22431 45917
rect 24854 45908 24860 45920
rect 24912 45908 24918 45960
rect 26697 45951 26755 45957
rect 26697 45917 26709 45951
rect 26743 45948 26755 45951
rect 26970 45948 26976 45960
rect 26743 45920 26976 45948
rect 26743 45917 26755 45920
rect 26697 45911 26755 45917
rect 26970 45908 26976 45920
rect 27028 45948 27034 45960
rect 27801 45951 27859 45957
rect 27801 45948 27813 45951
rect 27028 45920 27813 45948
rect 27028 45908 27034 45920
rect 27801 45917 27813 45920
rect 27847 45948 27859 45951
rect 28445 45951 28503 45957
rect 28445 45948 28457 45951
rect 27847 45920 28457 45948
rect 27847 45917 27859 45920
rect 27801 45911 27859 45917
rect 28445 45917 28457 45920
rect 28491 45917 28503 45951
rect 28445 45911 28503 45917
rect 28537 45951 28595 45957
rect 28537 45917 28549 45951
rect 28583 45917 28595 45951
rect 29730 45948 29736 45960
rect 29691 45920 29736 45948
rect 28537 45911 28595 45917
rect 14182 45880 14188 45892
rect 12952 45852 14188 45880
rect 12952 45840 12958 45852
rect 14182 45840 14188 45852
rect 14240 45840 14246 45892
rect 14360 45883 14418 45889
rect 14360 45849 14372 45883
rect 14406 45849 14418 45883
rect 14360 45843 14418 45849
rect 4982 45812 4988 45824
rect 3988 45784 4988 45812
rect 4982 45772 4988 45784
rect 5040 45772 5046 45824
rect 5810 45812 5816 45824
rect 5771 45784 5816 45812
rect 5810 45772 5816 45784
rect 5868 45772 5874 45824
rect 7742 45812 7748 45824
rect 7703 45784 7748 45812
rect 7742 45772 7748 45784
rect 7800 45772 7806 45824
rect 9858 45772 9864 45824
rect 9916 45812 9922 45824
rect 10321 45815 10379 45821
rect 10321 45812 10333 45815
rect 9916 45784 10333 45812
rect 9916 45772 9922 45784
rect 10321 45781 10333 45784
rect 10367 45781 10379 45815
rect 10321 45775 10379 45781
rect 14274 45772 14280 45824
rect 14332 45812 14338 45824
rect 14384 45812 14412 45843
rect 16574 45840 16580 45892
rect 16632 45880 16638 45892
rect 17046 45883 17104 45889
rect 17046 45880 17058 45883
rect 16632 45852 17058 45880
rect 16632 45840 16638 45852
rect 17046 45849 17058 45852
rect 17092 45849 17104 45883
rect 17046 45843 17104 45849
rect 19426 45840 19432 45892
rect 19484 45880 19490 45892
rect 19705 45883 19763 45889
rect 19705 45880 19717 45883
rect 19484 45852 19717 45880
rect 19484 45840 19490 45852
rect 19705 45849 19717 45852
rect 19751 45849 19763 45883
rect 19705 45843 19763 45849
rect 22640 45883 22698 45889
rect 22640 45849 22652 45883
rect 22686 45880 22698 45883
rect 22738 45880 22744 45892
rect 22686 45852 22744 45880
rect 22686 45849 22698 45852
rect 22640 45843 22698 45849
rect 22738 45840 22744 45852
rect 22796 45840 22802 45892
rect 25130 45889 25136 45892
rect 25124 45843 25136 45889
rect 25188 45880 25194 45892
rect 25188 45852 25224 45880
rect 25130 45840 25136 45843
rect 25188 45840 25194 45852
rect 26418 45840 26424 45892
rect 26476 45880 26482 45892
rect 28552 45880 28580 45911
rect 29730 45908 29736 45920
rect 29788 45948 29794 45960
rect 30377 45951 30435 45957
rect 30377 45948 30389 45951
rect 29788 45920 30389 45948
rect 29788 45908 29794 45920
rect 30377 45917 30389 45920
rect 30423 45917 30435 45951
rect 30377 45911 30435 45917
rect 26476 45852 28580 45880
rect 30392 45880 30420 45911
rect 30466 45908 30472 45960
rect 30524 45948 30530 45960
rect 31021 45951 31079 45957
rect 31021 45948 31033 45951
rect 30524 45920 31033 45948
rect 30524 45908 30530 45920
rect 31021 45917 31033 45920
rect 31067 45917 31079 45951
rect 31021 45911 31079 45917
rect 31386 45880 31392 45892
rect 30392 45852 31392 45880
rect 26476 45840 26482 45852
rect 31386 45840 31392 45852
rect 31444 45840 31450 45892
rect 14332 45784 14412 45812
rect 14332 45772 14338 45784
rect 14734 45772 14740 45824
rect 14792 45812 14798 45824
rect 15102 45812 15108 45824
rect 14792 45784 15108 45812
rect 14792 45772 14798 45784
rect 15102 45772 15108 45784
rect 15160 45812 15166 45824
rect 15473 45815 15531 45821
rect 15473 45812 15485 45815
rect 15160 45784 15485 45812
rect 15160 45772 15166 45784
rect 15473 45781 15485 45784
rect 15519 45781 15531 45815
rect 15930 45812 15936 45824
rect 15891 45784 15936 45812
rect 15473 45775 15531 45781
rect 15930 45772 15936 45784
rect 15988 45772 15994 45824
rect 23750 45812 23756 45824
rect 23711 45784 23756 45812
rect 23750 45772 23756 45784
rect 23808 45772 23814 45824
rect 26234 45812 26240 45824
rect 26195 45784 26240 45812
rect 26234 45772 26240 45784
rect 26292 45772 26298 45824
rect 28445 45815 28503 45821
rect 28445 45781 28457 45815
rect 28491 45812 28503 45815
rect 29730 45812 29736 45824
rect 28491 45784 29736 45812
rect 28491 45781 28503 45784
rect 28445 45775 28503 45781
rect 29730 45772 29736 45784
rect 29788 45772 29794 45824
rect 31726 45812 31754 45988
rect 31849 45951 31907 45957
rect 31849 45917 31861 45951
rect 31895 45948 31907 45951
rect 33226 45948 33232 45960
rect 31895 45920 33232 45948
rect 31895 45917 31907 45920
rect 31849 45911 31907 45917
rect 33226 45908 33232 45920
rect 33284 45908 33290 45960
rect 33318 45908 33324 45960
rect 33376 45948 33382 45960
rect 33781 45951 33839 45957
rect 33781 45948 33793 45951
rect 33376 45920 33793 45948
rect 33376 45908 33382 45920
rect 33781 45917 33793 45920
rect 33827 45948 33839 45951
rect 34330 45948 34336 45960
rect 33827 45920 34336 45948
rect 33827 45917 33839 45920
rect 33781 45911 33839 45917
rect 34330 45908 34336 45920
rect 34388 45948 34394 45960
rect 35345 45951 35403 45957
rect 35345 45948 35357 45951
rect 34388 45920 35357 45948
rect 34388 45908 34394 45920
rect 35345 45917 35357 45920
rect 35391 45948 35403 45951
rect 35820 45948 35848 46124
rect 39114 46112 39120 46124
rect 39172 46112 39178 46164
rect 39301 46155 39359 46161
rect 39301 46121 39313 46155
rect 39347 46152 39359 46155
rect 39850 46152 39856 46164
rect 39347 46124 39856 46152
rect 39347 46121 39359 46124
rect 39301 46115 39359 46121
rect 39850 46112 39856 46124
rect 39908 46112 39914 46164
rect 40957 46155 41015 46161
rect 40957 46121 40969 46155
rect 41003 46152 41015 46155
rect 41322 46152 41328 46164
rect 41003 46124 41328 46152
rect 41003 46121 41015 46124
rect 40957 46115 41015 46121
rect 41322 46112 41328 46124
rect 41380 46112 41386 46164
rect 41874 46152 41880 46164
rect 41835 46124 41880 46152
rect 41874 46112 41880 46124
rect 41932 46112 41938 46164
rect 43073 46155 43131 46161
rect 43073 46121 43085 46155
rect 43119 46152 43131 46155
rect 43162 46152 43168 46164
rect 43119 46124 43168 46152
rect 43119 46121 43131 46124
rect 43073 46115 43131 46121
rect 43162 46112 43168 46124
rect 43220 46112 43226 46164
rect 44174 46112 44180 46164
rect 44232 46152 44238 46164
rect 44269 46155 44327 46161
rect 44269 46152 44281 46155
rect 44232 46124 44281 46152
rect 44232 46112 44238 46124
rect 44269 46121 44281 46124
rect 44315 46121 44327 46155
rect 44269 46115 44327 46121
rect 45554 46112 45560 46164
rect 45612 46152 45618 46164
rect 45833 46155 45891 46161
rect 45833 46152 45845 46155
rect 45612 46124 45845 46152
rect 45612 46112 45618 46124
rect 45833 46121 45845 46124
rect 45879 46121 45891 46155
rect 45833 46115 45891 46121
rect 46474 46112 46480 46164
rect 46532 46152 46538 46164
rect 46569 46155 46627 46161
rect 46569 46152 46581 46155
rect 46532 46124 46581 46152
rect 46532 46112 46538 46124
rect 46569 46121 46581 46124
rect 46615 46121 46627 46155
rect 47302 46152 47308 46164
rect 47263 46124 47308 46152
rect 46569 46115 46627 46121
rect 47302 46112 47308 46124
rect 47360 46112 47366 46164
rect 39942 46084 39948 46096
rect 37016 46056 39948 46084
rect 35986 45948 35992 45960
rect 35391 45920 35848 45948
rect 35947 45920 35992 45948
rect 35391 45917 35403 45920
rect 35345 45911 35403 45917
rect 35986 45908 35992 45920
rect 36044 45908 36050 45960
rect 37016 45948 37044 46056
rect 39942 46044 39948 46056
rect 40000 46044 40006 46096
rect 40037 46087 40095 46093
rect 40037 46053 40049 46087
rect 40083 46053 40095 46087
rect 40037 46047 40095 46053
rect 40052 46016 40080 46047
rect 40126 46044 40132 46096
rect 40184 46084 40190 46096
rect 45094 46084 45100 46096
rect 40184 46056 45100 46084
rect 40184 46044 40190 46056
rect 45094 46044 45100 46056
rect 45152 46044 45158 46096
rect 45189 46087 45247 46093
rect 45189 46053 45201 46087
rect 45235 46084 45247 46087
rect 46750 46084 46756 46096
rect 45235 46056 46756 46084
rect 45235 46053 45247 46056
rect 45189 46047 45247 46053
rect 46750 46044 46756 46056
rect 46808 46044 46814 46096
rect 40052 45988 46428 46016
rect 36096 45920 37044 45948
rect 37921 45951 37979 45957
rect 31938 45840 31944 45892
rect 31996 45880 32002 45892
rect 32094 45883 32152 45889
rect 32094 45880 32106 45883
rect 31996 45852 32106 45880
rect 31996 45840 32002 45852
rect 32094 45849 32106 45852
rect 32140 45849 32152 45883
rect 36096 45880 36124 45920
rect 37921 45917 37933 45951
rect 37967 45948 37979 45951
rect 38473 45951 38531 45957
rect 38473 45948 38485 45951
rect 37967 45920 38485 45948
rect 37967 45917 37979 45920
rect 37921 45911 37979 45917
rect 38473 45917 38485 45920
rect 38519 45948 38531 45951
rect 39114 45948 39120 45960
rect 38519 45920 39120 45948
rect 38519 45917 38531 45920
rect 38473 45911 38531 45917
rect 39114 45908 39120 45920
rect 39172 45908 39178 45960
rect 39666 45908 39672 45960
rect 39724 45948 39730 45960
rect 39853 45951 39911 45957
rect 39853 45948 39865 45951
rect 39724 45920 39865 45948
rect 39724 45908 39730 45920
rect 39853 45917 39865 45920
rect 39899 45917 39911 45951
rect 39853 45911 39911 45917
rect 40773 45951 40831 45957
rect 40773 45917 40785 45951
rect 40819 45948 40831 45951
rect 41506 45948 41512 45960
rect 40819 45920 41512 45948
rect 40819 45917 40831 45920
rect 40773 45911 40831 45917
rect 41506 45908 41512 45920
rect 41564 45908 41570 45960
rect 41690 45908 41696 45960
rect 41748 45948 41754 45960
rect 42429 45951 42487 45957
rect 42429 45948 42441 45951
rect 41748 45920 42441 45948
rect 41748 45908 41754 45920
rect 42429 45917 42441 45920
rect 42475 45948 42487 45951
rect 42889 45951 42947 45957
rect 42889 45948 42901 45951
rect 42475 45920 42901 45948
rect 42475 45917 42487 45920
rect 42429 45911 42487 45917
rect 42889 45917 42901 45920
rect 42935 45948 42947 45951
rect 43625 45951 43683 45957
rect 43625 45948 43637 45951
rect 42935 45920 43637 45948
rect 42935 45917 42947 45920
rect 42889 45911 42947 45917
rect 43625 45917 43637 45920
rect 43671 45948 43683 45951
rect 43898 45948 43904 45960
rect 43671 45920 43904 45948
rect 43671 45917 43683 45920
rect 43625 45911 43683 45917
rect 43898 45908 43904 45920
rect 43956 45948 43962 45960
rect 46400 45957 46428 45988
rect 44085 45951 44143 45957
rect 44085 45948 44097 45951
rect 43956 45920 44097 45948
rect 43956 45908 43962 45920
rect 44085 45917 44097 45920
rect 44131 45948 44143 45951
rect 45649 45951 45707 45957
rect 45649 45948 45661 45951
rect 44131 45920 45661 45948
rect 44131 45917 44143 45920
rect 44085 45911 44143 45917
rect 45649 45917 45661 45920
rect 45695 45917 45707 45951
rect 45649 45911 45707 45917
rect 46385 45951 46443 45957
rect 46385 45917 46397 45951
rect 46431 45917 46443 45951
rect 46385 45911 46443 45917
rect 46474 45908 46480 45960
rect 46532 45948 46538 45960
rect 47121 45951 47179 45957
rect 47121 45948 47133 45951
rect 46532 45920 47133 45948
rect 46532 45908 46538 45920
rect 47121 45917 47133 45920
rect 47167 45917 47179 45951
rect 47854 45948 47860 45960
rect 47815 45920 47860 45948
rect 47121 45911 47179 45917
rect 47854 45908 47860 45920
rect 47912 45908 47918 45960
rect 32094 45843 32152 45849
rect 33060 45852 36124 45880
rect 36256 45883 36314 45889
rect 33060 45812 33088 45852
rect 36256 45849 36268 45883
rect 36302 45880 36314 45883
rect 36446 45880 36452 45892
rect 36302 45852 36452 45880
rect 36302 45849 36314 45852
rect 36256 45843 36314 45849
rect 36446 45840 36452 45852
rect 36504 45840 36510 45892
rect 44726 45880 44732 45892
rect 36556 45852 44732 45880
rect 31726 45784 33088 45812
rect 33134 45772 33140 45824
rect 33192 45812 33198 45824
rect 33229 45815 33287 45821
rect 33229 45812 33241 45815
rect 33192 45784 33241 45812
rect 33192 45772 33198 45784
rect 33229 45781 33241 45784
rect 33275 45781 33287 45815
rect 34790 45812 34796 45824
rect 34751 45784 34796 45812
rect 33229 45775 33287 45781
rect 34790 45772 34796 45784
rect 34848 45772 34854 45824
rect 35434 45772 35440 45824
rect 35492 45812 35498 45824
rect 36556 45812 36584 45852
rect 44726 45840 44732 45852
rect 44784 45880 44790 45892
rect 45278 45880 45284 45892
rect 44784 45852 45284 45880
rect 44784 45840 44790 45852
rect 45278 45840 45284 45852
rect 45336 45840 45342 45892
rect 37366 45812 37372 45824
rect 35492 45784 36584 45812
rect 37327 45784 37372 45812
rect 35492 45772 35498 45784
rect 37366 45772 37372 45784
rect 37424 45772 37430 45824
rect 48038 45812 48044 45824
rect 47999 45784 48044 45812
rect 48038 45772 48044 45784
rect 48096 45772 48102 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 5258 45608 5264 45620
rect 5219 45580 5264 45608
rect 5258 45568 5264 45580
rect 5316 45568 5322 45620
rect 6454 45608 6460 45620
rect 6415 45580 6460 45608
rect 6454 45568 6460 45580
rect 6512 45568 6518 45620
rect 9306 45608 9312 45620
rect 6564 45580 7880 45608
rect 9267 45580 9312 45608
rect 2774 45540 2780 45552
rect 1780 45512 2780 45540
rect 1780 45481 1808 45512
rect 2774 45500 2780 45512
rect 2832 45500 2838 45552
rect 1765 45475 1823 45481
rect 1765 45441 1777 45475
rect 1811 45441 1823 45475
rect 1765 45435 1823 45441
rect 2498 45432 2504 45484
rect 2556 45472 2562 45484
rect 3522 45475 3580 45481
rect 3522 45472 3534 45475
rect 2556 45444 3534 45472
rect 2556 45432 2562 45444
rect 3522 45441 3534 45444
rect 3568 45441 3580 45475
rect 4522 45472 4528 45484
rect 4483 45444 4528 45472
rect 3522 45435 3580 45441
rect 4522 45432 4528 45444
rect 4580 45432 4586 45484
rect 4706 45472 4712 45484
rect 4667 45444 4712 45472
rect 4706 45432 4712 45444
rect 4764 45432 4770 45484
rect 5077 45475 5135 45481
rect 5077 45441 5089 45475
rect 5123 45472 5135 45475
rect 5810 45472 5816 45484
rect 5123 45444 5816 45472
rect 5123 45441 5135 45444
rect 5077 45435 5135 45441
rect 5810 45432 5816 45444
rect 5868 45432 5874 45484
rect 6564 45472 6592 45580
rect 7742 45540 7748 45552
rect 6656 45512 7748 45540
rect 6656 45481 6684 45512
rect 7742 45500 7748 45512
rect 7800 45500 7806 45552
rect 7852 45540 7880 45580
rect 9306 45568 9312 45580
rect 9364 45568 9370 45620
rect 11514 45608 11520 45620
rect 11475 45580 11520 45608
rect 11514 45568 11520 45580
rect 11572 45568 11578 45620
rect 14274 45608 14280 45620
rect 14235 45580 14280 45608
rect 14274 45568 14280 45580
rect 14332 45568 14338 45620
rect 22738 45608 22744 45620
rect 22699 45580 22744 45608
rect 22738 45568 22744 45580
rect 22796 45568 22802 45620
rect 25041 45611 25099 45617
rect 25041 45577 25053 45611
rect 25087 45608 25099 45611
rect 25130 45608 25136 45620
rect 25087 45580 25136 45608
rect 25087 45577 25099 45580
rect 25041 45571 25099 45577
rect 25130 45568 25136 45580
rect 25188 45568 25194 45620
rect 28442 45568 28448 45620
rect 28500 45608 28506 45620
rect 29549 45611 29607 45617
rect 29549 45608 29561 45611
rect 28500 45580 29561 45608
rect 28500 45568 28506 45580
rect 29549 45577 29561 45580
rect 29595 45608 29607 45611
rect 30466 45608 30472 45620
rect 29595 45580 30472 45608
rect 29595 45577 29607 45580
rect 29549 45571 29607 45577
rect 30466 45568 30472 45580
rect 30524 45568 30530 45620
rect 31386 45568 31392 45620
rect 31444 45608 31450 45620
rect 31444 45580 32076 45608
rect 31444 45568 31450 45580
rect 8386 45540 8392 45552
rect 7852 45512 8392 45540
rect 6380 45444 6592 45472
rect 6641 45475 6699 45481
rect 3789 45407 3847 45413
rect 3789 45373 3801 45407
rect 3835 45404 3847 45407
rect 4614 45404 4620 45416
rect 3835 45376 4620 45404
rect 3835 45373 3847 45376
rect 3789 45367 3847 45373
rect 4614 45364 4620 45376
rect 4672 45364 4678 45416
rect 4798 45404 4804 45416
rect 4759 45376 4804 45404
rect 4798 45364 4804 45376
rect 4856 45364 4862 45416
rect 4893 45407 4951 45413
rect 4893 45373 4905 45407
rect 4939 45373 4951 45407
rect 4893 45367 4951 45373
rect 1946 45336 1952 45348
rect 1907 45308 1952 45336
rect 1946 45296 1952 45308
rect 2004 45296 2010 45348
rect 4154 45296 4160 45348
rect 4212 45296 4218 45348
rect 4908 45336 4936 45367
rect 4982 45364 4988 45416
rect 5040 45404 5046 45416
rect 5721 45407 5779 45413
rect 5721 45404 5733 45407
rect 5040 45376 5733 45404
rect 5040 45364 5046 45376
rect 5721 45373 5733 45376
rect 5767 45404 5779 45407
rect 6380 45404 6408 45444
rect 6641 45441 6653 45475
rect 6687 45441 6699 45475
rect 7009 45475 7067 45481
rect 7009 45472 7021 45475
rect 6641 45435 6699 45441
rect 6748 45444 7021 45472
rect 5767 45376 6408 45404
rect 5767 45373 5779 45376
rect 5721 45367 5779 45373
rect 6454 45364 6460 45416
rect 6512 45404 6518 45416
rect 6748 45404 6776 45444
rect 7009 45441 7021 45444
rect 7055 45441 7067 45475
rect 7009 45435 7067 45441
rect 7190 45432 7196 45484
rect 7248 45472 7254 45484
rect 7852 45481 7880 45512
rect 8386 45500 8392 45512
rect 8444 45500 8450 45552
rect 10042 45540 10048 45552
rect 8588 45512 10048 45540
rect 8588 45481 8616 45512
rect 10042 45500 10048 45512
rect 10100 45500 10106 45552
rect 12802 45540 12808 45552
rect 11716 45512 12808 45540
rect 7837 45475 7895 45481
rect 7248 45444 7341 45472
rect 7248 45432 7254 45444
rect 7837 45441 7849 45475
rect 7883 45441 7895 45475
rect 8573 45475 8631 45481
rect 8573 45472 8585 45475
rect 7837 45435 7895 45441
rect 7944 45444 8585 45472
rect 6512 45376 6776 45404
rect 6825 45407 6883 45413
rect 6512 45364 6518 45376
rect 6825 45373 6837 45407
rect 6871 45373 6883 45407
rect 6825 45367 6883 45373
rect 6917 45407 6975 45413
rect 6917 45373 6929 45407
rect 6963 45404 6975 45407
rect 7208 45404 7236 45432
rect 7944 45404 7972 45444
rect 8573 45441 8585 45444
rect 8619 45441 8631 45475
rect 8757 45475 8815 45481
rect 8757 45472 8769 45475
rect 8573 45435 8631 45441
rect 8680 45444 8769 45472
rect 6963 45376 7052 45404
rect 7208 45376 7972 45404
rect 6963 45373 6975 45376
rect 6917 45367 6975 45373
rect 6730 45336 6736 45348
rect 4908 45308 6736 45336
rect 6730 45296 6736 45308
rect 6788 45336 6794 45348
rect 6840 45336 6868 45367
rect 7024 45348 7052 45376
rect 8294 45364 8300 45416
rect 8352 45404 8358 45416
rect 8680 45404 8708 45444
rect 8757 45441 8769 45444
rect 8803 45441 8815 45475
rect 8757 45435 8815 45441
rect 8846 45432 8852 45484
rect 8904 45472 8910 45484
rect 9125 45475 9183 45481
rect 8904 45444 8949 45472
rect 8904 45432 8910 45444
rect 9125 45441 9137 45475
rect 9171 45472 9183 45475
rect 9858 45472 9864 45484
rect 9171 45444 9864 45472
rect 9171 45441 9183 45444
rect 9125 45435 9183 45441
rect 9858 45432 9864 45444
rect 9916 45432 9922 45484
rect 9953 45475 10011 45481
rect 9953 45441 9965 45475
rect 9999 45472 10011 45475
rect 10410 45472 10416 45484
rect 9999 45444 10416 45472
rect 9999 45441 10011 45444
rect 9953 45435 10011 45441
rect 8352 45376 8708 45404
rect 8941 45407 8999 45413
rect 8352 45364 8358 45376
rect 8941 45373 8953 45407
rect 8987 45373 8999 45407
rect 8941 45367 8999 45373
rect 6788 45308 6868 45336
rect 6788 45296 6794 45308
rect 2409 45271 2467 45277
rect 2409 45237 2421 45271
rect 2455 45268 2467 45271
rect 2682 45268 2688 45280
rect 2455 45240 2688 45268
rect 2455 45237 2467 45240
rect 2409 45231 2467 45237
rect 2682 45228 2688 45240
rect 2740 45268 2746 45280
rect 4172 45268 4200 45296
rect 2740 45240 4200 45268
rect 6840 45268 6868 45308
rect 7006 45296 7012 45348
rect 7064 45296 7070 45348
rect 8018 45336 8024 45348
rect 7979 45308 8024 45336
rect 8018 45296 8024 45308
rect 8076 45296 8082 45348
rect 8956 45336 8984 45367
rect 9398 45364 9404 45416
rect 9456 45404 9462 45416
rect 9968 45404 9996 45435
rect 10410 45432 10416 45444
rect 10468 45432 10474 45484
rect 11716 45481 11744 45512
rect 12802 45500 12808 45512
rect 12860 45500 12866 45552
rect 15565 45543 15623 45549
rect 13556 45512 14872 45540
rect 11701 45475 11759 45481
rect 11701 45441 11713 45475
rect 11747 45441 11759 45475
rect 12069 45475 12127 45481
rect 12069 45472 12081 45475
rect 11701 45435 11759 45441
rect 11808 45444 12081 45472
rect 9456 45376 9996 45404
rect 9456 45364 9462 45376
rect 11238 45364 11244 45416
rect 11296 45404 11302 45416
rect 11808 45404 11836 45444
rect 12069 45441 12081 45444
rect 12115 45441 12127 45475
rect 12069 45435 12127 45441
rect 12253 45475 12311 45481
rect 12253 45441 12265 45475
rect 12299 45472 12311 45475
rect 12894 45472 12900 45484
rect 12299 45444 12333 45472
rect 12855 45444 12900 45472
rect 12299 45441 12311 45444
rect 12253 45435 12311 45441
rect 11296 45376 11836 45404
rect 11885 45407 11943 45413
rect 11296 45364 11302 45376
rect 11885 45373 11897 45407
rect 11931 45373 11943 45407
rect 11885 45367 11943 45373
rect 9766 45336 9772 45348
rect 8864 45308 8984 45336
rect 9727 45308 9772 45336
rect 8864 45268 8892 45308
rect 9766 45296 9772 45308
rect 9824 45296 9830 45348
rect 10594 45336 10600 45348
rect 10555 45308 10600 45336
rect 10594 45296 10600 45308
rect 10652 45296 10658 45348
rect 11900 45336 11928 45367
rect 11974 45364 11980 45416
rect 12032 45404 12038 45416
rect 12032 45376 12077 45404
rect 12032 45364 12038 45376
rect 12158 45364 12164 45416
rect 12216 45404 12222 45416
rect 12268 45404 12296 45435
rect 12894 45432 12900 45444
rect 12952 45432 12958 45484
rect 13556 45481 13584 45512
rect 13541 45475 13599 45481
rect 13541 45441 13553 45475
rect 13587 45441 13599 45475
rect 13722 45472 13728 45484
rect 13683 45444 13728 45472
rect 13541 45435 13599 45441
rect 13556 45404 13584 45435
rect 13722 45432 13728 45444
rect 13780 45432 13786 45484
rect 14093 45475 14151 45481
rect 14093 45441 14105 45475
rect 14139 45472 14151 45475
rect 14734 45472 14740 45484
rect 14139 45444 14740 45472
rect 14139 45441 14151 45444
rect 14093 45435 14151 45441
rect 14734 45432 14740 45444
rect 14792 45432 14798 45484
rect 14844 45481 14872 45512
rect 15565 45509 15577 45543
rect 15611 45540 15623 45543
rect 16574 45540 16580 45552
rect 15611 45512 16580 45540
rect 15611 45509 15623 45512
rect 15565 45503 15623 45509
rect 16574 45500 16580 45512
rect 16632 45500 16638 45552
rect 17497 45543 17555 45549
rect 17497 45509 17509 45543
rect 17543 45540 17555 45543
rect 23750 45540 23756 45552
rect 17543 45512 22094 45540
rect 17543 45509 17555 45512
rect 17497 45503 17555 45509
rect 14829 45475 14887 45481
rect 14829 45441 14841 45475
rect 14875 45441 14887 45475
rect 15010 45472 15016 45484
rect 14971 45444 15016 45472
rect 14829 45435 14887 45441
rect 15010 45432 15016 45444
rect 15068 45472 15074 45484
rect 15381 45475 15439 45481
rect 15068 45444 15332 45472
rect 15068 45432 15074 45444
rect 12216 45376 13584 45404
rect 13817 45407 13875 45413
rect 12216 45364 12222 45376
rect 13817 45373 13829 45407
rect 13863 45373 13875 45407
rect 13817 45367 13875 45373
rect 13909 45407 13967 45413
rect 13909 45373 13921 45407
rect 13955 45373 13967 45407
rect 15102 45404 15108 45416
rect 15063 45376 15108 45404
rect 13909 45367 13967 45373
rect 12434 45336 12440 45348
rect 11900 45308 12440 45336
rect 12434 45296 12440 45308
rect 12492 45296 12498 45348
rect 13078 45336 13084 45348
rect 13039 45308 13084 45336
rect 13078 45296 13084 45308
rect 13136 45296 13142 45348
rect 6840 45240 8892 45268
rect 2740 45228 2746 45240
rect 11974 45228 11980 45280
rect 12032 45268 12038 45280
rect 12894 45268 12900 45280
rect 12032 45240 12900 45268
rect 12032 45228 12038 45240
rect 12894 45228 12900 45240
rect 12952 45268 12958 45280
rect 13832 45268 13860 45367
rect 13924 45336 13952 45367
rect 15102 45364 15108 45376
rect 15160 45364 15166 45416
rect 15197 45407 15255 45413
rect 15197 45373 15209 45407
rect 15243 45373 15255 45407
rect 15197 45367 15255 45373
rect 14458 45336 14464 45348
rect 13924 45308 14464 45336
rect 14458 45296 14464 45308
rect 14516 45336 14522 45348
rect 15212 45336 15240 45367
rect 14516 45308 15240 45336
rect 15304 45336 15332 45444
rect 15381 45441 15393 45475
rect 15427 45472 15439 45475
rect 15930 45472 15936 45484
rect 15427 45444 15936 45472
rect 15427 45441 15439 45444
rect 15381 45435 15439 45441
rect 15930 45432 15936 45444
rect 15988 45432 15994 45484
rect 18598 45481 18604 45484
rect 17313 45475 17371 45481
rect 17313 45441 17325 45475
rect 17359 45441 17371 45475
rect 17313 45435 17371 45441
rect 18592 45435 18604 45481
rect 18656 45472 18662 45484
rect 18656 45444 18692 45472
rect 16669 45339 16727 45345
rect 16669 45336 16681 45339
rect 15304 45308 16681 45336
rect 14516 45296 14522 45308
rect 16669 45305 16681 45308
rect 16715 45336 16727 45339
rect 17328 45336 17356 45435
rect 18598 45432 18604 45435
rect 18656 45432 18662 45444
rect 17402 45364 17408 45416
rect 17460 45404 17466 45416
rect 18322 45404 18328 45416
rect 17460 45376 18328 45404
rect 17460 45364 17466 45376
rect 18322 45364 18328 45376
rect 18380 45364 18386 45416
rect 19426 45336 19432 45348
rect 16715 45308 17356 45336
rect 19260 45308 19432 45336
rect 16715 45305 16727 45308
rect 16669 45299 16727 45305
rect 12952 45240 13860 45268
rect 16117 45271 16175 45277
rect 12952 45228 12958 45240
rect 16117 45237 16129 45271
rect 16163 45268 16175 45271
rect 16206 45268 16212 45280
rect 16163 45240 16212 45268
rect 16163 45237 16175 45240
rect 16117 45231 16175 45237
rect 16206 45228 16212 45240
rect 16264 45228 16270 45280
rect 17862 45228 17868 45280
rect 17920 45268 17926 45280
rect 19260 45268 19288 45308
rect 19426 45296 19432 45308
rect 19484 45336 19490 45348
rect 20165 45339 20223 45345
rect 20165 45336 20177 45339
rect 19484 45308 20177 45336
rect 19484 45296 19490 45308
rect 20165 45305 20177 45308
rect 20211 45305 20223 45339
rect 20165 45299 20223 45305
rect 20714 45296 20720 45348
rect 20772 45336 20778 45348
rect 20809 45339 20867 45345
rect 20809 45336 20821 45339
rect 20772 45308 20821 45336
rect 20772 45296 20778 45308
rect 20809 45305 20821 45308
rect 20855 45336 20867 45339
rect 21542 45336 21548 45348
rect 20855 45308 21548 45336
rect 20855 45305 20867 45308
rect 20809 45299 20867 45305
rect 21542 45296 21548 45308
rect 21600 45296 21606 45348
rect 19702 45268 19708 45280
rect 17920 45240 19288 45268
rect 19663 45240 19708 45268
rect 17920 45228 17926 45240
rect 19702 45228 19708 45240
rect 19760 45268 19766 45280
rect 19978 45268 19984 45280
rect 19760 45240 19984 45268
rect 19760 45228 19766 45240
rect 19978 45228 19984 45240
rect 20036 45228 20042 45280
rect 22066 45268 22094 45512
rect 22940 45512 23756 45540
rect 22940 45481 22968 45512
rect 23750 45500 23756 45512
rect 23808 45500 23814 45552
rect 23934 45500 23940 45552
rect 23992 45540 23998 45552
rect 26234 45540 26240 45552
rect 23992 45512 24532 45540
rect 23992 45500 23998 45512
rect 22925 45475 22983 45481
rect 22925 45441 22937 45475
rect 22971 45441 22983 45475
rect 22925 45435 22983 45441
rect 23014 45432 23020 45484
rect 23072 45472 23078 45484
rect 23293 45475 23351 45481
rect 23293 45472 23305 45475
rect 23072 45444 23305 45472
rect 23072 45432 23078 45444
rect 23293 45441 23305 45444
rect 23339 45441 23351 45475
rect 23293 45435 23351 45441
rect 23477 45475 23535 45481
rect 23477 45441 23489 45475
rect 23523 45472 23535 45475
rect 23842 45472 23848 45484
rect 23523 45444 23848 45472
rect 23523 45441 23535 45444
rect 23477 45435 23535 45441
rect 23842 45432 23848 45444
rect 23900 45472 23906 45484
rect 24504 45481 24532 45512
rect 24872 45512 26240 45540
rect 24872 45481 24900 45512
rect 26234 45500 26240 45512
rect 26292 45500 26298 45552
rect 28534 45500 28540 45552
rect 28592 45540 28598 45552
rect 30193 45543 30251 45549
rect 30193 45540 30205 45543
rect 28592 45512 30205 45540
rect 28592 45500 28598 45512
rect 30193 45509 30205 45512
rect 30239 45509 30251 45543
rect 31202 45540 31208 45552
rect 30193 45503 30251 45509
rect 30852 45512 31208 45540
rect 24305 45475 24363 45481
rect 24305 45472 24317 45475
rect 23900 45444 24317 45472
rect 23900 45432 23906 45444
rect 24305 45441 24317 45444
rect 24351 45441 24363 45475
rect 24305 45435 24363 45441
rect 24489 45475 24547 45481
rect 24489 45441 24501 45475
rect 24535 45472 24547 45475
rect 24857 45475 24915 45481
rect 24535 45444 24808 45472
rect 24535 45441 24547 45444
rect 24489 45435 24547 45441
rect 22281 45407 22339 45413
rect 22281 45373 22293 45407
rect 22327 45404 22339 45407
rect 23032 45404 23060 45432
rect 22327 45376 23060 45404
rect 23109 45407 23167 45413
rect 22327 45373 22339 45376
rect 22281 45367 22339 45373
rect 23109 45373 23121 45407
rect 23155 45373 23167 45407
rect 23109 45367 23167 45373
rect 23201 45407 23259 45413
rect 23201 45373 23213 45407
rect 23247 45404 23259 45407
rect 23658 45404 23664 45416
rect 23247 45376 23664 45404
rect 23247 45373 23259 45376
rect 23201 45367 23259 45373
rect 23124 45336 23152 45367
rect 23658 45364 23664 45376
rect 23716 45404 23722 45416
rect 24581 45407 24639 45413
rect 24581 45404 24593 45407
rect 23716 45376 24593 45404
rect 23716 45364 23722 45376
rect 24581 45373 24593 45376
rect 24627 45373 24639 45407
rect 24581 45367 24639 45373
rect 24673 45407 24731 45413
rect 24673 45373 24685 45407
rect 24719 45373 24731 45407
rect 24780 45404 24808 45444
rect 24857 45441 24869 45475
rect 24903 45441 24915 45475
rect 24857 45435 24915 45441
rect 25501 45475 25559 45481
rect 25501 45441 25513 45475
rect 25547 45472 25559 45475
rect 26326 45472 26332 45484
rect 25547 45444 26332 45472
rect 25547 45441 25559 45444
rect 25501 45435 25559 45441
rect 26326 45432 26332 45444
rect 26384 45432 26390 45484
rect 28258 45432 28264 45484
rect 28316 45472 28322 45484
rect 28425 45475 28483 45481
rect 28425 45472 28437 45475
rect 28316 45444 28437 45472
rect 28316 45432 28322 45444
rect 28425 45441 28437 45444
rect 28471 45441 28483 45475
rect 28425 45435 28483 45441
rect 28994 45432 29000 45484
rect 29052 45472 29058 45484
rect 30852 45481 30880 45512
rect 31202 45500 31208 45512
rect 31260 45500 31266 45552
rect 31573 45543 31631 45549
rect 31573 45509 31585 45543
rect 31619 45540 31631 45543
rect 31938 45540 31944 45552
rect 31619 45512 31944 45540
rect 31619 45509 31631 45512
rect 31573 45503 31631 45509
rect 31938 45500 31944 45512
rect 31996 45500 32002 45552
rect 32048 45540 32076 45580
rect 32122 45568 32128 45620
rect 32180 45608 32186 45620
rect 40218 45608 40224 45620
rect 32180 45580 40224 45608
rect 32180 45568 32186 45580
rect 40218 45568 40224 45580
rect 40276 45568 40282 45620
rect 41049 45611 41107 45617
rect 41049 45577 41061 45611
rect 41095 45608 41107 45611
rect 41230 45608 41236 45620
rect 41095 45580 41236 45608
rect 41095 45577 41107 45580
rect 41049 45571 41107 45577
rect 32217 45543 32275 45549
rect 32217 45540 32229 45543
rect 32048 45512 32229 45540
rect 32217 45509 32229 45512
rect 32263 45540 32275 45543
rect 32769 45543 32827 45549
rect 32769 45540 32781 45543
rect 32263 45512 32781 45540
rect 32263 45509 32275 45512
rect 32217 45503 32275 45509
rect 32769 45509 32781 45512
rect 32815 45540 32827 45543
rect 33318 45540 33324 45552
rect 32815 45512 33324 45540
rect 32815 45509 32827 45512
rect 32769 45503 32827 45509
rect 33318 45500 33324 45512
rect 33376 45500 33382 45552
rect 35986 45540 35992 45552
rect 33428 45512 35992 45540
rect 30837 45475 30895 45481
rect 30837 45472 30849 45475
rect 29052 45444 30849 45472
rect 29052 45432 29058 45444
rect 30837 45441 30849 45444
rect 30883 45441 30895 45475
rect 30837 45435 30895 45441
rect 30926 45432 30932 45484
rect 30984 45472 30990 45484
rect 31021 45475 31079 45481
rect 31021 45472 31033 45475
rect 30984 45444 31033 45472
rect 30984 45432 30990 45444
rect 31021 45441 31033 45444
rect 31067 45441 31079 45475
rect 31021 45435 31079 45441
rect 31389 45475 31447 45481
rect 31389 45441 31401 45475
rect 31435 45472 31447 45475
rect 33134 45472 33140 45484
rect 31435 45444 33140 45472
rect 31435 45441 31447 45444
rect 31389 45435 31447 45441
rect 33134 45432 33140 45444
rect 33192 45432 33198 45484
rect 33226 45432 33232 45484
rect 33284 45472 33290 45484
rect 33428 45472 33456 45512
rect 35986 45500 35992 45512
rect 36044 45500 36050 45552
rect 36170 45500 36176 45552
rect 36228 45540 36234 45552
rect 36633 45543 36691 45549
rect 36228 45512 36308 45540
rect 36228 45500 36234 45512
rect 33502 45481 33508 45484
rect 33284 45444 33456 45472
rect 33284 45432 33290 45444
rect 33496 45435 33508 45481
rect 33560 45472 33566 45484
rect 33560 45444 33596 45472
rect 33502 45432 33508 45435
rect 33560 45432 33566 45444
rect 35710 45432 35716 45484
rect 35768 45472 35774 45484
rect 36280 45481 36308 45512
rect 36633 45509 36645 45543
rect 36679 45540 36691 45543
rect 37522 45543 37580 45549
rect 37522 45540 37534 45543
rect 36679 45512 37534 45540
rect 36679 45509 36691 45512
rect 36633 45503 36691 45509
rect 37522 45509 37534 45512
rect 37568 45509 37580 45543
rect 37522 45503 37580 45509
rect 39114 45500 39120 45552
rect 39172 45540 39178 45552
rect 39209 45543 39267 45549
rect 39209 45540 39221 45543
rect 39172 45512 39221 45540
rect 39172 45500 39178 45512
rect 39209 45509 39221 45512
rect 39255 45540 39267 45543
rect 41064 45540 41092 45571
rect 41230 45568 41236 45580
rect 41288 45608 41294 45620
rect 41690 45608 41696 45620
rect 41288 45580 41696 45608
rect 41288 45568 41294 45580
rect 41690 45568 41696 45580
rect 41748 45568 41754 45620
rect 42426 45608 42432 45620
rect 42387 45580 42432 45608
rect 42426 45568 42432 45580
rect 42484 45568 42490 45620
rect 43441 45611 43499 45617
rect 43441 45577 43453 45611
rect 43487 45608 43499 45611
rect 43530 45608 43536 45620
rect 43487 45580 43536 45608
rect 43487 45577 43499 45580
rect 43441 45571 43499 45577
rect 43530 45568 43536 45580
rect 43588 45568 43594 45620
rect 43898 45608 43904 45620
rect 43859 45580 43904 45608
rect 43898 45568 43904 45580
rect 43956 45568 43962 45620
rect 44542 45568 44548 45620
rect 44600 45608 44606 45620
rect 44637 45611 44695 45617
rect 44637 45608 44649 45611
rect 44600 45580 44649 45608
rect 44600 45568 44606 45580
rect 44637 45577 44649 45580
rect 44683 45577 44695 45611
rect 44637 45571 44695 45577
rect 48041 45611 48099 45617
rect 48041 45577 48053 45611
rect 48087 45608 48099 45611
rect 49694 45608 49700 45620
rect 48087 45580 49700 45608
rect 48087 45577 48099 45580
rect 48041 45571 48099 45577
rect 49694 45568 49700 45580
rect 49752 45568 49758 45620
rect 39255 45512 41092 45540
rect 41156 45512 47900 45540
rect 39255 45509 39267 45512
rect 39209 45503 39267 45509
rect 35897 45475 35955 45481
rect 35897 45472 35909 45475
rect 35768 45444 35909 45472
rect 35768 45432 35774 45444
rect 35897 45441 35909 45444
rect 35943 45441 35955 45475
rect 36081 45475 36139 45481
rect 36081 45472 36093 45475
rect 35897 45435 35955 45441
rect 36004 45444 36093 45472
rect 27157 45407 27215 45413
rect 27157 45404 27169 45407
rect 24780 45376 27169 45404
rect 24673 45367 24731 45373
rect 27157 45373 27169 45376
rect 27203 45404 27215 45407
rect 27430 45404 27436 45416
rect 27203 45376 27436 45404
rect 27203 45373 27215 45376
rect 27157 45367 27215 45373
rect 23750 45336 23756 45348
rect 23124 45308 23756 45336
rect 23750 45296 23756 45308
rect 23808 45336 23814 45348
rect 24688 45336 24716 45367
rect 27430 45364 27436 45376
rect 27488 45364 27494 45416
rect 27982 45364 27988 45416
rect 28040 45404 28046 45416
rect 28169 45407 28227 45413
rect 28169 45404 28181 45407
rect 28040 45376 28181 45404
rect 28040 45364 28046 45376
rect 28169 45373 28181 45376
rect 28215 45373 28227 45407
rect 28169 45367 28227 45373
rect 30377 45407 30435 45413
rect 30377 45373 30389 45407
rect 30423 45404 30435 45407
rect 30944 45404 30972 45432
rect 31110 45404 31116 45416
rect 30423 45376 30972 45404
rect 31071 45376 31116 45404
rect 30423 45373 30435 45376
rect 30377 45367 30435 45373
rect 31110 45364 31116 45376
rect 31168 45364 31174 45416
rect 31205 45407 31263 45413
rect 31205 45373 31217 45407
rect 31251 45373 31263 45407
rect 31205 45367 31263 45373
rect 25682 45336 25688 45348
rect 23808 45308 24716 45336
rect 25643 45308 25688 45336
rect 23808 45296 23814 45308
rect 25682 45296 25688 45308
rect 25740 45296 25746 45348
rect 30190 45336 30196 45348
rect 25792 45308 27108 45336
rect 30103 45308 30196 45336
rect 25792 45268 25820 45308
rect 22066 45240 25820 45268
rect 26237 45271 26295 45277
rect 26237 45237 26249 45271
rect 26283 45268 26295 45271
rect 26326 45268 26332 45280
rect 26283 45240 26332 45268
rect 26283 45237 26295 45240
rect 26237 45231 26295 45237
rect 26326 45228 26332 45240
rect 26384 45268 26390 45280
rect 26970 45268 26976 45280
rect 26384 45240 26976 45268
rect 26384 45228 26390 45240
rect 26970 45228 26976 45240
rect 27028 45228 27034 45280
rect 27080 45268 27108 45308
rect 30190 45296 30196 45308
rect 30248 45336 30254 45348
rect 31220 45336 31248 45367
rect 35342 45364 35348 45416
rect 35400 45404 35406 45416
rect 36004 45404 36032 45444
rect 36081 45441 36093 45444
rect 36127 45441 36139 45475
rect 36081 45435 36139 45441
rect 36265 45475 36323 45481
rect 36265 45441 36277 45475
rect 36311 45441 36323 45475
rect 36265 45435 36323 45441
rect 36449 45475 36507 45481
rect 36449 45441 36461 45475
rect 36495 45472 36507 45475
rect 38654 45472 38660 45484
rect 36495 45444 38660 45472
rect 36495 45441 36507 45444
rect 36449 45435 36507 45441
rect 38654 45432 38660 45444
rect 38712 45432 38718 45484
rect 36170 45404 36176 45416
rect 35400 45376 36032 45404
rect 36131 45376 36176 45404
rect 35400 45364 35406 45376
rect 36170 45364 36176 45376
rect 36228 45364 36234 45416
rect 37277 45407 37335 45413
rect 37277 45373 37289 45407
rect 37323 45373 37335 45407
rect 37277 45367 37335 45373
rect 33134 45336 33140 45348
rect 30248 45308 33140 45336
rect 30248 45296 30254 45308
rect 33134 45296 33140 45308
rect 33192 45296 33198 45348
rect 34532 45308 35480 45336
rect 34532 45268 34560 45308
rect 27080 45240 34560 45268
rect 34606 45228 34612 45280
rect 34664 45268 34670 45280
rect 35342 45268 35348 45280
rect 34664 45240 34709 45268
rect 35303 45240 35348 45268
rect 34664 45228 34670 45240
rect 35342 45228 35348 45240
rect 35400 45228 35406 45280
rect 35452 45268 35480 45308
rect 35986 45296 35992 45348
rect 36044 45336 36050 45348
rect 37292 45336 37320 45367
rect 40034 45364 40040 45416
rect 40092 45404 40098 45416
rect 41156 45404 41184 45512
rect 41506 45432 41512 45484
rect 41564 45472 41570 45484
rect 42613 45475 42671 45481
rect 42613 45472 42625 45475
rect 41564 45444 42625 45472
rect 41564 45432 41570 45444
rect 42613 45441 42625 45444
rect 42659 45472 42671 45475
rect 43257 45475 43315 45481
rect 43257 45472 43269 45475
rect 42659 45444 43269 45472
rect 42659 45441 42671 45444
rect 42613 45435 42671 45441
rect 43257 45441 43269 45444
rect 43303 45472 43315 45475
rect 44450 45472 44456 45484
rect 43303 45444 44456 45472
rect 43303 45441 43315 45444
rect 43257 45435 43315 45441
rect 44450 45432 44456 45444
rect 44508 45432 44514 45484
rect 45094 45472 45100 45484
rect 45055 45444 45100 45472
rect 45094 45432 45100 45444
rect 45152 45432 45158 45484
rect 46014 45472 46020 45484
rect 45975 45444 46020 45472
rect 46014 45432 46020 45444
rect 46072 45432 46078 45484
rect 47872 45481 47900 45512
rect 46753 45475 46811 45481
rect 46753 45441 46765 45475
rect 46799 45441 46811 45475
rect 46753 45435 46811 45441
rect 47857 45475 47915 45481
rect 47857 45441 47869 45475
rect 47903 45441 47915 45475
rect 47857 45435 47915 45441
rect 40092 45376 41184 45404
rect 40092 45364 40098 45376
rect 45646 45364 45652 45416
rect 45704 45404 45710 45416
rect 46768 45404 46796 45435
rect 45704 45376 46796 45404
rect 45704 45364 45710 45376
rect 45830 45336 45836 45348
rect 36044 45308 37320 45336
rect 38212 45308 45836 45336
rect 36044 45296 36050 45308
rect 38212 45268 38240 45308
rect 45830 45296 45836 45308
rect 45888 45296 45894 45348
rect 45922 45296 45928 45348
rect 45980 45336 45986 45348
rect 46201 45339 46259 45345
rect 46201 45336 46213 45339
rect 45980 45308 46213 45336
rect 45980 45296 45986 45308
rect 46201 45305 46213 45308
rect 46247 45305 46259 45339
rect 46201 45299 46259 45305
rect 38654 45268 38660 45280
rect 35452 45240 38240 45268
rect 38615 45240 38660 45268
rect 38654 45228 38660 45240
rect 38712 45228 38718 45280
rect 39666 45268 39672 45280
rect 39627 45240 39672 45268
rect 39666 45228 39672 45240
rect 39724 45228 39730 45280
rect 45281 45271 45339 45277
rect 45281 45237 45293 45271
rect 45327 45268 45339 45271
rect 46474 45268 46480 45280
rect 45327 45240 46480 45268
rect 45327 45237 45339 45240
rect 45281 45231 45339 45237
rect 46474 45228 46480 45240
rect 46532 45228 46538 45280
rect 46842 45228 46848 45280
rect 46900 45268 46906 45280
rect 46937 45271 46995 45277
rect 46937 45268 46949 45271
rect 46900 45240 46949 45268
rect 46900 45228 46906 45240
rect 46937 45237 46949 45240
rect 46983 45237 46995 45271
rect 46937 45231 46995 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 2498 45064 2504 45076
rect 2459 45036 2504 45064
rect 2498 45024 2504 45036
rect 2556 45024 2562 45076
rect 4614 45024 4620 45076
rect 4672 45064 4678 45076
rect 5442 45064 5448 45076
rect 4672 45036 5448 45064
rect 4672 45024 4678 45036
rect 5442 45024 5448 45036
rect 5500 45064 5506 45076
rect 5537 45067 5595 45073
rect 5537 45064 5549 45067
rect 5500 45036 5549 45064
rect 5500 45024 5506 45036
rect 5537 45033 5549 45036
rect 5583 45033 5595 45067
rect 6914 45064 6920 45076
rect 6875 45036 6920 45064
rect 5537 45027 5595 45033
rect 6914 45024 6920 45036
rect 6972 45024 6978 45076
rect 7837 45067 7895 45073
rect 7837 45033 7849 45067
rect 7883 45064 7895 45067
rect 8386 45064 8392 45076
rect 7883 45036 8392 45064
rect 7883 45033 7895 45036
rect 7837 45027 7895 45033
rect 8386 45024 8392 45036
rect 8444 45024 8450 45076
rect 14366 45064 14372 45076
rect 14327 45036 14372 45064
rect 14366 45024 14372 45036
rect 14424 45024 14430 45076
rect 15654 45064 15660 45076
rect 15615 45036 15660 45064
rect 15654 45024 15660 45036
rect 15712 45024 15718 45076
rect 18322 45024 18328 45076
rect 18380 45064 18386 45076
rect 19797 45067 19855 45073
rect 19797 45064 19809 45067
rect 18380 45036 19809 45064
rect 18380 45024 18386 45036
rect 19797 45033 19809 45036
rect 19843 45033 19855 45067
rect 20714 45064 20720 45076
rect 19797 45027 19855 45033
rect 19904 45036 20720 45064
rect 4982 44996 4988 45008
rect 4943 44968 4988 44996
rect 4982 44956 4988 44968
rect 5040 44956 5046 45008
rect 10137 44999 10195 45005
rect 10137 44965 10149 44999
rect 10183 44996 10195 44999
rect 10410 44996 10416 45008
rect 10183 44968 10416 44996
rect 10183 44965 10195 44968
rect 10137 44959 10195 44965
rect 10410 44956 10416 44968
rect 10468 44996 10474 45008
rect 10468 44968 12664 44996
rect 10468 44956 10474 44968
rect 2961 44931 3019 44937
rect 2961 44897 2973 44931
rect 3007 44928 3019 44931
rect 4798 44928 4804 44940
rect 3007 44900 4804 44928
rect 3007 44897 3019 44900
rect 2961 44891 3019 44897
rect 4798 44888 4804 44900
rect 4856 44928 4862 44940
rect 7006 44928 7012 44940
rect 4856 44900 7012 44928
rect 4856 44888 4862 44900
rect 7006 44888 7012 44900
rect 7064 44888 7070 44940
rect 12526 44928 12532 44940
rect 9646 44900 12532 44928
rect 2682 44860 2688 44872
rect 2643 44832 2688 44860
rect 2682 44820 2688 44832
rect 2740 44820 2746 44872
rect 2869 44863 2927 44869
rect 2869 44829 2881 44863
rect 2915 44829 2927 44863
rect 2869 44823 2927 44829
rect 2038 44724 2044 44736
rect 1999 44696 2044 44724
rect 2038 44684 2044 44696
rect 2096 44684 2102 44736
rect 2682 44684 2688 44736
rect 2740 44724 2746 44736
rect 2884 44724 2912 44823
rect 3050 44820 3056 44872
rect 3108 44860 3114 44872
rect 3237 44863 3295 44869
rect 3108 44832 3153 44860
rect 3108 44820 3114 44832
rect 3237 44829 3249 44863
rect 3283 44829 3295 44863
rect 3237 44823 3295 44829
rect 3252 44792 3280 44823
rect 3602 44820 3608 44872
rect 3660 44860 3666 44872
rect 9646 44860 9674 44900
rect 12526 44888 12532 44900
rect 12584 44888 12590 44940
rect 12636 44869 12664 44968
rect 13722 44956 13728 45008
rect 13780 44996 13786 45008
rect 16666 44996 16672 45008
rect 13780 44968 16672 44996
rect 13780 44956 13786 44968
rect 16666 44956 16672 44968
rect 16724 44956 16730 45008
rect 17126 44956 17132 45008
rect 17184 44996 17190 45008
rect 17184 44968 18276 44996
rect 17184 44956 17190 44968
rect 17310 44888 17316 44940
rect 17368 44928 17374 44940
rect 17862 44928 17868 44940
rect 17368 44900 17868 44928
rect 17368 44888 17374 44900
rect 17862 44888 17868 44900
rect 17920 44928 17926 44940
rect 18248 44937 18276 44968
rect 18598 44956 18604 45008
rect 18656 44996 18662 45008
rect 18693 44999 18751 45005
rect 18693 44996 18705 44999
rect 18656 44968 18705 44996
rect 18656 44956 18662 44968
rect 18693 44965 18705 44968
rect 18739 44965 18751 44999
rect 18693 44959 18751 44965
rect 18782 44956 18788 45008
rect 18840 44996 18846 45008
rect 19337 44999 19395 45005
rect 19337 44996 19349 44999
rect 18840 44968 19349 44996
rect 18840 44956 18846 44968
rect 19337 44965 19349 44968
rect 19383 44996 19395 44999
rect 19904 44996 19932 45036
rect 20714 45024 20720 45036
rect 20772 45024 20778 45076
rect 21729 45067 21787 45073
rect 21729 45033 21741 45067
rect 21775 45064 21787 45067
rect 22094 45064 22100 45076
rect 21775 45036 22100 45064
rect 21775 45033 21787 45036
rect 21729 45027 21787 45033
rect 22094 45024 22100 45036
rect 22152 45064 22158 45076
rect 22554 45064 22560 45076
rect 22152 45036 22560 45064
rect 22152 45024 22158 45036
rect 22554 45024 22560 45036
rect 22612 45024 22618 45076
rect 22925 45067 22983 45073
rect 22925 45033 22937 45067
rect 22971 45064 22983 45067
rect 23106 45064 23112 45076
rect 22971 45036 23112 45064
rect 22971 45033 22983 45036
rect 22925 45027 22983 45033
rect 23106 45024 23112 45036
rect 23164 45024 23170 45076
rect 24578 45024 24584 45076
rect 24636 45064 24642 45076
rect 25133 45067 25191 45073
rect 25133 45064 25145 45067
rect 24636 45036 25145 45064
rect 24636 45024 24642 45036
rect 25133 45033 25145 45036
rect 25179 45064 25191 45067
rect 25685 45067 25743 45073
rect 25685 45064 25697 45067
rect 25179 45036 25697 45064
rect 25179 45033 25191 45036
rect 25133 45027 25191 45033
rect 25685 45033 25697 45036
rect 25731 45064 25743 45067
rect 26970 45064 26976 45076
rect 25731 45036 26976 45064
rect 25731 45033 25743 45036
rect 25685 45027 25743 45033
rect 26970 45024 26976 45036
rect 27028 45024 27034 45076
rect 28258 45064 28264 45076
rect 28219 45036 28264 45064
rect 28258 45024 28264 45036
rect 28316 45024 28322 45076
rect 28350 45024 28356 45076
rect 28408 45064 28414 45076
rect 28810 45064 28816 45076
rect 28408 45036 28816 45064
rect 28408 45024 28414 45036
rect 28810 45024 28816 45036
rect 28868 45024 28874 45076
rect 33226 45064 33232 45076
rect 30392 45036 33232 45064
rect 19383 44968 19932 44996
rect 21376 44968 24532 44996
rect 19383 44965 19395 44968
rect 19337 44959 19395 44965
rect 18233 44931 18291 44937
rect 17920 44900 18184 44928
rect 17920 44888 17926 44900
rect 11793 44863 11851 44869
rect 11793 44860 11805 44863
rect 3660 44832 9674 44860
rect 10796 44832 11805 44860
rect 3660 44820 3666 44832
rect 4338 44792 4344 44804
rect 3252 44764 4344 44792
rect 4338 44752 4344 44764
rect 4396 44752 4402 44804
rect 4433 44795 4491 44801
rect 4433 44761 4445 44795
rect 4479 44792 4491 44795
rect 4706 44792 4712 44804
rect 4479 44764 4712 44792
rect 4479 44761 4491 44764
rect 4433 44755 4491 44761
rect 4706 44752 4712 44764
rect 4764 44792 4770 44804
rect 5258 44792 5264 44804
rect 4764 44764 5264 44792
rect 4764 44752 4770 44764
rect 5258 44752 5264 44764
rect 5316 44752 5322 44804
rect 10796 44736 10824 44832
rect 11793 44829 11805 44832
rect 11839 44829 11851 44863
rect 11793 44823 11851 44829
rect 12621 44863 12679 44869
rect 12621 44829 12633 44863
rect 12667 44860 12679 44863
rect 14182 44860 14188 44872
rect 12667 44832 14188 44860
rect 12667 44829 12679 44832
rect 12621 44823 12679 44829
rect 14182 44820 14188 44832
rect 14240 44860 14246 44872
rect 14918 44860 14924 44872
rect 14240 44832 14924 44860
rect 14240 44820 14246 44832
rect 14918 44820 14924 44832
rect 14976 44860 14982 44872
rect 15473 44863 15531 44869
rect 15473 44860 15485 44863
rect 14976 44832 15485 44860
rect 14976 44820 14982 44832
rect 15473 44829 15485 44832
rect 15519 44860 15531 44863
rect 16206 44860 16212 44872
rect 15519 44832 16212 44860
rect 15519 44829 15531 44832
rect 15473 44823 15531 44829
rect 16206 44820 16212 44832
rect 16264 44820 16270 44872
rect 17957 44863 18015 44869
rect 17957 44829 17969 44863
rect 18003 44860 18015 44863
rect 18046 44860 18052 44872
rect 18003 44832 18052 44860
rect 18003 44829 18015 44832
rect 17957 44823 18015 44829
rect 18046 44820 18052 44832
rect 18104 44820 18110 44872
rect 18156 44871 18184 44900
rect 18233 44897 18245 44931
rect 18279 44897 18291 44931
rect 18233 44891 18291 44897
rect 18141 44865 18199 44871
rect 18141 44831 18153 44865
rect 18187 44831 18199 44865
rect 18141 44825 18199 44831
rect 18322 44820 18328 44872
rect 18380 44860 18386 44872
rect 18509 44863 18567 44869
rect 18380 44832 18425 44860
rect 18380 44820 18386 44832
rect 18509 44829 18521 44863
rect 18555 44860 18567 44863
rect 19702 44860 19708 44872
rect 18555 44832 19708 44860
rect 18555 44829 18567 44832
rect 18509 44823 18567 44829
rect 19702 44820 19708 44832
rect 19760 44820 19766 44872
rect 20346 44860 20352 44872
rect 20307 44832 20352 44860
rect 20346 44820 20352 44832
rect 20404 44820 20410 44872
rect 21376 44860 21404 44968
rect 21542 44888 21548 44940
rect 21600 44928 21606 44940
rect 24504 44928 24532 44968
rect 24762 44956 24768 45008
rect 24820 44996 24826 45008
rect 30285 44999 30343 45005
rect 30285 44996 30297 44999
rect 24820 44968 30297 44996
rect 24820 44956 24826 44968
rect 30285 44965 30297 44968
rect 30331 44965 30343 44999
rect 30285 44959 30343 44965
rect 27709 44931 27767 44937
rect 27709 44928 27721 44931
rect 21600 44900 22324 44928
rect 24504 44900 27721 44928
rect 21600 44888 21606 44900
rect 22296 44869 22324 44900
rect 27709 44897 27721 44900
rect 27755 44928 27767 44931
rect 28350 44928 28356 44940
rect 27755 44900 28356 44928
rect 27755 44897 27767 44900
rect 27709 44891 27767 44897
rect 28350 44888 28356 44900
rect 28408 44888 28414 44940
rect 28534 44888 28540 44940
rect 28592 44928 28598 44940
rect 30392 44937 30420 45036
rect 33226 45024 33232 45036
rect 33284 45024 33290 45076
rect 33502 45064 33508 45076
rect 33463 45036 33508 45064
rect 33502 45024 33508 45036
rect 33560 45024 33566 45076
rect 34057 45067 34115 45073
rect 34057 45033 34069 45067
rect 34103 45064 34115 45067
rect 34330 45064 34336 45076
rect 34103 45036 34336 45064
rect 34103 45033 34115 45036
rect 34057 45027 34115 45033
rect 34330 45024 34336 45036
rect 34388 45024 34394 45076
rect 35342 45024 35348 45076
rect 35400 45064 35406 45076
rect 36446 45064 36452 45076
rect 35400 45036 36308 45064
rect 36407 45036 36452 45064
rect 35400 45024 35406 45036
rect 31754 44996 31760 45008
rect 31715 44968 31760 44996
rect 31754 44956 31760 44968
rect 31812 44956 31818 45008
rect 34790 44996 34796 45008
rect 32968 44968 34796 44996
rect 28629 44931 28687 44937
rect 28629 44928 28641 44931
rect 28592 44900 28641 44928
rect 28592 44888 28598 44900
rect 28629 44897 28641 44900
rect 28675 44897 28687 44931
rect 30377 44931 30435 44937
rect 30377 44928 30389 44931
rect 28629 44891 28687 44897
rect 29564 44900 30389 44928
rect 20456 44832 21404 44860
rect 22281 44863 22339 44869
rect 12406 44764 18368 44792
rect 3878 44724 3884 44736
rect 2740 44696 3884 44724
rect 2740 44684 2746 44696
rect 3878 44684 3884 44696
rect 3936 44684 3942 44736
rect 6365 44727 6423 44733
rect 6365 44693 6377 44727
rect 6411 44724 6423 44727
rect 6454 44724 6460 44736
rect 6411 44696 6460 44724
rect 6411 44693 6423 44696
rect 6365 44687 6423 44693
rect 6454 44684 6460 44696
rect 6512 44684 6518 44736
rect 8294 44724 8300 44736
rect 8255 44696 8300 44724
rect 8294 44684 8300 44696
rect 8352 44684 8358 44736
rect 9493 44727 9551 44733
rect 9493 44693 9505 44727
rect 9539 44724 9551 44727
rect 9674 44724 9680 44736
rect 9539 44696 9680 44724
rect 9539 44693 9551 44696
rect 9493 44687 9551 44693
rect 9674 44684 9680 44696
rect 9732 44684 9738 44736
rect 10778 44724 10784 44736
rect 10739 44696 10784 44724
rect 10778 44684 10784 44696
rect 10836 44684 10842 44736
rect 11238 44724 11244 44736
rect 11199 44696 11244 44724
rect 11238 44684 11244 44696
rect 11296 44684 11302 44736
rect 11977 44727 12035 44733
rect 11977 44693 11989 44727
rect 12023 44724 12035 44727
rect 12406 44724 12434 44764
rect 12023 44696 12434 44724
rect 13449 44727 13507 44733
rect 12023 44693 12035 44696
rect 11977 44687 12035 44693
rect 13449 44693 13461 44727
rect 13495 44724 13507 44727
rect 13722 44724 13728 44736
rect 13495 44696 13728 44724
rect 13495 44693 13507 44696
rect 13449 44687 13507 44693
rect 13722 44684 13728 44696
rect 13780 44684 13786 44736
rect 14921 44727 14979 44733
rect 14921 44693 14933 44727
rect 14967 44724 14979 44727
rect 15010 44724 15016 44736
rect 14967 44696 15016 44724
rect 14967 44693 14979 44696
rect 14921 44687 14979 44693
rect 15010 44684 15016 44696
rect 15068 44684 15074 44736
rect 16206 44724 16212 44736
rect 16167 44696 16212 44724
rect 16206 44684 16212 44696
rect 16264 44684 16270 44736
rect 17310 44684 17316 44736
rect 17368 44724 17374 44736
rect 17405 44727 17463 44733
rect 17405 44724 17417 44727
rect 17368 44696 17417 44724
rect 17368 44684 17374 44696
rect 17405 44693 17417 44696
rect 17451 44693 17463 44727
rect 18340 44724 18368 44764
rect 19426 44752 19432 44804
rect 19484 44792 19490 44804
rect 20456 44792 20484 44832
rect 22281 44829 22293 44863
rect 22327 44860 22339 44863
rect 22741 44863 22799 44869
rect 22741 44860 22753 44863
rect 22327 44832 22753 44860
rect 22327 44829 22339 44832
rect 22281 44823 22339 44829
rect 22741 44829 22753 44832
rect 22787 44860 22799 44863
rect 22787 44858 24532 44860
rect 24578 44858 24584 44872
rect 22787 44832 24584 44858
rect 22787 44829 22799 44832
rect 24504 44830 24584 44832
rect 22741 44823 22799 44829
rect 24578 44820 24584 44830
rect 24636 44860 24642 44872
rect 24636 44832 24681 44860
rect 24636 44820 24642 44832
rect 28442 44820 28448 44872
rect 28500 44860 28506 44872
rect 28721 44863 28779 44869
rect 28500 44832 28545 44860
rect 28500 44820 28506 44832
rect 28721 44829 28733 44863
rect 28767 44829 28779 44863
rect 28721 44823 28779 44829
rect 19484 44764 20484 44792
rect 20616 44795 20674 44801
rect 19484 44752 19490 44764
rect 20616 44761 20628 44795
rect 20662 44792 20674 44795
rect 20898 44792 20904 44804
rect 20662 44764 20904 44792
rect 20662 44761 20674 44764
rect 20616 44755 20674 44761
rect 20898 44752 20904 44764
rect 20956 44752 20962 44804
rect 23566 44752 23572 44804
rect 23624 44792 23630 44804
rect 27338 44792 27344 44804
rect 23624 44764 27344 44792
rect 23624 44752 23630 44764
rect 27338 44752 27344 44764
rect 27396 44752 27402 44804
rect 20990 44724 20996 44736
rect 18340 44696 20996 44724
rect 17405 44687 17463 44693
rect 20990 44684 20996 44696
rect 21048 44684 21054 44736
rect 23845 44727 23903 44733
rect 23845 44693 23857 44727
rect 23891 44724 23903 44727
rect 23934 44724 23940 44736
rect 23891 44696 23940 44724
rect 23891 44693 23903 44696
rect 23845 44687 23903 44693
rect 23934 44684 23940 44696
rect 23992 44684 23998 44736
rect 24394 44724 24400 44736
rect 24355 44696 24400 44724
rect 24394 44684 24400 44696
rect 24452 44684 24458 44736
rect 28534 44684 28540 44736
rect 28592 44724 28598 44736
rect 28736 44724 28764 44823
rect 28810 44820 28816 44872
rect 28868 44860 28874 44872
rect 28994 44860 29000 44872
rect 28868 44832 28913 44860
rect 28955 44832 29000 44860
rect 28868 44820 28874 44832
rect 28994 44820 29000 44832
rect 29052 44820 29058 44872
rect 28902 44752 28908 44804
rect 28960 44792 28966 44804
rect 29564 44792 29592 44900
rect 30377 44897 30389 44900
rect 30423 44897 30435 44931
rect 30377 44891 30435 44897
rect 32214 44888 32220 44940
rect 32272 44928 32278 44940
rect 32968 44928 32996 44968
rect 34790 44956 34796 44968
rect 34848 44956 34854 45008
rect 35894 44956 35900 45008
rect 35952 44956 35958 45008
rect 36280 44996 36308 45036
rect 36446 45024 36452 45036
rect 36504 45024 36510 45076
rect 39025 45067 39083 45073
rect 39025 45033 39037 45067
rect 39071 45064 39083 45067
rect 39114 45064 39120 45076
rect 39071 45036 39120 45064
rect 39071 45033 39083 45036
rect 39025 45027 39083 45033
rect 39114 45024 39120 45036
rect 39172 45024 39178 45076
rect 43898 45064 43904 45076
rect 43859 45036 43904 45064
rect 43898 45024 43904 45036
rect 43956 45024 43962 45076
rect 45094 45064 45100 45076
rect 45055 45036 45100 45064
rect 45094 45024 45100 45036
rect 45152 45024 45158 45076
rect 46014 45064 46020 45076
rect 45975 45036 46020 45064
rect 46014 45024 46020 45036
rect 46072 45024 46078 45076
rect 47578 45024 47584 45076
rect 47636 45064 47642 45076
rect 47857 45067 47915 45073
rect 47857 45064 47869 45067
rect 47636 45036 47869 45064
rect 47636 45024 47642 45036
rect 47857 45033 47869 45036
rect 47903 45033 47915 45067
rect 47857 45027 47915 45033
rect 39666 44996 39672 45008
rect 36280 44968 39672 44996
rect 39666 44956 39672 44968
rect 39724 44956 39730 45008
rect 33134 44928 33140 44940
rect 32272 44900 32996 44928
rect 33095 44900 33140 44928
rect 32272 44888 32278 44900
rect 30285 44863 30343 44869
rect 30285 44829 30297 44863
rect 30331 44860 30343 44863
rect 30331 44832 30788 44860
rect 30331 44829 30343 44832
rect 30285 44823 30343 44829
rect 28960 44764 29592 44792
rect 29641 44795 29699 44801
rect 28960 44752 28966 44764
rect 29641 44761 29653 44795
rect 29687 44792 29699 44795
rect 29730 44792 29736 44804
rect 29687 44764 29736 44792
rect 29687 44761 29699 44764
rect 29641 44755 29699 44761
rect 29730 44752 29736 44764
rect 29788 44752 29794 44804
rect 30466 44752 30472 44804
rect 30524 44792 30530 44804
rect 30622 44795 30680 44801
rect 30622 44792 30634 44795
rect 30524 44764 30634 44792
rect 30524 44752 30530 44764
rect 30622 44761 30634 44764
rect 30668 44761 30680 44795
rect 30760 44792 30788 44832
rect 31202 44820 31208 44872
rect 31260 44860 31266 44872
rect 32968 44869 32996 44900
rect 33134 44888 33140 44900
rect 33192 44888 33198 44940
rect 35912 44928 35940 44956
rect 35989 44931 36047 44937
rect 35989 44928 36001 44931
rect 35912 44900 36001 44928
rect 35989 44897 36001 44900
rect 36035 44928 36047 44931
rect 36170 44928 36176 44940
rect 36035 44900 36176 44928
rect 36035 44897 36047 44900
rect 35989 44891 36047 44897
rect 36170 44888 36176 44900
rect 36228 44888 36234 44940
rect 44450 44888 44456 44940
rect 44508 44928 44514 44940
rect 47302 44928 47308 44940
rect 44508 44900 47308 44928
rect 44508 44888 44514 44900
rect 32769 44863 32827 44869
rect 32769 44860 32781 44863
rect 31260 44832 32781 44860
rect 31260 44820 31266 44832
rect 32769 44829 32781 44832
rect 32815 44829 32827 44863
rect 32769 44823 32827 44829
rect 32953 44863 33011 44869
rect 32953 44829 32965 44863
rect 32999 44829 33011 44863
rect 32953 44823 33011 44829
rect 33045 44863 33103 44869
rect 33045 44829 33057 44863
rect 33091 44860 33103 44863
rect 33226 44860 33232 44872
rect 33091 44832 33232 44860
rect 33091 44829 33103 44832
rect 33045 44823 33103 44829
rect 33226 44820 33232 44832
rect 33284 44820 33290 44872
rect 33321 44863 33379 44869
rect 33321 44829 33333 44863
rect 33367 44860 33379 44863
rect 34606 44860 34612 44872
rect 33367 44832 34612 44860
rect 33367 44829 33379 44832
rect 33321 44823 33379 44829
rect 34606 44820 34612 44832
rect 34664 44820 34670 44872
rect 35710 44860 35716 44872
rect 35671 44832 35716 44860
rect 35710 44820 35716 44832
rect 35768 44820 35774 44872
rect 35802 44820 35808 44872
rect 35860 44860 35866 44872
rect 35897 44863 35955 44869
rect 35897 44860 35909 44863
rect 35860 44832 35909 44860
rect 35860 44820 35866 44832
rect 35897 44829 35909 44832
rect 35943 44829 35955 44863
rect 36078 44860 36084 44872
rect 36039 44832 36084 44860
rect 35897 44823 35955 44829
rect 36078 44820 36084 44832
rect 36136 44820 36142 44872
rect 36265 44863 36323 44869
rect 36265 44829 36277 44863
rect 36311 44860 36323 44863
rect 37366 44860 37372 44872
rect 36311 44832 37372 44860
rect 36311 44829 36323 44832
rect 36265 44823 36323 44829
rect 37366 44820 37372 44832
rect 37424 44820 37430 44872
rect 45738 44860 45744 44872
rect 41386 44832 45744 44860
rect 41386 44792 41414 44832
rect 45738 44820 45744 44832
rect 45796 44820 45802 44872
rect 45848 44869 45876 44900
rect 47302 44888 47308 44900
rect 47360 44888 47366 44940
rect 45833 44863 45891 44869
rect 45833 44829 45845 44863
rect 45879 44829 45891 44863
rect 45833 44823 45891 44829
rect 46937 44863 46995 44869
rect 46937 44829 46949 44863
rect 46983 44829 46995 44863
rect 47670 44860 47676 44872
rect 47631 44832 47676 44860
rect 46937 44823 46995 44829
rect 46952 44792 46980 44823
rect 47670 44820 47676 44832
rect 47728 44820 47734 44872
rect 30760 44764 41414 44792
rect 44376 44764 46980 44792
rect 30622 44755 30680 44761
rect 44376 44736 44404 44764
rect 31018 44724 31024 44736
rect 28592 44696 31024 44724
rect 28592 44684 28598 44696
rect 31018 44684 31024 44696
rect 31076 44684 31082 44736
rect 32214 44724 32220 44736
rect 32175 44696 32220 44724
rect 32214 44684 32220 44696
rect 32272 44684 32278 44736
rect 34698 44684 34704 44736
rect 34756 44724 34762 44736
rect 35161 44727 35219 44733
rect 35161 44724 35173 44727
rect 34756 44696 35173 44724
rect 34756 44684 34762 44696
rect 35161 44693 35173 44696
rect 35207 44724 35219 44727
rect 35802 44724 35808 44736
rect 35207 44696 35808 44724
rect 35207 44693 35219 44696
rect 35161 44687 35219 44693
rect 35802 44684 35808 44696
rect 35860 44724 35866 44736
rect 40494 44724 40500 44736
rect 35860 44696 40500 44724
rect 35860 44684 35866 44696
rect 40494 44684 40500 44696
rect 40552 44684 40558 44736
rect 44358 44724 44364 44736
rect 44319 44696 44364 44724
rect 44358 44684 44364 44696
rect 44416 44684 44422 44736
rect 46842 44684 46848 44736
rect 46900 44724 46906 44736
rect 47121 44727 47179 44733
rect 47121 44724 47133 44727
rect 46900 44696 47133 44724
rect 46900 44684 46906 44696
rect 47121 44693 47133 44696
rect 47167 44693 47179 44727
rect 47121 44687 47179 44693
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 8846 44480 8852 44532
rect 8904 44520 8910 44532
rect 9953 44523 10011 44529
rect 9953 44520 9965 44523
rect 8904 44492 9965 44520
rect 8904 44480 8910 44492
rect 9953 44489 9965 44492
rect 9999 44520 10011 44523
rect 10137 44523 10195 44529
rect 10137 44520 10149 44523
rect 9999 44492 10149 44520
rect 9999 44489 10011 44492
rect 9953 44483 10011 44489
rect 10137 44489 10149 44492
rect 10183 44489 10195 44523
rect 10137 44483 10195 44489
rect 10704 44492 12572 44520
rect 6730 44412 6736 44464
rect 6788 44452 6794 44464
rect 9033 44455 9091 44461
rect 9033 44452 9045 44455
rect 6788 44424 9045 44452
rect 6788 44412 6794 44424
rect 9033 44421 9045 44424
rect 9079 44421 9091 44455
rect 9033 44415 9091 44421
rect 9217 44455 9275 44461
rect 9217 44421 9229 44455
rect 9263 44452 9275 44455
rect 9674 44452 9680 44464
rect 9263 44424 9680 44452
rect 9263 44421 9275 44424
rect 9217 44415 9275 44421
rect 9674 44412 9680 44424
rect 9732 44452 9738 44464
rect 10704 44452 10732 44492
rect 9732 44424 10732 44452
rect 9732 44412 9738 44424
rect 10778 44412 10784 44464
rect 10836 44452 10842 44464
rect 10836 44424 12112 44452
rect 10836 44412 10842 44424
rect 7929 44387 7987 44393
rect 7929 44384 7941 44387
rect 7392 44356 7941 44384
rect 2133 44319 2191 44325
rect 2133 44285 2145 44319
rect 2179 44316 2191 44319
rect 2593 44319 2651 44325
rect 2593 44316 2605 44319
rect 2179 44288 2605 44316
rect 2179 44285 2191 44288
rect 2133 44279 2191 44285
rect 2593 44285 2605 44288
rect 2639 44316 2651 44319
rect 2774 44316 2780 44328
rect 2639 44288 2780 44316
rect 2639 44285 2651 44288
rect 2593 44279 2651 44285
rect 2774 44276 2780 44288
rect 2832 44276 2838 44328
rect 4338 44316 4344 44328
rect 4251 44288 4344 44316
rect 4338 44276 4344 44288
rect 4396 44316 4402 44328
rect 4798 44316 4804 44328
rect 4396 44288 4804 44316
rect 4396 44276 4402 44288
rect 4798 44276 4804 44288
rect 4856 44276 4862 44328
rect 3050 44208 3056 44260
rect 3108 44248 3114 44260
rect 3697 44251 3755 44257
rect 3697 44248 3709 44251
rect 3108 44220 3709 44248
rect 3108 44208 3114 44220
rect 3697 44217 3709 44220
rect 3743 44217 3755 44251
rect 3697 44211 3755 44217
rect 2774 44140 2780 44192
rect 2832 44180 2838 44192
rect 3145 44183 3203 44189
rect 3145 44180 3157 44183
rect 2832 44152 3157 44180
rect 2832 44140 2838 44152
rect 3145 44149 3157 44152
rect 3191 44149 3203 44183
rect 3145 44143 3203 44149
rect 4893 44183 4951 44189
rect 4893 44149 4905 44183
rect 4939 44180 4951 44183
rect 4982 44180 4988 44192
rect 4939 44152 4988 44180
rect 4939 44149 4951 44152
rect 4893 44143 4951 44149
rect 4982 44140 4988 44152
rect 5040 44140 5046 44192
rect 6454 44140 6460 44192
rect 6512 44180 6518 44192
rect 7392 44189 7420 44356
rect 7929 44353 7941 44356
rect 7975 44353 7987 44387
rect 10226 44384 10232 44396
rect 10187 44356 10232 44384
rect 7929 44347 7987 44353
rect 10226 44344 10232 44356
rect 10284 44344 10290 44396
rect 11698 44384 11704 44396
rect 11659 44356 11704 44384
rect 11698 44344 11704 44356
rect 11756 44344 11762 44396
rect 11974 44384 11980 44396
rect 11808 44356 11980 44384
rect 9953 44319 10011 44325
rect 9953 44285 9965 44319
rect 9999 44316 10011 44319
rect 11808 44316 11836 44356
rect 11974 44344 11980 44356
rect 12032 44344 12038 44396
rect 12084 44393 12112 44424
rect 12069 44387 12127 44393
rect 12069 44353 12081 44387
rect 12115 44353 12127 44387
rect 12069 44347 12127 44353
rect 12158 44344 12164 44396
rect 12216 44384 12222 44396
rect 12253 44387 12311 44393
rect 12253 44384 12265 44387
rect 12216 44356 12265 44384
rect 12216 44344 12222 44356
rect 12253 44353 12265 44356
rect 12299 44353 12311 44387
rect 12544 44384 12572 44492
rect 13170 44480 13176 44532
rect 13228 44520 13234 44532
rect 14458 44520 14464 44532
rect 13228 44492 14464 44520
rect 13228 44480 13234 44492
rect 14458 44480 14464 44492
rect 14516 44480 14522 44532
rect 14918 44480 14924 44532
rect 14976 44520 14982 44532
rect 15013 44523 15071 44529
rect 15013 44520 15025 44523
rect 14976 44492 15025 44520
rect 14976 44480 14982 44492
rect 15013 44489 15025 44492
rect 15059 44489 15071 44523
rect 15838 44520 15844 44532
rect 15799 44492 15844 44520
rect 15013 44483 15071 44489
rect 15838 44480 15844 44492
rect 15896 44480 15902 44532
rect 16206 44480 16212 44532
rect 16264 44520 16270 44532
rect 17957 44523 18015 44529
rect 17957 44520 17969 44523
rect 16264 44492 17969 44520
rect 16264 44480 16270 44492
rect 17957 44489 17969 44492
rect 18003 44489 18015 44523
rect 17957 44483 18015 44489
rect 18322 44480 18328 44532
rect 18380 44520 18386 44532
rect 19613 44523 19671 44529
rect 19613 44520 19625 44523
rect 18380 44492 19625 44520
rect 18380 44480 18386 44492
rect 19613 44489 19625 44492
rect 19659 44520 19671 44523
rect 20530 44520 20536 44532
rect 19659 44492 20536 44520
rect 19659 44489 19671 44492
rect 19613 44483 19671 44489
rect 20530 44480 20536 44492
rect 20588 44480 20594 44532
rect 20898 44520 20904 44532
rect 20859 44492 20904 44520
rect 20898 44480 20904 44492
rect 20956 44480 20962 44532
rect 20990 44480 20996 44532
rect 21048 44520 21054 44532
rect 45646 44520 45652 44532
rect 21048 44492 45652 44520
rect 21048 44480 21054 44492
rect 45646 44480 45652 44492
rect 45704 44480 45710 44532
rect 45830 44480 45836 44532
rect 45888 44520 45894 44532
rect 46385 44523 46443 44529
rect 46385 44520 46397 44523
rect 45888 44492 46397 44520
rect 45888 44480 45894 44492
rect 46385 44489 46397 44492
rect 46431 44520 46443 44523
rect 47854 44520 47860 44532
rect 46431 44492 47860 44520
rect 46431 44489 46443 44492
rect 46385 44483 46443 44489
rect 47854 44480 47860 44492
rect 47912 44480 47918 44532
rect 12618 44412 12624 44464
rect 12676 44452 12682 44464
rect 27709 44455 27767 44461
rect 12676 44424 27660 44452
rect 12676 44412 12682 44424
rect 13817 44387 13875 44393
rect 13817 44384 13829 44387
rect 12544 44356 13829 44384
rect 12253 44347 12311 44353
rect 13817 44353 13829 44356
rect 13863 44384 13875 44387
rect 14369 44387 14427 44393
rect 14369 44384 14381 44387
rect 13863 44356 14381 44384
rect 13863 44353 13875 44356
rect 13817 44347 13875 44353
rect 14369 44353 14381 44356
rect 14415 44384 14427 44387
rect 19518 44384 19524 44396
rect 14415 44356 19524 44384
rect 14415 44353 14427 44356
rect 14369 44347 14427 44353
rect 19518 44344 19524 44356
rect 19576 44344 19582 44396
rect 20162 44384 20168 44396
rect 20123 44356 20168 44384
rect 20162 44344 20168 44356
rect 20220 44344 20226 44396
rect 20254 44344 20260 44396
rect 20312 44384 20318 44396
rect 20349 44387 20407 44393
rect 20349 44384 20361 44387
rect 20312 44356 20361 44384
rect 20312 44344 20318 44356
rect 20349 44353 20361 44356
rect 20395 44353 20407 44387
rect 20349 44347 20407 44353
rect 20441 44387 20499 44393
rect 20441 44353 20453 44387
rect 20487 44384 20499 44387
rect 20717 44387 20775 44393
rect 20487 44356 20668 44384
rect 20487 44353 20499 44356
rect 20441 44347 20499 44353
rect 9999 44288 11836 44316
rect 11885 44319 11943 44325
rect 9999 44285 10011 44288
rect 9953 44279 10011 44285
rect 11885 44285 11897 44319
rect 11931 44316 11943 44319
rect 12434 44316 12440 44328
rect 11931 44288 12440 44316
rect 11931 44285 11943 44288
rect 11885 44279 11943 44285
rect 12434 44276 12440 44288
rect 12492 44316 12498 44328
rect 13170 44316 13176 44328
rect 12492 44288 13176 44316
rect 12492 44276 12498 44288
rect 13170 44276 13176 44288
rect 13228 44276 13234 44328
rect 15930 44276 15936 44328
rect 15988 44316 15994 44328
rect 19426 44316 19432 44328
rect 15988 44288 19432 44316
rect 15988 44276 15994 44288
rect 19426 44276 19432 44288
rect 19484 44276 19490 44328
rect 20530 44316 20536 44328
rect 19628 44288 19840 44316
rect 20491 44288 20536 44316
rect 8113 44251 8171 44257
rect 8113 44217 8125 44251
rect 8159 44248 8171 44251
rect 19628 44248 19656 44288
rect 8159 44220 19656 44248
rect 19812 44248 19840 44288
rect 20530 44276 20536 44288
rect 20588 44276 20594 44328
rect 20640 44316 20668 44356
rect 20717 44353 20729 44387
rect 20763 44384 20775 44387
rect 22094 44384 22100 44396
rect 20763 44356 22100 44384
rect 20763 44353 20775 44356
rect 20717 44347 20775 44353
rect 22094 44344 22100 44356
rect 22152 44344 22158 44396
rect 22278 44384 22284 44396
rect 22239 44356 22284 44384
rect 22278 44344 22284 44356
rect 22336 44344 22342 44396
rect 23017 44387 23075 44393
rect 23017 44353 23029 44387
rect 23063 44384 23075 44387
rect 23566 44384 23572 44396
rect 23063 44356 23572 44384
rect 23063 44353 23075 44356
rect 23017 44347 23075 44353
rect 21266 44316 21272 44328
rect 20640 44288 21272 44316
rect 21266 44276 21272 44288
rect 21324 44276 21330 44328
rect 22186 44276 22192 44328
rect 22244 44316 22250 44328
rect 23032 44316 23060 44347
rect 23566 44344 23572 44356
rect 23624 44344 23630 44396
rect 23750 44384 23756 44396
rect 23711 44356 23756 44384
rect 23750 44344 23756 44356
rect 23808 44384 23814 44396
rect 24762 44384 24768 44396
rect 23808 44356 24768 44384
rect 23808 44344 23814 44356
rect 24762 44344 24768 44356
rect 24820 44344 24826 44396
rect 24854 44344 24860 44396
rect 24912 44384 24918 44396
rect 25041 44387 25099 44393
rect 25041 44384 25053 44387
rect 24912 44356 25053 44384
rect 24912 44344 24918 44356
rect 25041 44353 25053 44356
rect 25087 44353 25099 44387
rect 25041 44347 25099 44353
rect 25130 44344 25136 44396
rect 25188 44384 25194 44396
rect 25297 44387 25355 44393
rect 25297 44384 25309 44387
rect 25188 44356 25309 44384
rect 25188 44344 25194 44356
rect 25297 44353 25309 44356
rect 25343 44353 25355 44387
rect 25297 44347 25355 44353
rect 27338 44344 27344 44396
rect 27396 44384 27402 44396
rect 27525 44387 27583 44393
rect 27525 44384 27537 44387
rect 27396 44356 27537 44384
rect 27396 44344 27402 44356
rect 27525 44353 27537 44356
rect 27571 44353 27583 44387
rect 27632 44384 27660 44424
rect 27709 44421 27721 44455
rect 27755 44452 27767 44455
rect 28718 44452 28724 44464
rect 27755 44424 28724 44452
rect 27755 44421 27767 44424
rect 27709 44415 27767 44421
rect 28718 44412 28724 44424
rect 28776 44412 28782 44464
rect 30466 44452 30472 44464
rect 30427 44424 30472 44452
rect 30466 44412 30472 44424
rect 30524 44412 30530 44464
rect 31754 44452 31760 44464
rect 30760 44424 31760 44452
rect 29086 44386 29092 44396
rect 28966 44384 29092 44386
rect 27632 44358 29092 44384
rect 27632 44356 28994 44358
rect 27525 44347 27583 44353
rect 29086 44344 29092 44358
rect 29144 44344 29150 44396
rect 30670 44387 30728 44393
rect 30670 44384 30682 44387
rect 30668 44354 30682 44384
rect 30670 44353 30682 44354
rect 30716 44382 30728 44387
rect 30760 44382 30788 44424
rect 31754 44412 31760 44424
rect 31812 44412 31818 44464
rect 34241 44455 34299 44461
rect 34241 44421 34253 44455
rect 34287 44452 34299 44455
rect 34330 44452 34336 44464
rect 34287 44424 34336 44452
rect 34287 44421 34299 44424
rect 34241 44415 34299 44421
rect 34330 44412 34336 44424
rect 34388 44412 34394 44464
rect 44726 44452 44732 44464
rect 44687 44424 44732 44452
rect 44726 44412 44732 44424
rect 44784 44412 44790 44464
rect 47670 44452 47676 44464
rect 45296 44424 47676 44452
rect 30926 44384 30932 44396
rect 30716 44354 30788 44382
rect 30887 44356 30932 44384
rect 30716 44353 30728 44354
rect 30670 44347 30728 44353
rect 30926 44344 30932 44356
rect 30984 44344 30990 44396
rect 31033 44390 31091 44395
rect 31033 44389 31156 44390
rect 31033 44355 31045 44389
rect 31079 44362 31156 44389
rect 31079 44355 31091 44362
rect 31033 44349 31091 44355
rect 31128 44328 31156 44362
rect 31202 44344 31208 44396
rect 31260 44384 31266 44396
rect 31260 44356 31305 44384
rect 31260 44344 31266 44356
rect 31386 44344 31392 44396
rect 31444 44384 31450 44396
rect 45296 44393 45324 44424
rect 47670 44412 47676 44424
rect 47728 44412 47734 44464
rect 45281 44387 45339 44393
rect 45281 44384 45293 44387
rect 31444 44356 45293 44384
rect 31444 44344 31450 44356
rect 45281 44353 45293 44356
rect 45327 44353 45339 44387
rect 45281 44347 45339 44353
rect 45738 44344 45744 44396
rect 45796 44384 45802 44396
rect 45833 44387 45891 44393
rect 45833 44384 45845 44387
rect 45796 44356 45845 44384
rect 45796 44344 45802 44356
rect 45833 44353 45845 44356
rect 45879 44353 45891 44387
rect 45833 44347 45891 44353
rect 46934 44344 46940 44396
rect 46992 44384 46998 44396
rect 47857 44387 47915 44393
rect 47857 44384 47869 44387
rect 46992 44356 47869 44384
rect 46992 44344 46998 44356
rect 47857 44353 47869 44356
rect 47903 44353 47915 44387
rect 47857 44347 47915 44353
rect 22244 44288 23060 44316
rect 22244 44276 22250 44288
rect 23474 44276 23480 44328
rect 23532 44316 23538 44328
rect 24670 44316 24676 44328
rect 23532 44288 24676 44316
rect 23532 44276 23538 44288
rect 24670 44276 24676 44288
rect 24728 44276 24734 44328
rect 28074 44276 28080 44328
rect 28132 44316 28138 44328
rect 28353 44319 28411 44325
rect 28353 44316 28365 44319
rect 28132 44288 28365 44316
rect 28132 44276 28138 44288
rect 28353 44285 28365 44288
rect 28399 44285 28411 44319
rect 28353 44279 28411 44285
rect 28629 44319 28687 44325
rect 28629 44285 28641 44319
rect 28675 44316 28687 44319
rect 28994 44316 29000 44328
rect 28675 44288 29000 44316
rect 28675 44285 28687 44288
rect 28629 44279 28687 44285
rect 28994 44276 29000 44288
rect 29052 44276 29058 44328
rect 30190 44276 30196 44328
rect 30248 44316 30254 44328
rect 30837 44319 30895 44325
rect 30837 44316 30849 44319
rect 30248 44288 30849 44316
rect 30248 44276 30254 44288
rect 30837 44285 30849 44288
rect 30883 44285 30895 44319
rect 30837 44279 30895 44285
rect 31110 44276 31116 44328
rect 31168 44316 31174 44328
rect 31294 44316 31300 44328
rect 31168 44288 31300 44316
rect 31168 44276 31174 44288
rect 31294 44276 31300 44288
rect 31352 44276 31358 44328
rect 30742 44248 30748 44260
rect 19812 44220 25084 44248
rect 8159 44217 8171 44220
rect 8113 44211 8171 44217
rect 7377 44183 7435 44189
rect 7377 44180 7389 44183
rect 6512 44152 7389 44180
rect 6512 44140 6518 44152
rect 7377 44149 7389 44152
rect 7423 44149 7435 44183
rect 7377 44143 7435 44149
rect 10778 44140 10784 44192
rect 10836 44180 10842 44192
rect 10873 44183 10931 44189
rect 10873 44180 10885 44183
rect 10836 44152 10885 44180
rect 10836 44140 10842 44152
rect 10873 44149 10885 44152
rect 10919 44149 10931 44183
rect 10873 44143 10931 44149
rect 11517 44183 11575 44189
rect 11517 44149 11529 44183
rect 11563 44180 11575 44183
rect 11606 44180 11612 44192
rect 11563 44152 11612 44180
rect 11563 44149 11575 44152
rect 11517 44143 11575 44149
rect 11606 44140 11612 44152
rect 11664 44140 11670 44192
rect 12805 44183 12863 44189
rect 12805 44149 12817 44183
rect 12851 44180 12863 44183
rect 13262 44180 13268 44192
rect 12851 44152 13268 44180
rect 12851 44149 12863 44152
rect 12805 44143 12863 44149
rect 13262 44140 13268 44152
rect 13320 44140 13326 44192
rect 16761 44183 16819 44189
rect 16761 44149 16773 44183
rect 16807 44180 16819 44183
rect 17218 44180 17224 44192
rect 16807 44152 17224 44180
rect 16807 44149 16819 44152
rect 16761 44143 16819 44149
rect 17218 44140 17224 44152
rect 17276 44140 17282 44192
rect 17957 44183 18015 44189
rect 17957 44149 17969 44183
rect 18003 44180 18015 44183
rect 18141 44183 18199 44189
rect 18141 44180 18153 44183
rect 18003 44152 18153 44180
rect 18003 44149 18015 44152
rect 17957 44143 18015 44149
rect 18141 44149 18153 44152
rect 18187 44180 18199 44183
rect 18782 44180 18788 44192
rect 18187 44152 18788 44180
rect 18187 44149 18199 44152
rect 18141 44143 18199 44149
rect 18782 44140 18788 44152
rect 18840 44140 18846 44192
rect 18969 44183 19027 44189
rect 18969 44149 18981 44183
rect 19015 44180 19027 44183
rect 19518 44180 19524 44192
rect 19015 44152 19524 44180
rect 19015 44149 19027 44152
rect 18969 44143 19027 44149
rect 19518 44140 19524 44152
rect 19576 44180 19582 44192
rect 22002 44180 22008 44192
rect 19576 44152 22008 44180
rect 19576 44140 19582 44152
rect 22002 44140 22008 44152
rect 22060 44140 22066 44192
rect 22373 44183 22431 44189
rect 22373 44149 22385 44183
rect 22419 44180 22431 44183
rect 23474 44180 23480 44192
rect 22419 44152 23480 44180
rect 22419 44149 22431 44152
rect 22373 44143 22431 44149
rect 23474 44140 23480 44152
rect 23532 44140 23538 44192
rect 23658 44140 23664 44192
rect 23716 44180 23722 44192
rect 23934 44180 23940 44192
rect 23716 44152 23940 44180
rect 23716 44140 23722 44152
rect 23934 44140 23940 44152
rect 23992 44140 23998 44192
rect 24305 44183 24363 44189
rect 24305 44149 24317 44183
rect 24351 44180 24363 44183
rect 24578 44180 24584 44192
rect 24351 44152 24584 44180
rect 24351 44149 24363 44152
rect 24305 44143 24363 44149
rect 24578 44140 24584 44152
rect 24636 44140 24642 44192
rect 25056 44180 25084 44220
rect 25976 44220 30748 44248
rect 25976 44180 26004 44220
rect 30742 44208 30748 44220
rect 30800 44208 30806 44260
rect 31202 44208 31208 44260
rect 31260 44248 31266 44260
rect 44358 44248 44364 44260
rect 31260 44220 44364 44248
rect 31260 44208 31266 44220
rect 44358 44208 44364 44220
rect 44416 44208 44422 44260
rect 26418 44180 26424 44192
rect 25056 44152 26004 44180
rect 26379 44152 26424 44180
rect 26418 44140 26424 44152
rect 26476 44140 26482 44192
rect 28074 44140 28080 44192
rect 28132 44180 28138 44192
rect 29641 44183 29699 44189
rect 29641 44180 29653 44183
rect 28132 44152 29653 44180
rect 28132 44140 28138 44152
rect 29641 44149 29653 44152
rect 29687 44180 29699 44183
rect 30098 44180 30104 44192
rect 29687 44152 30104 44180
rect 29687 44149 29699 44152
rect 29641 44143 29699 44149
rect 30098 44140 30104 44152
rect 30156 44140 30162 44192
rect 34885 44183 34943 44189
rect 34885 44149 34897 44183
rect 34931 44180 34943 44183
rect 35618 44180 35624 44192
rect 34931 44152 35624 44180
rect 34931 44149 34943 44152
rect 34885 44143 34943 44149
rect 35618 44140 35624 44152
rect 35676 44140 35682 44192
rect 46934 44180 46940 44192
rect 46895 44152 46940 44180
rect 46934 44140 46940 44152
rect 46992 44140 46998 44192
rect 48038 44180 48044 44192
rect 47999 44152 48044 44180
rect 48038 44140 48044 44152
rect 48096 44140 48102 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 1857 43979 1915 43985
rect 1857 43945 1869 43979
rect 1903 43976 1915 43979
rect 2866 43976 2872 43988
rect 1903 43948 2872 43976
rect 1903 43945 1915 43948
rect 1857 43939 1915 43945
rect 2866 43936 2872 43948
rect 2924 43936 2930 43988
rect 5442 43936 5448 43988
rect 5500 43976 5506 43988
rect 5905 43979 5963 43985
rect 5905 43976 5917 43979
rect 5500 43948 5917 43976
rect 5500 43936 5506 43948
rect 5905 43945 5917 43948
rect 5951 43976 5963 43979
rect 11146 43976 11152 43988
rect 5951 43948 11152 43976
rect 5951 43945 5963 43948
rect 5905 43939 5963 43945
rect 11146 43936 11152 43948
rect 11204 43976 11210 43988
rect 12713 43979 12771 43985
rect 11204 43948 11928 43976
rect 11204 43936 11210 43948
rect 3878 43908 3884 43920
rect 3791 43880 3884 43908
rect 3878 43868 3884 43880
rect 3936 43908 3942 43920
rect 4614 43908 4620 43920
rect 3936 43880 4620 43908
rect 3936 43868 3942 43880
rect 4614 43868 4620 43880
rect 4672 43868 4678 43920
rect 7006 43868 7012 43920
rect 7064 43908 7070 43920
rect 7561 43911 7619 43917
rect 7561 43908 7573 43911
rect 7064 43880 7573 43908
rect 7064 43868 7070 43880
rect 7561 43877 7573 43880
rect 7607 43877 7619 43911
rect 7561 43871 7619 43877
rect 7668 43880 9536 43908
rect 3237 43843 3295 43849
rect 3237 43809 3249 43843
rect 3283 43840 3295 43843
rect 4982 43840 4988 43852
rect 3283 43812 4988 43840
rect 3283 43809 3295 43812
rect 3237 43803 3295 43809
rect 4982 43800 4988 43812
rect 5040 43800 5046 43852
rect 2038 43732 2044 43784
rect 2096 43772 2102 43784
rect 7668 43772 7696 43880
rect 8202 43800 8208 43852
rect 8260 43840 8266 43852
rect 8297 43843 8355 43849
rect 8297 43840 8309 43843
rect 8260 43812 8309 43840
rect 8260 43800 8266 43812
rect 8297 43809 8309 43812
rect 8343 43840 8355 43843
rect 8343 43812 9444 43840
rect 8343 43809 8355 43812
rect 8297 43803 8355 43809
rect 2096 43744 7696 43772
rect 2096 43732 2102 43744
rect 2958 43704 2964 43716
rect 3016 43713 3022 43716
rect 2928 43676 2964 43704
rect 2958 43664 2964 43676
rect 3016 43667 3028 43713
rect 3016 43664 3022 43667
rect 3510 43664 3516 43716
rect 3568 43704 3574 43716
rect 9416 43713 9444 43812
rect 4893 43707 4951 43713
rect 4893 43704 4905 43707
rect 3568 43676 4905 43704
rect 3568 43664 3574 43676
rect 4893 43673 4905 43676
rect 4939 43673 4951 43707
rect 4893 43667 4951 43673
rect 7745 43707 7803 43713
rect 7745 43673 7757 43707
rect 7791 43704 7803 43707
rect 9401 43707 9459 43713
rect 7791 43676 8340 43704
rect 7791 43673 7803 43676
rect 7745 43667 7803 43673
rect 4433 43639 4491 43645
rect 4433 43605 4445 43639
rect 4479 43636 4491 43639
rect 4798 43636 4804 43648
rect 4479 43608 4804 43636
rect 4479 43605 4491 43608
rect 4433 43599 4491 43605
rect 4798 43596 4804 43608
rect 4856 43596 4862 43648
rect 8312 43636 8340 43676
rect 9401 43673 9413 43707
rect 9447 43673 9459 43707
rect 9508 43704 9536 43880
rect 11900 43849 11928 43948
rect 12713 43945 12725 43979
rect 12759 43976 12771 43979
rect 46934 43976 46940 43988
rect 12759 43948 46940 43976
rect 12759 43945 12771 43948
rect 12713 43939 12771 43945
rect 46934 43936 46940 43948
rect 46992 43936 46998 43988
rect 47210 43936 47216 43988
rect 47268 43976 47274 43988
rect 47489 43979 47547 43985
rect 47489 43976 47501 43979
rect 47268 43948 47501 43976
rect 47268 43936 47274 43948
rect 47489 43945 47501 43948
rect 47535 43945 47547 43979
rect 47489 43939 47547 43945
rect 47946 43936 47952 43988
rect 48004 43976 48010 43988
rect 48041 43979 48099 43985
rect 48041 43976 48053 43979
rect 48004 43948 48053 43976
rect 48004 43936 48010 43948
rect 48041 43945 48053 43948
rect 48087 43945 48099 43979
rect 48041 43939 48099 43945
rect 35066 43908 35072 43920
rect 12406 43880 35072 43908
rect 11885 43843 11943 43849
rect 11885 43809 11897 43843
rect 11931 43840 11943 43843
rect 11974 43840 11980 43852
rect 11931 43812 11980 43840
rect 11931 43809 11943 43812
rect 11885 43803 11943 43809
rect 11974 43800 11980 43812
rect 12032 43800 12038 43852
rect 12406 43840 12434 43880
rect 35066 43868 35072 43880
rect 35124 43868 35130 43920
rect 37737 43911 37795 43917
rect 37737 43877 37749 43911
rect 37783 43908 37795 43911
rect 38654 43908 38660 43920
rect 37783 43880 38660 43908
rect 37783 43877 37795 43880
rect 37737 43871 37795 43877
rect 38654 43868 38660 43880
rect 38712 43908 38718 43920
rect 39758 43908 39764 43920
rect 38712 43880 39764 43908
rect 38712 43868 38718 43880
rect 39758 43868 39764 43880
rect 39816 43868 39822 43920
rect 45646 43908 45652 43920
rect 45607 43880 45652 43908
rect 45646 43868 45652 43880
rect 45704 43868 45710 43920
rect 46198 43908 46204 43920
rect 46159 43880 46204 43908
rect 46198 43868 46204 43880
rect 46256 43868 46262 43920
rect 46658 43868 46664 43920
rect 46716 43908 46722 43920
rect 46753 43911 46811 43917
rect 46753 43908 46765 43911
rect 46716 43880 46765 43908
rect 46716 43868 46722 43880
rect 46753 43877 46765 43880
rect 46799 43877 46811 43911
rect 46753 43871 46811 43877
rect 12084 43812 12434 43840
rect 11606 43732 11612 43784
rect 11664 43781 11670 43784
rect 11664 43772 11676 43781
rect 11664 43744 11709 43772
rect 11664 43735 11676 43744
rect 11664 43732 11670 43735
rect 12084 43704 12112 43812
rect 12894 43800 12900 43852
rect 12952 43840 12958 43852
rect 13081 43843 13139 43849
rect 13081 43840 13093 43843
rect 12952 43812 13093 43840
rect 12952 43800 12958 43812
rect 13081 43809 13093 43812
rect 13127 43809 13139 43843
rect 13081 43803 13139 43809
rect 13170 43800 13176 43852
rect 13228 43840 13234 43852
rect 13228 43812 13273 43840
rect 13228 43800 13234 43812
rect 15102 43800 15108 43852
rect 15160 43840 15166 43852
rect 15565 43843 15623 43849
rect 15565 43840 15577 43843
rect 15160 43812 15577 43840
rect 15160 43800 15166 43812
rect 15565 43809 15577 43812
rect 15611 43809 15623 43843
rect 15565 43803 15623 43809
rect 12158 43732 12164 43784
rect 12216 43772 12222 43784
rect 12805 43775 12863 43781
rect 12805 43772 12817 43775
rect 12216 43744 12817 43772
rect 12216 43732 12222 43744
rect 12805 43741 12817 43744
rect 12851 43741 12863 43775
rect 12805 43735 12863 43741
rect 12989 43775 13047 43781
rect 12989 43741 13001 43775
rect 13035 43741 13047 43775
rect 12989 43735 13047 43741
rect 13357 43775 13415 43781
rect 13357 43741 13369 43775
rect 13403 43772 13415 43775
rect 13814 43772 13820 43784
rect 13403 43744 13820 43772
rect 13403 43741 13415 43744
rect 13357 43735 13415 43741
rect 9508 43676 12112 43704
rect 13004 43704 13032 43735
rect 13814 43732 13820 43744
rect 13872 43732 13878 43784
rect 15580 43772 15608 43803
rect 16666 43800 16672 43852
rect 16724 43840 16730 43852
rect 17037 43843 17095 43849
rect 16724 43812 16896 43840
rect 16724 43800 16730 43812
rect 16758 43772 16764 43784
rect 15580 43744 16764 43772
rect 16758 43732 16764 43744
rect 16816 43732 16822 43784
rect 16868 43781 16896 43812
rect 17037 43809 17049 43843
rect 17083 43840 17095 43843
rect 18322 43840 18328 43852
rect 17083 43812 18328 43840
rect 17083 43809 17095 43812
rect 17037 43803 17095 43809
rect 18322 43800 18328 43812
rect 18380 43800 18386 43852
rect 18598 43800 18604 43852
rect 18656 43840 18662 43852
rect 20073 43843 20131 43849
rect 20073 43840 20085 43843
rect 18656 43812 20085 43840
rect 18656 43800 18662 43812
rect 20073 43809 20085 43812
rect 20119 43840 20131 43843
rect 21174 43840 21180 43852
rect 20119 43812 21180 43840
rect 20119 43809 20131 43812
rect 20073 43803 20131 43809
rect 21174 43800 21180 43812
rect 21232 43800 21238 43852
rect 21266 43800 21272 43852
rect 21324 43840 21330 43852
rect 23477 43843 23535 43849
rect 21324 43812 23428 43840
rect 21324 43800 21330 43812
rect 16853 43775 16911 43781
rect 16853 43741 16865 43775
rect 16899 43741 16911 43775
rect 17126 43772 17132 43784
rect 17087 43744 17132 43772
rect 16853 43735 16911 43741
rect 17126 43732 17132 43744
rect 17184 43732 17190 43784
rect 17218 43732 17224 43784
rect 17276 43772 17282 43784
rect 17276 43744 17321 43772
rect 17276 43732 17282 43744
rect 17402 43732 17408 43784
rect 17460 43772 17466 43784
rect 18046 43772 18052 43784
rect 17460 43744 18052 43772
rect 17460 43732 17466 43744
rect 18046 43732 18052 43744
rect 18104 43772 18110 43784
rect 19797 43775 19855 43781
rect 19797 43772 19809 43775
rect 18104 43744 19809 43772
rect 18104 43732 18110 43744
rect 19797 43741 19809 43744
rect 19843 43772 19855 43775
rect 20162 43772 20168 43784
rect 19843 43744 20168 43772
rect 19843 43741 19855 43744
rect 19797 43735 19855 43741
rect 20162 43732 20168 43744
rect 20220 43732 20226 43784
rect 20254 43732 20260 43784
rect 20312 43772 20318 43784
rect 20625 43775 20683 43781
rect 20625 43772 20637 43775
rect 20312 43744 20637 43772
rect 20312 43732 20318 43744
rect 20625 43741 20637 43744
rect 20671 43772 20683 43775
rect 22186 43772 22192 43784
rect 20671 43744 22192 43772
rect 20671 43741 20683 43744
rect 20625 43735 20683 43741
rect 22186 43732 22192 43744
rect 22244 43732 22250 43784
rect 22922 43732 22928 43784
rect 22980 43772 22986 43784
rect 23293 43775 23351 43781
rect 23293 43772 23305 43775
rect 22980 43744 23305 43772
rect 22980 43732 22986 43744
rect 23293 43741 23305 43744
rect 23339 43741 23351 43775
rect 23293 43735 23351 43741
rect 23400 43766 23428 43812
rect 23477 43809 23489 43843
rect 23523 43840 23535 43843
rect 24762 43840 24768 43852
rect 23523 43812 24768 43840
rect 23523 43809 23535 43812
rect 23477 43803 23535 43809
rect 24762 43800 24768 43812
rect 24820 43800 24826 43852
rect 25130 43840 25136 43852
rect 25091 43812 25136 43840
rect 25130 43800 25136 43812
rect 25188 43800 25194 43852
rect 27338 43840 27344 43852
rect 27299 43812 27344 43840
rect 27338 43800 27344 43812
rect 27396 43800 27402 43852
rect 29822 43840 29828 43852
rect 28460 43812 29828 43840
rect 23566 43772 23572 43784
rect 23492 43766 23572 43772
rect 23400 43744 23572 43766
rect 23400 43738 23520 43744
rect 23566 43732 23572 43744
rect 23624 43732 23630 43784
rect 23661 43775 23719 43781
rect 23661 43741 23673 43775
rect 23707 43772 23719 43775
rect 23750 43772 23756 43784
rect 23707 43744 23756 43772
rect 23707 43741 23719 43744
rect 23661 43735 23719 43741
rect 13262 43704 13268 43716
rect 13004 43676 13268 43704
rect 9401 43667 9459 43673
rect 13262 43664 13268 43676
rect 13320 43664 13326 43716
rect 15746 43704 15752 43716
rect 15707 43676 15752 43704
rect 15746 43664 15752 43676
rect 15804 43664 15810 43716
rect 17494 43664 17500 43716
rect 17552 43704 17558 43716
rect 21361 43707 21419 43713
rect 21361 43704 21373 43707
rect 17552 43676 21373 43704
rect 17552 43664 17558 43676
rect 21361 43673 21373 43676
rect 21407 43704 21419 43707
rect 22278 43704 22284 43716
rect 21407 43676 22284 43704
rect 21407 43673 21419 43676
rect 21361 43667 21419 43673
rect 22278 43664 22284 43676
rect 22336 43664 22342 43716
rect 22649 43707 22707 43713
rect 22649 43673 22661 43707
rect 22695 43704 22707 43707
rect 23676 43704 23704 43735
rect 23750 43732 23756 43744
rect 23808 43732 23814 43784
rect 23842 43732 23848 43784
rect 23900 43772 23906 43784
rect 24397 43775 24455 43781
rect 24397 43772 24409 43775
rect 23900 43744 24409 43772
rect 23900 43732 23906 43744
rect 24397 43741 24409 43744
rect 24443 43741 24455 43775
rect 24578 43772 24584 43784
rect 24539 43744 24584 43772
rect 24397 43735 24455 43741
rect 24578 43732 24584 43744
rect 24636 43732 24642 43784
rect 24670 43732 24676 43784
rect 24728 43772 24734 43784
rect 24949 43775 25007 43781
rect 24728 43744 24773 43772
rect 24728 43732 24734 43744
rect 24949 43741 24961 43775
rect 24995 43772 25007 43775
rect 26418 43772 26424 43784
rect 24995 43744 26424 43772
rect 24995 43741 25007 43744
rect 24949 43735 25007 43741
rect 26418 43732 26424 43744
rect 26476 43732 26482 43784
rect 28460 43781 28488 43812
rect 29822 43800 29828 43812
rect 29880 43800 29886 43852
rect 32398 43800 32404 43852
rect 32456 43840 32462 43852
rect 32944 43843 33002 43849
rect 32944 43840 32956 43843
rect 32456 43812 32956 43840
rect 32456 43800 32462 43812
rect 32944 43809 32956 43812
rect 32990 43809 33002 43843
rect 32944 43803 33002 43809
rect 33318 43800 33324 43852
rect 33376 43840 33382 43852
rect 35437 43843 35495 43849
rect 35437 43840 35449 43843
rect 33376 43812 35449 43840
rect 33376 43800 33382 43812
rect 35437 43809 35449 43812
rect 35483 43840 35495 43843
rect 35894 43840 35900 43852
rect 35483 43812 35900 43840
rect 35483 43809 35495 43812
rect 35437 43803 35495 43809
rect 35894 43800 35900 43812
rect 35952 43800 35958 43852
rect 35986 43800 35992 43852
rect 36044 43840 36050 43852
rect 36357 43843 36415 43849
rect 36357 43840 36369 43843
rect 36044 43812 36369 43840
rect 36044 43800 36050 43812
rect 36357 43809 36369 43812
rect 36403 43809 36415 43843
rect 36357 43803 36415 43809
rect 28445 43775 28503 43781
rect 28445 43741 28457 43775
rect 28491 43741 28503 43775
rect 28626 43772 28632 43784
rect 28587 43744 28632 43772
rect 28445 43735 28503 43741
rect 28626 43732 28632 43744
rect 28684 43732 28690 43784
rect 28718 43775 28776 43781
rect 28718 43741 28730 43775
rect 28764 43741 28776 43775
rect 28718 43735 28776 43741
rect 28813 43777 28871 43783
rect 28813 43743 28825 43777
rect 28859 43743 28871 43777
rect 28994 43772 29000 43784
rect 28955 43744 29000 43772
rect 28813 43737 28871 43743
rect 22695 43676 23704 43704
rect 24688 43704 24716 43732
rect 28534 43704 28540 43716
rect 24688 43676 28540 43704
rect 22695 43673 22707 43676
rect 22649 43667 22707 43673
rect 28534 43664 28540 43676
rect 28592 43704 28598 43716
rect 28733 43704 28761 43735
rect 28592 43676 28761 43704
rect 28828 43704 28856 43737
rect 28994 43732 29000 43744
rect 29052 43732 29058 43784
rect 31570 43732 31576 43784
rect 31628 43772 31634 43784
rect 32677 43775 32735 43781
rect 32677 43772 32689 43775
rect 31628 43744 32689 43772
rect 31628 43732 31634 43744
rect 32677 43741 32689 43744
rect 32723 43741 32735 43775
rect 32858 43774 32864 43784
rect 32677 43735 32735 43741
rect 32784 43746 32864 43774
rect 32784 43704 32812 43746
rect 32858 43732 32864 43746
rect 32916 43772 32922 43784
rect 33045 43775 33103 43781
rect 32916 43744 33009 43772
rect 32916 43732 32922 43744
rect 33045 43741 33057 43775
rect 33091 43741 33103 43775
rect 33045 43735 33103 43741
rect 28828 43676 29316 43704
rect 28592 43664 28598 43676
rect 29288 43648 29316 43676
rect 31956 43676 32812 43704
rect 33060 43704 33088 43735
rect 33134 43732 33140 43784
rect 33192 43772 33198 43784
rect 33229 43775 33287 43781
rect 33229 43772 33241 43775
rect 33192 43744 33241 43772
rect 33192 43732 33198 43744
rect 33229 43741 33241 43744
rect 33275 43741 33287 43775
rect 35161 43775 35219 43781
rect 35161 43774 35173 43775
rect 33229 43735 33287 43741
rect 35084 43746 35173 43774
rect 34054 43704 34060 43716
rect 33060 43676 34060 43704
rect 9493 43639 9551 43645
rect 9493 43636 9505 43639
rect 8312 43608 9505 43636
rect 9493 43605 9505 43608
rect 9539 43636 9551 43639
rect 10226 43636 10232 43648
rect 9539 43608 10232 43636
rect 9539 43605 9551 43608
rect 9493 43599 9551 43605
rect 10226 43596 10232 43608
rect 10284 43596 10290 43648
rect 10505 43639 10563 43645
rect 10505 43605 10517 43639
rect 10551 43636 10563 43639
rect 11698 43636 11704 43648
rect 10551 43608 11704 43636
rect 10551 43605 10563 43608
rect 10505 43599 10563 43605
rect 11698 43596 11704 43608
rect 11756 43596 11762 43648
rect 11790 43596 11796 43648
rect 11848 43636 11854 43648
rect 12713 43639 12771 43645
rect 12713 43636 12725 43639
rect 11848 43608 12725 43636
rect 11848 43596 11854 43608
rect 12713 43605 12725 43608
rect 12759 43605 12771 43639
rect 12713 43599 12771 43605
rect 13354 43596 13360 43648
rect 13412 43636 13418 43648
rect 13541 43639 13599 43645
rect 13541 43636 13553 43639
rect 13412 43608 13553 43636
rect 13412 43596 13418 43608
rect 13541 43605 13553 43608
rect 13587 43605 13599 43639
rect 13541 43599 13599 43605
rect 13630 43596 13636 43648
rect 13688 43636 13694 43648
rect 14185 43639 14243 43645
rect 14185 43636 14197 43639
rect 13688 43608 14197 43636
rect 13688 43596 13694 43608
rect 14185 43605 14197 43608
rect 14231 43636 14243 43639
rect 15194 43636 15200 43648
rect 14231 43608 15200 43636
rect 14231 43605 14243 43608
rect 14185 43599 14243 43605
rect 15194 43596 15200 43608
rect 15252 43596 15258 43648
rect 16669 43639 16727 43645
rect 16669 43605 16681 43639
rect 16715 43636 16727 43639
rect 16942 43636 16948 43648
rect 16715 43608 16948 43636
rect 16715 43605 16727 43608
rect 16669 43599 16727 43605
rect 16942 43596 16948 43608
rect 17000 43596 17006 43648
rect 21266 43636 21272 43648
rect 21227 43608 21272 43636
rect 21266 43596 21272 43608
rect 21324 43596 21330 43648
rect 23109 43639 23167 43645
rect 23109 43605 23121 43639
rect 23155 43636 23167 43639
rect 23198 43636 23204 43648
rect 23155 43608 23204 43636
rect 23155 43605 23167 43608
rect 23109 43599 23167 43605
rect 23198 43596 23204 43608
rect 23256 43596 23262 43648
rect 23290 43596 23296 43648
rect 23348 43636 23354 43648
rect 28074 43636 28080 43648
rect 23348 43608 28080 43636
rect 23348 43596 23354 43608
rect 28074 43596 28080 43608
rect 28132 43596 28138 43648
rect 28258 43636 28264 43648
rect 28219 43608 28264 43636
rect 28258 43596 28264 43608
rect 28316 43596 28322 43648
rect 29270 43596 29276 43648
rect 29328 43636 29334 43648
rect 29549 43639 29607 43645
rect 29549 43636 29561 43639
rect 29328 43608 29561 43636
rect 29328 43596 29334 43608
rect 29549 43605 29561 43608
rect 29595 43605 29607 43639
rect 30374 43636 30380 43648
rect 30335 43608 30380 43636
rect 29549 43599 29607 43605
rect 30374 43596 30380 43608
rect 30432 43636 30438 43648
rect 31110 43636 31116 43648
rect 30432 43608 31116 43636
rect 30432 43596 30438 43608
rect 31110 43596 31116 43608
rect 31168 43596 31174 43648
rect 31846 43596 31852 43648
rect 31904 43636 31910 43648
rect 31956 43645 31984 43676
rect 34054 43664 34060 43676
rect 34112 43664 34118 43716
rect 35084 43704 35112 43746
rect 35161 43741 35173 43746
rect 35207 43741 35219 43775
rect 35161 43735 35219 43741
rect 35250 43732 35256 43784
rect 35308 43772 35314 43784
rect 35345 43775 35403 43781
rect 35345 43772 35357 43775
rect 35308 43744 35357 43772
rect 35308 43732 35314 43744
rect 35345 43741 35357 43744
rect 35391 43741 35403 43775
rect 35345 43735 35403 43741
rect 35529 43775 35587 43781
rect 35529 43741 35541 43775
rect 35575 43772 35587 43775
rect 35618 43772 35624 43784
rect 35575 43744 35624 43772
rect 35575 43741 35587 43744
rect 35529 43735 35587 43741
rect 35618 43732 35624 43744
rect 35676 43732 35682 43784
rect 35710 43732 35716 43784
rect 35768 43772 35774 43784
rect 47302 43772 47308 43784
rect 35768 43744 35813 43772
rect 47263 43744 47308 43772
rect 35768 43732 35774 43744
rect 47302 43732 47308 43744
rect 47360 43732 47366 43784
rect 36262 43704 36268 43716
rect 35084 43676 36268 43704
rect 36262 43664 36268 43676
rect 36320 43664 36326 43716
rect 36354 43664 36360 43716
rect 36412 43704 36418 43716
rect 36602 43707 36660 43713
rect 36602 43704 36614 43707
rect 36412 43676 36614 43704
rect 36412 43664 36418 43676
rect 36602 43673 36614 43676
rect 36648 43673 36660 43707
rect 36602 43667 36660 43673
rect 31941 43639 31999 43645
rect 31941 43636 31953 43639
rect 31904 43608 31953 43636
rect 31904 43596 31910 43608
rect 31941 43605 31953 43608
rect 31987 43605 31999 43639
rect 32490 43636 32496 43648
rect 32451 43608 32496 43636
rect 31941 43599 31999 43605
rect 32490 43596 32496 43608
rect 32548 43596 32554 43648
rect 34790 43596 34796 43648
rect 34848 43636 34854 43648
rect 34977 43639 35035 43645
rect 34977 43636 34989 43639
rect 34848 43608 34989 43636
rect 34848 43596 34854 43608
rect 34977 43605 34989 43608
rect 35023 43605 35035 43639
rect 34977 43599 35035 43605
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 2516 43404 2774 43432
rect 2314 43296 2320 43308
rect 2275 43268 2320 43296
rect 2314 43256 2320 43268
rect 2372 43256 2378 43308
rect 2516 43305 2544 43404
rect 2746 43364 2774 43404
rect 2958 43392 2964 43444
rect 3016 43432 3022 43444
rect 3053 43435 3111 43441
rect 3053 43432 3065 43435
rect 3016 43404 3065 43432
rect 3016 43392 3022 43404
rect 3053 43401 3065 43404
rect 3099 43401 3111 43435
rect 3053 43395 3111 43401
rect 3697 43435 3755 43441
rect 3697 43401 3709 43435
rect 3743 43432 3755 43435
rect 5810 43432 5816 43444
rect 3743 43404 5672 43432
rect 5723 43404 5816 43432
rect 3743 43401 3755 43404
rect 3697 43395 3755 43401
rect 5442 43364 5448 43376
rect 2746 43336 3556 43364
rect 3528 43308 3556 43336
rect 4448 43336 5448 43364
rect 2501 43299 2559 43305
rect 2501 43265 2513 43299
rect 2547 43265 2559 43299
rect 2682 43296 2688 43308
rect 2643 43268 2688 43296
rect 2501 43259 2559 43265
rect 2516 43228 2544 43259
rect 2682 43256 2688 43268
rect 2740 43256 2746 43308
rect 2866 43296 2872 43308
rect 2827 43268 2872 43296
rect 2866 43256 2872 43268
rect 2924 43256 2930 43308
rect 3510 43296 3516 43308
rect 3471 43268 3516 43296
rect 3510 43256 3516 43268
rect 3568 43256 3574 43308
rect 4448 43305 4476 43336
rect 5442 43324 5448 43336
rect 5500 43324 5506 43376
rect 5644 43364 5672 43404
rect 5810 43392 5816 43404
rect 5868 43432 5874 43444
rect 6362 43432 6368 43444
rect 5868 43404 6368 43432
rect 5868 43392 5874 43404
rect 6362 43392 6368 43404
rect 6420 43392 6426 43444
rect 8110 43432 8116 43444
rect 8071 43404 8116 43432
rect 8110 43392 8116 43404
rect 8168 43392 8174 43444
rect 9674 43392 9680 43444
rect 9732 43432 9738 43444
rect 9953 43435 10011 43441
rect 9953 43432 9965 43435
rect 9732 43404 9965 43432
rect 9732 43392 9738 43404
rect 9953 43401 9965 43404
rect 9999 43401 10011 43435
rect 9953 43395 10011 43401
rect 10042 43392 10048 43444
rect 10100 43432 10106 43444
rect 10597 43435 10655 43441
rect 10597 43432 10609 43435
rect 10100 43404 10609 43432
rect 10100 43392 10106 43404
rect 10597 43401 10609 43404
rect 10643 43401 10655 43435
rect 10597 43395 10655 43401
rect 11992 43404 13768 43432
rect 11790 43364 11796 43376
rect 5644 43336 11796 43364
rect 11790 43324 11796 43336
rect 11848 43324 11854 43376
rect 4706 43305 4712 43308
rect 4433 43299 4491 43305
rect 4433 43265 4445 43299
rect 4479 43265 4491 43299
rect 4433 43259 4491 43265
rect 4700 43259 4712 43305
rect 4764 43296 4770 43308
rect 4764 43268 4800 43296
rect 4706 43256 4712 43259
rect 4764 43256 4770 43268
rect 4982 43256 4988 43308
rect 5040 43296 5046 43308
rect 6733 43299 6791 43305
rect 6733 43296 6745 43299
rect 5040 43268 6745 43296
rect 5040 43256 5046 43268
rect 6733 43265 6745 43268
rect 6779 43296 6791 43299
rect 6822 43296 6828 43308
rect 6779 43268 6828 43296
rect 6779 43265 6791 43268
rect 6733 43259 6791 43265
rect 6822 43256 6828 43268
rect 6880 43256 6886 43308
rect 7006 43305 7012 43308
rect 7000 43259 7012 43305
rect 7064 43296 7070 43308
rect 8938 43296 8944 43308
rect 7064 43268 7100 43296
rect 8899 43268 8944 43296
rect 7006 43256 7012 43259
rect 7064 43256 7070 43268
rect 8938 43256 8944 43268
rect 8996 43296 9002 43308
rect 9861 43299 9919 43305
rect 9861 43296 9873 43299
rect 8996 43268 9873 43296
rect 8996 43256 9002 43268
rect 9861 43265 9873 43268
rect 9907 43265 9919 43299
rect 9861 43259 9919 43265
rect 10502 43256 10508 43308
rect 10560 43296 10566 43308
rect 11992 43305 12020 43404
rect 12158 43364 12164 43376
rect 12119 43336 12164 43364
rect 12158 43324 12164 43336
rect 12216 43324 12222 43376
rect 13630 43364 13636 43376
rect 13096 43336 13636 43364
rect 10689 43299 10747 43305
rect 10689 43296 10701 43299
rect 10560 43268 10701 43296
rect 10560 43256 10566 43268
rect 10689 43265 10701 43268
rect 10735 43296 10747 43299
rect 11977 43299 12035 43305
rect 11977 43296 11989 43299
rect 10735 43268 11989 43296
rect 10735 43265 10747 43268
rect 10689 43259 10747 43265
rect 11977 43265 11989 43268
rect 12023 43265 12035 43299
rect 11977 43259 12035 43265
rect 12066 43256 12072 43308
rect 12124 43296 12130 43308
rect 13096 43305 13124 43336
rect 13630 43324 13636 43336
rect 13688 43324 13694 43376
rect 13354 43305 13360 43308
rect 13081 43299 13139 43305
rect 13081 43296 13093 43299
rect 12124 43268 13093 43296
rect 12124 43256 12130 43268
rect 13081 43265 13093 43268
rect 13127 43265 13139 43299
rect 13348 43296 13360 43305
rect 13315 43268 13360 43296
rect 13081 43259 13139 43265
rect 13348 43259 13360 43268
rect 13354 43256 13360 43259
rect 13412 43256 13418 43308
rect 13740 43296 13768 43404
rect 13814 43392 13820 43444
rect 13872 43432 13878 43444
rect 14461 43435 14519 43441
rect 14461 43432 14473 43435
rect 13872 43404 14473 43432
rect 13872 43392 13878 43404
rect 14461 43401 14473 43404
rect 14507 43401 14519 43435
rect 14461 43395 14519 43401
rect 15013 43435 15071 43441
rect 15013 43401 15025 43435
rect 15059 43432 15071 43435
rect 15194 43432 15200 43444
rect 15059 43404 15200 43432
rect 15059 43401 15071 43404
rect 15013 43395 15071 43401
rect 15194 43392 15200 43404
rect 15252 43432 15258 43444
rect 15838 43432 15844 43444
rect 15252 43404 15844 43432
rect 15252 43392 15258 43404
rect 15838 43392 15844 43404
rect 15896 43432 15902 43444
rect 16025 43435 16083 43441
rect 16025 43432 16037 43435
rect 15896 43404 16037 43432
rect 15896 43392 15902 43404
rect 16025 43401 16037 43404
rect 16071 43401 16083 43435
rect 16025 43395 16083 43401
rect 16040 43296 16068 43395
rect 16666 43392 16672 43444
rect 16724 43432 16730 43444
rect 17954 43432 17960 43444
rect 16724 43404 17960 43432
rect 16724 43392 16730 43404
rect 17954 43392 17960 43404
rect 18012 43432 18018 43444
rect 18049 43435 18107 43441
rect 18049 43432 18061 43435
rect 18012 43404 18061 43432
rect 18012 43392 18018 43404
rect 18049 43401 18061 43404
rect 18095 43401 18107 43435
rect 18049 43395 18107 43401
rect 18509 43435 18567 43441
rect 18509 43401 18521 43435
rect 18555 43432 18567 43435
rect 18690 43432 18696 43444
rect 18555 43404 18696 43432
rect 18555 43401 18567 43404
rect 18509 43395 18567 43401
rect 18690 43392 18696 43404
rect 18748 43392 18754 43444
rect 22005 43435 22063 43441
rect 22005 43432 22017 43435
rect 18800 43404 22017 43432
rect 16942 43373 16948 43376
rect 16936 43364 16948 43373
rect 16903 43336 16948 43364
rect 16936 43327 16948 43336
rect 16942 43324 16948 43327
rect 17000 43324 17006 43376
rect 16669 43299 16727 43305
rect 16669 43296 16681 43299
rect 13740 43268 15976 43296
rect 16040 43268 16681 43296
rect 1780 43200 2544 43228
rect 2593 43231 2651 43237
rect 842 43052 848 43104
rect 900 43092 906 43104
rect 1780 43101 1808 43200
rect 2593 43197 2605 43231
rect 2639 43197 2651 43231
rect 15948 43228 15976 43268
rect 16669 43265 16681 43268
rect 16715 43265 16727 43299
rect 18598 43296 18604 43308
rect 16669 43259 16727 43265
rect 16776 43268 18604 43296
rect 16776 43228 16804 43268
rect 18598 43256 18604 43268
rect 18656 43256 18662 43308
rect 15948 43200 16804 43228
rect 2593 43191 2651 43197
rect 2608 43160 2636 43191
rect 2774 43160 2780 43172
rect 2608 43132 2780 43160
rect 2774 43120 2780 43132
rect 2832 43120 2838 43172
rect 7668 43132 12434 43160
rect 1765 43095 1823 43101
rect 1765 43092 1777 43095
rect 900 43064 1777 43092
rect 900 43052 906 43064
rect 1765 43061 1777 43064
rect 1811 43061 1823 43095
rect 1765 43055 1823 43061
rect 4798 43052 4804 43104
rect 4856 43092 4862 43104
rect 7668 43092 7696 43132
rect 9214 43092 9220 43104
rect 4856 43064 7696 43092
rect 9175 43064 9220 43092
rect 4856 43052 4862 43064
rect 9214 43052 9220 43064
rect 9272 43052 9278 43104
rect 12406 43092 12434 43132
rect 18800 43092 18828 43404
rect 22005 43401 22017 43404
rect 22051 43432 22063 43435
rect 23106 43432 23112 43444
rect 22051 43404 23112 43432
rect 22051 43401 22063 43404
rect 22005 43395 22063 43401
rect 23106 43392 23112 43404
rect 23164 43392 23170 43444
rect 23382 43392 23388 43444
rect 23440 43432 23446 43444
rect 24305 43435 24363 43441
rect 24305 43432 24317 43435
rect 23440 43404 24317 43432
rect 23440 43392 23446 43404
rect 24305 43401 24317 43404
rect 24351 43432 24363 43435
rect 24946 43432 24952 43444
rect 24351 43404 24952 43432
rect 24351 43401 24363 43404
rect 24305 43395 24363 43401
rect 24946 43392 24952 43404
rect 25004 43392 25010 43444
rect 26326 43432 26332 43444
rect 26239 43404 26332 43432
rect 26326 43392 26332 43404
rect 26384 43432 26390 43444
rect 27522 43432 27528 43444
rect 26384 43404 27528 43432
rect 26384 43392 26390 43404
rect 27522 43392 27528 43404
rect 27580 43392 27586 43444
rect 29549 43435 29607 43441
rect 29549 43401 29561 43435
rect 29595 43432 29607 43435
rect 29822 43432 29828 43444
rect 29595 43404 29828 43432
rect 29595 43401 29607 43404
rect 29549 43395 29607 43401
rect 29822 43392 29828 43404
rect 29880 43392 29886 43444
rect 30193 43435 30251 43441
rect 30193 43401 30205 43435
rect 30239 43432 30251 43435
rect 33134 43432 33140 43444
rect 30239 43404 33140 43432
rect 30239 43401 30251 43404
rect 30193 43395 30251 43401
rect 33134 43392 33140 43404
rect 33192 43392 33198 43444
rect 33226 43392 33232 43444
rect 33284 43432 33290 43444
rect 33597 43435 33655 43441
rect 33597 43432 33609 43435
rect 33284 43404 33609 43432
rect 33284 43392 33290 43404
rect 33597 43401 33609 43404
rect 33643 43401 33655 43435
rect 35066 43432 35072 43444
rect 35027 43404 35072 43432
rect 33597 43395 33655 43401
rect 35066 43392 35072 43404
rect 35124 43392 35130 43444
rect 36354 43432 36360 43444
rect 36315 43404 36360 43432
rect 36354 43392 36360 43404
rect 36412 43392 36418 43444
rect 20622 43324 20628 43376
rect 20680 43364 20686 43376
rect 23290 43364 23296 43376
rect 20680 43336 20760 43364
rect 20680 43324 20686 43336
rect 19334 43256 19340 43308
rect 19392 43296 19398 43308
rect 19622 43299 19680 43305
rect 19622 43296 19634 43299
rect 19392 43268 19634 43296
rect 19392 43256 19398 43268
rect 19622 43265 19634 43268
rect 19668 43265 19680 43299
rect 19622 43259 19680 43265
rect 20162 43256 20168 43308
rect 20220 43296 20226 43308
rect 20349 43299 20407 43305
rect 20349 43296 20361 43299
rect 20220 43268 20361 43296
rect 20220 43256 20226 43268
rect 20349 43265 20361 43268
rect 20395 43265 20407 43299
rect 20530 43296 20536 43308
rect 20491 43268 20536 43296
rect 20349 43259 20407 43265
rect 20530 43256 20536 43268
rect 20588 43256 20594 43308
rect 20732 43305 20760 43336
rect 22940 43336 23296 43364
rect 20717 43299 20775 43305
rect 20717 43265 20729 43299
rect 20763 43265 20775 43299
rect 20717 43259 20775 43265
rect 20901 43299 20959 43305
rect 20901 43265 20913 43299
rect 20947 43296 20959 43299
rect 21082 43296 21088 43308
rect 20947 43268 21088 43296
rect 20947 43265 20959 43268
rect 20901 43259 20959 43265
rect 21082 43256 21088 43268
rect 21140 43256 21146 43308
rect 21174 43256 21180 43308
rect 21232 43296 21238 43308
rect 21821 43299 21879 43305
rect 21821 43296 21833 43299
rect 21232 43268 21833 43296
rect 21232 43256 21238 43268
rect 21821 43265 21833 43268
rect 21867 43296 21879 43299
rect 21910 43296 21916 43308
rect 21867 43268 21916 43296
rect 21867 43265 21879 43268
rect 21821 43259 21879 43265
rect 21910 43256 21916 43268
rect 21968 43256 21974 43308
rect 22940 43305 22968 43336
rect 23290 43324 23296 43336
rect 23348 43364 23354 43376
rect 24854 43364 24860 43376
rect 23348 43336 24860 43364
rect 23348 43324 23354 43336
rect 24854 43324 24860 43336
rect 24912 43324 24918 43376
rect 28258 43324 28264 43376
rect 28316 43364 28322 43376
rect 28414 43367 28472 43373
rect 28414 43364 28426 43367
rect 28316 43336 28426 43364
rect 28316 43324 28322 43336
rect 28414 43333 28426 43336
rect 28460 43333 28472 43367
rect 30098 43364 30104 43376
rect 30059 43336 30104 43364
rect 28414 43327 28472 43333
rect 30098 43324 30104 43336
rect 30156 43324 30162 43376
rect 32858 43324 32864 43376
rect 32916 43364 32922 43376
rect 33505 43367 33563 43373
rect 33505 43364 33517 43367
rect 32916 43336 33517 43364
rect 32916 43324 32922 43336
rect 33505 43333 33517 43336
rect 33551 43364 33563 43367
rect 34149 43367 34207 43373
rect 34149 43364 34161 43367
rect 33551 43336 34161 43364
rect 33551 43333 33563 43336
rect 33505 43327 33563 43333
rect 34149 43333 34161 43336
rect 34195 43333 34207 43367
rect 35084 43364 35112 43392
rect 35084 43336 35848 43364
rect 34149 43327 34207 43333
rect 23198 43305 23204 43308
rect 22925 43299 22983 43305
rect 22925 43296 22937 43299
rect 22066 43268 22937 43296
rect 19889 43231 19947 43237
rect 19889 43197 19901 43231
rect 19935 43197 19947 43231
rect 20622 43228 20628 43240
rect 20583 43200 20628 43228
rect 19889 43191 19947 43197
rect 19904 43160 19932 43191
rect 20622 43188 20628 43200
rect 20680 43188 20686 43240
rect 20346 43160 20352 43172
rect 19904 43132 20352 43160
rect 12406 43064 18828 43092
rect 19610 43052 19616 43104
rect 19668 43092 19674 43104
rect 19904 43092 19932 43132
rect 20346 43120 20352 43132
rect 20404 43160 20410 43172
rect 22066 43160 22094 43268
rect 22925 43265 22937 43268
rect 22971 43265 22983 43299
rect 23192 43296 23204 43305
rect 23159 43268 23204 43296
rect 22925 43259 22983 43265
rect 23192 43259 23204 43268
rect 23198 43256 23204 43259
rect 23256 43256 23262 43308
rect 24872 43296 24900 43324
rect 25222 43305 25228 43308
rect 24949 43299 25007 43305
rect 24949 43296 24961 43299
rect 24872 43268 24961 43296
rect 24949 43265 24961 43268
rect 24995 43265 25007 43299
rect 24949 43259 25007 43265
rect 25216 43259 25228 43305
rect 25280 43296 25286 43308
rect 28902 43296 28908 43308
rect 25280 43268 25316 43296
rect 28184 43268 28908 43296
rect 25222 43256 25228 43259
rect 25280 43256 25286 43268
rect 27982 43188 27988 43240
rect 28040 43228 28046 43240
rect 28184 43237 28212 43268
rect 28902 43256 28908 43268
rect 28960 43256 28966 43308
rect 31570 43296 31576 43308
rect 31531 43268 31576 43296
rect 31570 43256 31576 43268
rect 31628 43256 31634 43308
rect 32398 43296 32404 43308
rect 32359 43268 32404 43296
rect 32398 43256 32404 43268
rect 32456 43256 32462 43308
rect 33134 43256 33140 43308
rect 33192 43296 33198 43308
rect 35621 43299 35679 43305
rect 35621 43296 35633 43299
rect 33192 43268 35633 43296
rect 33192 43256 33198 43268
rect 35621 43265 35633 43268
rect 35667 43296 35679 43299
rect 35710 43296 35716 43308
rect 35667 43268 35716 43296
rect 35667 43265 35679 43268
rect 35621 43259 35679 43265
rect 35710 43256 35716 43268
rect 35768 43256 35774 43308
rect 35820 43305 35848 43336
rect 35805 43299 35863 43305
rect 35805 43265 35817 43299
rect 35851 43265 35863 43299
rect 35805 43259 35863 43265
rect 35894 43256 35900 43308
rect 35952 43296 35958 43308
rect 36173 43299 36231 43305
rect 35952 43268 35997 43296
rect 35952 43256 35958 43268
rect 36173 43265 36185 43299
rect 36219 43296 36231 43299
rect 38654 43296 38660 43308
rect 36219 43268 38660 43296
rect 36219 43265 36231 43268
rect 36173 43259 36231 43265
rect 38654 43256 38660 43268
rect 38712 43256 38718 43308
rect 46934 43256 46940 43308
rect 46992 43296 46998 43308
rect 47857 43299 47915 43305
rect 47857 43296 47869 43299
rect 46992 43268 47869 43296
rect 46992 43256 46998 43268
rect 47857 43265 47869 43268
rect 47903 43265 47915 43299
rect 47857 43259 47915 43265
rect 28169 43231 28227 43237
rect 28169 43228 28181 43231
rect 28040 43200 28181 43228
rect 28040 43188 28046 43200
rect 28169 43197 28181 43200
rect 28215 43197 28227 43231
rect 28169 43191 28227 43197
rect 31938 43188 31944 43240
rect 31996 43228 32002 43240
rect 32125 43231 32183 43237
rect 32125 43228 32137 43231
rect 31996 43200 32137 43228
rect 31996 43188 32002 43200
rect 32125 43197 32137 43200
rect 32171 43197 32183 43231
rect 32416 43228 32444 43256
rect 35250 43228 35256 43240
rect 32416 43200 35256 43228
rect 32125 43191 32183 43197
rect 35250 43188 35256 43200
rect 35308 43228 35314 43240
rect 35989 43231 36047 43237
rect 35989 43228 36001 43231
rect 35308 43200 36001 43228
rect 35308 43188 35314 43200
rect 35989 43197 36001 43200
rect 36035 43228 36047 43231
rect 36078 43228 36084 43240
rect 36035 43200 36084 43228
rect 36035 43197 36047 43200
rect 35989 43191 36047 43197
rect 36078 43188 36084 43200
rect 36136 43188 36142 43240
rect 35342 43160 35348 43172
rect 20404 43132 22094 43160
rect 24228 43132 24440 43160
rect 20404 43120 20410 43132
rect 21082 43092 21088 43104
rect 19668 43064 19932 43092
rect 21043 43064 21088 43092
rect 19668 43052 19674 43064
rect 21082 43052 21088 43064
rect 21140 43052 21146 43104
rect 21358 43052 21364 43104
rect 21416 43092 21422 43104
rect 24228 43092 24256 43132
rect 21416 43064 24256 43092
rect 24412 43092 24440 43132
rect 26252 43132 26464 43160
rect 26252 43092 26280 43132
rect 24412 43064 26280 43092
rect 26436 43092 26464 43132
rect 29104 43132 35348 43160
rect 29104 43092 29132 43132
rect 35342 43120 35348 43132
rect 35400 43120 35406 43172
rect 48038 43160 48044 43172
rect 47999 43132 48044 43160
rect 48038 43120 48044 43132
rect 48096 43120 48102 43172
rect 26436 43064 29132 43092
rect 21416 43052 21422 43064
rect 31294 43052 31300 43104
rect 31352 43092 31358 43104
rect 31481 43095 31539 43101
rect 31481 43092 31493 43095
rect 31352 43064 31493 43092
rect 31352 43052 31358 43064
rect 31481 43061 31493 43064
rect 31527 43061 31539 43095
rect 46934 43092 46940 43104
rect 46895 43064 46940 43092
rect 31481 43055 31539 43061
rect 46934 43052 46940 43064
rect 46992 43052 46998 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 4706 42848 4712 42900
rect 4764 42888 4770 42900
rect 5537 42891 5595 42897
rect 5537 42888 5549 42891
rect 4764 42860 5549 42888
rect 4764 42848 4770 42860
rect 5537 42857 5549 42860
rect 5583 42857 5595 42891
rect 5537 42851 5595 42857
rect 7006 42848 7012 42900
rect 7064 42888 7070 42900
rect 7101 42891 7159 42897
rect 7101 42888 7113 42891
rect 7064 42860 7113 42888
rect 7064 42848 7070 42860
rect 7101 42857 7113 42860
rect 7147 42857 7159 42891
rect 7101 42851 7159 42857
rect 8297 42891 8355 42897
rect 8297 42857 8309 42891
rect 8343 42888 8355 42891
rect 8938 42888 8944 42900
rect 8343 42860 8944 42888
rect 8343 42857 8355 42860
rect 8297 42851 8355 42857
rect 8938 42848 8944 42860
rect 8996 42848 9002 42900
rect 10502 42888 10508 42900
rect 10463 42860 10508 42888
rect 10502 42848 10508 42860
rect 10560 42848 10566 42900
rect 11974 42888 11980 42900
rect 11935 42860 11980 42888
rect 11974 42848 11980 42860
rect 12032 42848 12038 42900
rect 20622 42888 20628 42900
rect 17880 42860 20628 42888
rect 2314 42780 2320 42832
rect 2372 42820 2378 42832
rect 2372 42792 3096 42820
rect 2372 42780 2378 42792
rect 2682 42752 2688 42764
rect 2643 42724 2688 42752
rect 2682 42712 2688 42724
rect 2740 42712 2746 42764
rect 2501 42687 2559 42693
rect 2501 42653 2513 42687
rect 2547 42684 2559 42687
rect 2590 42684 2596 42696
rect 2547 42656 2596 42684
rect 2547 42653 2559 42656
rect 2501 42647 2559 42653
rect 2590 42644 2596 42656
rect 2648 42644 2654 42696
rect 3068 42693 3096 42792
rect 4246 42780 4252 42832
rect 4304 42820 4310 42832
rect 4614 42820 4620 42832
rect 4304 42792 4620 42820
rect 4304 42780 4310 42792
rect 4614 42780 4620 42792
rect 4672 42820 4678 42832
rect 9214 42820 9220 42832
rect 4672 42792 9220 42820
rect 4672 42780 4678 42792
rect 9214 42780 9220 42792
rect 9272 42780 9278 42832
rect 4341 42755 4399 42761
rect 4341 42721 4353 42755
rect 4387 42752 4399 42755
rect 4522 42752 4528 42764
rect 4387 42724 4528 42752
rect 4387 42721 4399 42724
rect 4341 42715 4399 42721
rect 4522 42712 4528 42724
rect 4580 42752 4586 42764
rect 5169 42755 5227 42761
rect 4580 42724 5028 42752
rect 4580 42712 4586 42724
rect 2768 42687 2826 42693
rect 3053 42687 3111 42693
rect 2768 42647 2780 42687
rect 2814 42674 2826 42687
rect 2869 42681 2927 42687
rect 1857 42619 1915 42625
rect 2774 42622 2780 42647
rect 2832 42622 2838 42674
rect 2869 42647 2881 42681
rect 2915 42647 2927 42681
rect 3053 42653 3065 42687
rect 3099 42684 3111 42687
rect 4706 42684 4712 42696
rect 3099 42656 4712 42684
rect 3099 42653 3111 42656
rect 3053 42647 3111 42653
rect 2869 42641 2927 42647
rect 4706 42644 4712 42656
rect 4764 42644 4770 42696
rect 4801 42687 4859 42693
rect 4801 42653 4813 42687
rect 4847 42684 4859 42687
rect 4890 42684 4896 42696
rect 4847 42656 4896 42684
rect 4847 42653 4859 42656
rect 4801 42647 4859 42653
rect 4890 42644 4896 42656
rect 4948 42644 4954 42696
rect 5000 42693 5028 42724
rect 5169 42721 5181 42755
rect 5215 42752 5227 42755
rect 6730 42752 6736 42764
rect 5215 42724 6736 42752
rect 5215 42721 5227 42724
rect 5169 42715 5227 42721
rect 6730 42712 6736 42724
rect 6788 42712 6794 42764
rect 8110 42752 8116 42764
rect 6932 42724 8116 42752
rect 4985 42687 5043 42693
rect 4985 42653 4997 42687
rect 5031 42653 5043 42687
rect 4985 42647 5043 42653
rect 5077 42687 5135 42693
rect 5077 42653 5089 42687
rect 5123 42653 5135 42687
rect 5077 42647 5135 42653
rect 5353 42687 5411 42693
rect 5353 42653 5365 42687
rect 5399 42684 5411 42687
rect 5810 42684 5816 42696
rect 5399 42656 5816 42684
rect 5399 42653 5411 42656
rect 5353 42647 5411 42653
rect 1857 42585 1869 42619
rect 1903 42616 1915 42619
rect 1903 42588 2452 42616
rect 1903 42585 1915 42588
rect 1857 42579 1915 42585
rect 2314 42548 2320 42560
rect 2275 42520 2320 42548
rect 2314 42508 2320 42520
rect 2372 42508 2378 42560
rect 2424 42548 2452 42588
rect 2884 42548 2912 42641
rect 3234 42548 3240 42560
rect 2424 42520 3240 42548
rect 3234 42508 3240 42520
rect 3292 42508 3298 42560
rect 4908 42548 4936 42644
rect 5092 42616 5120 42647
rect 5810 42644 5816 42656
rect 5868 42644 5874 42696
rect 6362 42684 6368 42696
rect 6323 42656 6368 42684
rect 6362 42644 6368 42656
rect 6420 42644 6426 42696
rect 6546 42684 6552 42696
rect 6507 42656 6552 42684
rect 6546 42644 6552 42656
rect 6604 42644 6610 42696
rect 6932 42693 6960 42724
rect 8110 42712 8116 42724
rect 8168 42712 8174 42764
rect 17126 42712 17132 42764
rect 17184 42752 17190 42764
rect 17880 42761 17908 42860
rect 20622 42848 20628 42860
rect 20680 42848 20686 42900
rect 20990 42888 20996 42900
rect 20951 42860 20996 42888
rect 20990 42848 20996 42860
rect 21048 42848 21054 42900
rect 23290 42888 23296 42900
rect 23251 42860 23296 42888
rect 23290 42848 23296 42860
rect 23348 42848 23354 42900
rect 25133 42891 25191 42897
rect 25133 42857 25145 42891
rect 25179 42888 25191 42891
rect 25222 42888 25228 42900
rect 25179 42860 25228 42888
rect 25179 42857 25191 42860
rect 25133 42851 25191 42857
rect 25222 42848 25228 42860
rect 25280 42848 25286 42900
rect 29917 42891 29975 42897
rect 29917 42857 29929 42891
rect 29963 42888 29975 42891
rect 30098 42888 30104 42900
rect 29963 42860 30104 42888
rect 29963 42857 29975 42860
rect 29917 42851 29975 42857
rect 30098 42848 30104 42860
rect 30156 42848 30162 42900
rect 34054 42888 34060 42900
rect 33967 42860 34060 42888
rect 34054 42848 34060 42860
rect 34112 42888 34118 42900
rect 41506 42888 41512 42900
rect 34112 42860 41512 42888
rect 34112 42848 34118 42860
rect 41506 42848 41512 42860
rect 41564 42848 41570 42900
rect 36262 42820 36268 42832
rect 36223 42792 36268 42820
rect 36262 42780 36268 42792
rect 36320 42780 36326 42832
rect 17865 42755 17923 42761
rect 17865 42752 17877 42755
rect 17184 42724 17877 42752
rect 17184 42712 17190 42724
rect 17865 42721 17877 42724
rect 17911 42721 17923 42755
rect 17865 42715 17923 42721
rect 18325 42755 18383 42761
rect 18325 42721 18337 42755
rect 18371 42752 18383 42755
rect 19334 42752 19340 42764
rect 18371 42724 19340 42752
rect 18371 42721 18383 42724
rect 18325 42715 18383 42721
rect 19334 42712 19340 42724
rect 19392 42712 19398 42764
rect 19610 42752 19616 42764
rect 19571 42724 19616 42752
rect 19610 42712 19616 42724
rect 19668 42712 19674 42764
rect 21910 42752 21916 42764
rect 21871 42724 21916 42752
rect 21910 42712 21916 42724
rect 21968 42712 21974 42764
rect 24762 42752 24768 42764
rect 24723 42724 24768 42752
rect 24762 42712 24768 42724
rect 24820 42712 24826 42764
rect 6641 42687 6699 42693
rect 6641 42653 6653 42687
rect 6687 42653 6699 42687
rect 6641 42647 6699 42653
rect 6917 42687 6975 42693
rect 6917 42653 6929 42687
rect 6963 42653 6975 42687
rect 8202 42684 8208 42696
rect 6917 42647 6975 42653
rect 7760 42656 8208 42684
rect 6656 42616 6684 42647
rect 7098 42616 7104 42628
rect 5092 42588 7104 42616
rect 7098 42576 7104 42588
rect 7156 42576 7162 42628
rect 7760 42560 7788 42656
rect 8202 42644 8208 42656
rect 8260 42684 8266 42696
rect 9122 42684 9128 42696
rect 8260 42656 9128 42684
rect 8260 42644 8266 42656
rect 9122 42644 9128 42656
rect 9180 42684 9186 42696
rect 9401 42687 9459 42693
rect 9401 42684 9413 42687
rect 9180 42656 9413 42684
rect 9180 42644 9186 42656
rect 9401 42653 9413 42656
rect 9447 42653 9459 42687
rect 10502 42684 10508 42696
rect 10463 42656 10508 42684
rect 9401 42647 9459 42653
rect 10502 42644 10508 42656
rect 10560 42644 10566 42696
rect 17402 42644 17408 42696
rect 17460 42684 17466 42696
rect 17589 42687 17647 42693
rect 17589 42684 17601 42687
rect 17460 42656 17601 42684
rect 17460 42644 17466 42656
rect 17589 42653 17601 42656
rect 17635 42653 17647 42687
rect 17589 42647 17647 42653
rect 17773 42687 17831 42693
rect 17773 42653 17785 42687
rect 17819 42653 17831 42687
rect 17773 42647 17831 42653
rect 17957 42687 18015 42693
rect 17957 42653 17969 42687
rect 18003 42653 18015 42687
rect 17957 42647 18015 42653
rect 18141 42687 18199 42693
rect 18141 42653 18153 42687
rect 18187 42684 18199 42687
rect 18690 42684 18696 42696
rect 18187 42656 18696 42684
rect 18187 42653 18199 42656
rect 18141 42647 18199 42653
rect 6362 42548 6368 42560
rect 4908 42520 6368 42548
rect 6362 42508 6368 42520
rect 6420 42508 6426 42560
rect 7742 42548 7748 42560
rect 7703 42520 7748 42548
rect 7742 42508 7748 42520
rect 7800 42508 7806 42560
rect 9674 42548 9680 42560
rect 9635 42520 9680 42548
rect 9674 42508 9680 42520
rect 9732 42508 9738 42560
rect 17129 42551 17187 42557
rect 17129 42517 17141 42551
rect 17175 42548 17187 42551
rect 17788 42548 17816 42647
rect 17972 42616 18000 42647
rect 18690 42644 18696 42656
rect 18748 42644 18754 42696
rect 19880 42687 19938 42693
rect 19880 42653 19892 42687
rect 19926 42684 19938 42687
rect 21082 42684 21088 42696
rect 19926 42656 21088 42684
rect 19926 42653 19938 42656
rect 19880 42647 19938 42653
rect 21082 42644 21088 42656
rect 21140 42644 21146 42696
rect 22189 42687 22247 42693
rect 22189 42653 22201 42687
rect 22235 42684 22247 42687
rect 23842 42684 23848 42696
rect 22235 42656 23848 42684
rect 22235 42653 22247 42656
rect 22189 42647 22247 42653
rect 23842 42644 23848 42656
rect 23900 42684 23906 42696
rect 24397 42687 24455 42693
rect 24397 42684 24409 42687
rect 23900 42656 24409 42684
rect 23900 42644 23906 42656
rect 24397 42653 24409 42656
rect 24443 42653 24455 42687
rect 24397 42647 24455 42653
rect 24581 42687 24639 42693
rect 24581 42653 24593 42687
rect 24627 42653 24639 42687
rect 24581 42647 24639 42653
rect 24673 42687 24731 42693
rect 24673 42653 24685 42687
rect 24719 42653 24731 42687
rect 24673 42647 24731 42653
rect 24949 42687 25007 42693
rect 24949 42653 24961 42687
rect 24995 42684 25007 42687
rect 26326 42684 26332 42696
rect 24995 42656 26332 42684
rect 24995 42653 25007 42656
rect 24949 42647 25007 42653
rect 18322 42616 18328 42628
rect 17972 42588 18328 42616
rect 18322 42576 18328 42588
rect 18380 42576 18386 42628
rect 23382 42616 23388 42628
rect 23343 42588 23388 42616
rect 23382 42576 23388 42588
rect 23440 42576 23446 42628
rect 24210 42576 24216 42628
rect 24268 42616 24274 42628
rect 24596 42616 24624 42647
rect 24268 42588 24624 42616
rect 24268 42576 24274 42588
rect 18506 42548 18512 42560
rect 17175 42520 18512 42548
rect 17175 42517 17187 42520
rect 17129 42511 17187 42517
rect 18506 42508 18512 42520
rect 18564 42508 18570 42560
rect 23566 42508 23572 42560
rect 23624 42548 23630 42560
rect 24688 42548 24716 42647
rect 26326 42644 26332 42656
rect 26384 42644 26390 42696
rect 26786 42644 26792 42696
rect 26844 42684 26850 42696
rect 30561 42687 30619 42693
rect 30561 42684 30573 42687
rect 26844 42656 30573 42684
rect 26844 42644 26850 42656
rect 30561 42653 30573 42656
rect 30607 42653 30619 42687
rect 30561 42647 30619 42653
rect 30745 42687 30803 42693
rect 30745 42653 30757 42687
rect 30791 42684 30803 42687
rect 31110 42684 31116 42696
rect 30791 42656 31116 42684
rect 30791 42653 30803 42656
rect 30745 42647 30803 42653
rect 30576 42616 30604 42647
rect 31110 42644 31116 42656
rect 31168 42644 31174 42696
rect 32674 42684 32680 42696
rect 32587 42656 32680 42684
rect 32674 42644 32680 42656
rect 32732 42684 32738 42696
rect 34885 42687 34943 42693
rect 34885 42684 34897 42687
rect 32732 42656 34897 42684
rect 32732 42644 32738 42656
rect 34885 42653 34897 42656
rect 34931 42653 34943 42687
rect 47857 42687 47915 42693
rect 47857 42684 47869 42687
rect 34885 42647 34943 42653
rect 47320 42656 47869 42684
rect 31205 42619 31263 42625
rect 31205 42616 31217 42619
rect 30576 42588 31217 42616
rect 31205 42585 31217 42588
rect 31251 42585 31263 42619
rect 31205 42579 31263 42585
rect 32490 42576 32496 42628
rect 32548 42616 32554 42628
rect 32922 42619 32980 42625
rect 32922 42616 32934 42619
rect 32548 42588 32934 42616
rect 32548 42576 32554 42588
rect 32922 42585 32934 42588
rect 32968 42585 32980 42619
rect 32922 42579 32980 42585
rect 34790 42576 34796 42628
rect 34848 42616 34854 42628
rect 35130 42619 35188 42625
rect 35130 42616 35142 42619
rect 34848 42588 35142 42616
rect 34848 42576 34854 42588
rect 35130 42585 35142 42588
rect 35176 42585 35188 42619
rect 35130 42579 35188 42585
rect 47320 42560 47348 42656
rect 47857 42653 47869 42656
rect 47903 42653 47915 42687
rect 47857 42647 47915 42653
rect 23624 42520 24716 42548
rect 23624 42508 23630 42520
rect 30466 42508 30472 42560
rect 30524 42548 30530 42560
rect 30653 42551 30711 42557
rect 30653 42548 30665 42551
rect 30524 42520 30665 42548
rect 30524 42508 30530 42520
rect 30653 42517 30665 42520
rect 30699 42517 30711 42551
rect 31938 42548 31944 42560
rect 31899 42520 31944 42548
rect 30653 42511 30711 42517
rect 31938 42508 31944 42520
rect 31996 42508 32002 42560
rect 47302 42548 47308 42560
rect 47263 42520 47308 42548
rect 47302 42508 47308 42520
rect 47360 42508 47366 42560
rect 48038 42548 48044 42560
rect 47999 42520 48044 42548
rect 48038 42508 48044 42520
rect 48096 42508 48102 42560
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 4246 42344 4252 42356
rect 4207 42316 4252 42344
rect 4246 42304 4252 42316
rect 4304 42304 4310 42356
rect 4801 42347 4859 42353
rect 4801 42313 4813 42347
rect 4847 42344 4859 42347
rect 4982 42344 4988 42356
rect 4847 42316 4988 42344
rect 4847 42313 4859 42316
rect 4801 42307 4859 42313
rect 2314 42236 2320 42288
rect 2372 42276 2378 42288
rect 3430 42279 3488 42285
rect 3430 42276 3442 42279
rect 2372 42248 3442 42276
rect 2372 42236 2378 42248
rect 3430 42245 3442 42248
rect 3476 42245 3488 42279
rect 3430 42239 3488 42245
rect 1673 42211 1731 42217
rect 1673 42177 1685 42211
rect 1719 42208 1731 42211
rect 1946 42208 1952 42220
rect 1719 42180 1952 42208
rect 1719 42177 1731 42180
rect 1673 42171 1731 42177
rect 1946 42168 1952 42180
rect 2004 42168 2010 42220
rect 3697 42211 3755 42217
rect 3697 42177 3709 42211
rect 3743 42208 3755 42211
rect 4816 42208 4844 42307
rect 4982 42304 4988 42316
rect 5040 42304 5046 42356
rect 6914 42304 6920 42356
rect 6972 42344 6978 42356
rect 8297 42347 8355 42353
rect 8297 42344 8309 42347
rect 6972 42316 8309 42344
rect 6972 42304 6978 42316
rect 8297 42313 8309 42316
rect 8343 42344 8355 42347
rect 9950 42344 9956 42356
rect 8343 42316 9956 42344
rect 8343 42313 8355 42316
rect 8297 42307 8355 42313
rect 9950 42304 9956 42316
rect 10008 42304 10014 42356
rect 10134 42304 10140 42356
rect 10192 42344 10198 42356
rect 10229 42347 10287 42353
rect 10229 42344 10241 42347
rect 10192 42316 10241 42344
rect 10192 42304 10198 42316
rect 10229 42313 10241 42316
rect 10275 42344 10287 42347
rect 10502 42344 10508 42356
rect 10275 42316 10508 42344
rect 10275 42313 10287 42316
rect 10229 42307 10287 42313
rect 10502 42304 10508 42316
rect 10560 42344 10566 42356
rect 26786 42344 26792 42356
rect 10560 42316 26792 42344
rect 10560 42304 10566 42316
rect 26786 42304 26792 42316
rect 26844 42304 26850 42356
rect 46937 42347 46995 42353
rect 46937 42344 46949 42347
rect 26896 42316 46949 42344
rect 9122 42276 9128 42288
rect 9083 42248 9128 42276
rect 9122 42236 9128 42248
rect 9180 42236 9186 42288
rect 20070 42236 20076 42288
rect 20128 42276 20134 42288
rect 20257 42279 20315 42285
rect 20257 42276 20269 42279
rect 20128 42248 20269 42276
rect 20128 42236 20134 42248
rect 20257 42245 20269 42248
rect 20303 42276 20315 42279
rect 20530 42276 20536 42288
rect 20303 42248 20536 42276
rect 20303 42245 20315 42248
rect 20257 42239 20315 42245
rect 20530 42236 20536 42248
rect 20588 42236 20594 42288
rect 24121 42279 24179 42285
rect 24121 42276 24133 42279
rect 20640 42248 24133 42276
rect 3743 42180 4844 42208
rect 3743 42177 3755 42180
rect 3697 42171 3755 42177
rect 14458 42168 14464 42220
rect 14516 42208 14522 42220
rect 20640 42208 20668 42248
rect 24121 42245 24133 42248
rect 24167 42245 24179 42279
rect 26896 42276 26924 42316
rect 46937 42313 46949 42316
rect 46983 42313 46995 42347
rect 46937 42307 46995 42313
rect 32674 42276 32680 42288
rect 24121 42239 24179 42245
rect 26436 42248 26924 42276
rect 30208 42248 32680 42276
rect 26436 42208 26464 42248
rect 14516 42180 20668 42208
rect 22066 42180 26464 42208
rect 14516 42168 14522 42180
rect 12434 42100 12440 42152
rect 12492 42140 12498 42152
rect 22066 42140 22094 42180
rect 27982 42168 27988 42220
rect 28040 42208 28046 42220
rect 30208 42217 30236 42248
rect 32674 42236 32680 42248
rect 32732 42236 32738 42288
rect 30466 42217 30472 42220
rect 30193 42211 30251 42217
rect 30193 42208 30205 42211
rect 28040 42180 30205 42208
rect 28040 42168 28046 42180
rect 30193 42177 30205 42180
rect 30239 42177 30251 42211
rect 30460 42208 30472 42217
rect 30427 42180 30472 42208
rect 30193 42171 30251 42177
rect 30460 42171 30472 42180
rect 30466 42168 30472 42171
rect 30524 42168 30530 42220
rect 46952 42208 46980 42307
rect 47857 42211 47915 42217
rect 47857 42208 47869 42211
rect 46952 42180 47869 42208
rect 47857 42177 47869 42180
rect 47903 42177 47915 42211
rect 47857 42171 47915 42177
rect 12492 42112 22094 42140
rect 12492 42100 12498 42112
rect 2317 42075 2375 42081
rect 2317 42041 2329 42075
rect 2363 42072 2375 42075
rect 2590 42072 2596 42084
rect 2363 42044 2596 42072
rect 2363 42041 2375 42044
rect 2317 42035 2375 42041
rect 2590 42032 2596 42044
rect 2648 42032 2654 42084
rect 24121 42075 24179 42081
rect 24121 42041 24133 42075
rect 24167 42072 24179 42075
rect 24167 42044 24348 42072
rect 24167 42041 24179 42044
rect 24121 42035 24179 42041
rect 1486 42004 1492 42016
rect 1447 41976 1492 42004
rect 1486 41964 1492 41976
rect 1544 41964 1550 42016
rect 6457 42007 6515 42013
rect 6457 41973 6469 42007
rect 6503 42004 6515 42007
rect 6546 42004 6552 42016
rect 6503 41976 6552 42004
rect 6503 41973 6515 41976
rect 6457 41967 6515 41973
rect 6546 41964 6552 41976
rect 6604 41964 6610 42016
rect 24210 42004 24216 42016
rect 24171 41976 24216 42004
rect 24210 41964 24216 41976
rect 24268 41964 24274 42016
rect 24320 42004 24348 42044
rect 31128 42044 31754 42072
rect 31128 42004 31156 42044
rect 31570 42004 31576 42016
rect 24320 41976 31156 42004
rect 31531 41976 31576 42004
rect 31570 41964 31576 41976
rect 31628 41964 31634 42016
rect 31726 42004 31754 42044
rect 34698 42004 34704 42016
rect 31726 41976 34704 42004
rect 34698 41964 34704 41976
rect 34756 41964 34762 42016
rect 48038 42004 48044 42016
rect 47999 41976 48044 42004
rect 48038 41964 48044 41976
rect 48096 41964 48102 42016
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1946 41800 1952 41812
rect 1907 41772 1952 41800
rect 1946 41760 1952 41772
rect 2004 41760 2010 41812
rect 3881 41803 3939 41809
rect 3881 41769 3893 41803
rect 3927 41800 3939 41803
rect 4706 41800 4712 41812
rect 3927 41772 4712 41800
rect 3927 41769 3939 41772
rect 3881 41763 3939 41769
rect 4706 41760 4712 41772
rect 4764 41760 4770 41812
rect 12250 41760 12256 41812
rect 12308 41800 12314 41812
rect 47302 41800 47308 41812
rect 12308 41772 47308 41800
rect 12308 41760 12314 41772
rect 47302 41760 47308 41772
rect 47360 41760 47366 41812
rect 2774 41692 2780 41744
rect 2832 41732 2838 41744
rect 3237 41735 3295 41741
rect 3237 41732 3249 41735
rect 2832 41704 3249 41732
rect 2832 41692 2838 41704
rect 3237 41701 3249 41704
rect 3283 41732 3295 41735
rect 9674 41732 9680 41744
rect 3283 41704 9680 41732
rect 3283 41701 3295 41704
rect 3237 41695 3295 41701
rect 9674 41692 9680 41704
rect 9732 41732 9738 41744
rect 30561 41735 30619 41741
rect 30561 41732 30573 41735
rect 9732 41704 30573 41732
rect 9732 41692 9738 41704
rect 30561 41701 30573 41704
rect 30607 41701 30619 41735
rect 31110 41732 31116 41744
rect 31071 41704 31116 41732
rect 30561 41695 30619 41701
rect 30576 41664 30604 41695
rect 31110 41692 31116 41704
rect 31168 41692 31174 41744
rect 31573 41667 31631 41673
rect 31573 41664 31585 41667
rect 30576 41636 31585 41664
rect 31573 41633 31585 41636
rect 31619 41664 31631 41667
rect 31846 41664 31852 41676
rect 31619 41636 31852 41664
rect 31619 41633 31631 41636
rect 31573 41627 31631 41633
rect 31846 41624 31852 41636
rect 31904 41624 31910 41676
rect 2133 41599 2191 41605
rect 2133 41565 2145 41599
rect 2179 41596 2191 41599
rect 2590 41596 2596 41608
rect 2179 41568 2596 41596
rect 2179 41565 2191 41568
rect 2133 41559 2191 41565
rect 2590 41556 2596 41568
rect 2648 41596 2654 41608
rect 2685 41599 2743 41605
rect 2685 41596 2697 41599
rect 2648 41568 2697 41596
rect 2648 41556 2654 41568
rect 2685 41565 2697 41568
rect 2731 41565 2743 41599
rect 2685 41559 2743 41565
rect 2700 41528 2728 41559
rect 9214 41556 9220 41608
rect 9272 41596 9278 41608
rect 30742 41596 30748 41608
rect 9272 41568 30748 41596
rect 9272 41556 9278 41568
rect 30742 41556 30748 41568
rect 30800 41556 30806 41608
rect 31294 41596 31300 41608
rect 31255 41568 31300 41596
rect 31294 41556 31300 41568
rect 31352 41556 31358 41608
rect 31389 41599 31447 41605
rect 31389 41565 31401 41599
rect 31435 41565 31447 41599
rect 31662 41596 31668 41608
rect 31623 41568 31668 41596
rect 31389 41559 31447 41565
rect 30760 41528 30788 41556
rect 31404 41528 31432 41559
rect 31662 41556 31668 41568
rect 31720 41556 31726 41608
rect 47397 41599 47455 41605
rect 47397 41565 47409 41599
rect 47443 41596 47455 41599
rect 48038 41596 48044 41608
rect 47443 41568 48044 41596
rect 47443 41565 47455 41568
rect 47397 41559 47455 41565
rect 48038 41556 48044 41568
rect 48096 41556 48102 41608
rect 31938 41528 31944 41540
rect 2700 41500 12434 41528
rect 30760 41500 31944 41528
rect 12406 41460 12434 41500
rect 31938 41488 31944 41500
rect 31996 41488 32002 41540
rect 46290 41488 46296 41540
rect 46348 41528 46354 41540
rect 47857 41531 47915 41537
rect 47857 41528 47869 41531
rect 46348 41500 47869 41528
rect 46348 41488 46354 41500
rect 47857 41497 47869 41500
rect 47903 41497 47915 41531
rect 47857 41491 47915 41497
rect 24578 41460 24584 41472
rect 12406 41432 24584 41460
rect 24578 41420 24584 41432
rect 24636 41420 24642 41472
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 30742 41256 30748 41268
rect 30703 41228 30748 41256
rect 30742 41216 30748 41228
rect 30800 41216 30806 41268
rect 48038 41120 48044 41132
rect 47999 41092 48044 41120
rect 48038 41080 48044 41092
rect 48096 41080 48102 41132
rect 47026 40944 47032 40996
rect 47084 40984 47090 40996
rect 47857 40987 47915 40993
rect 47857 40984 47869 40987
rect 47084 40956 47869 40984
rect 47084 40944 47090 40956
rect 47857 40953 47869 40956
rect 47903 40953 47915 40987
rect 47857 40947 47915 40953
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 18598 40672 18604 40724
rect 18656 40712 18662 40724
rect 46934 40712 46940 40724
rect 18656 40684 46940 40712
rect 18656 40672 18662 40684
rect 46934 40672 46940 40684
rect 46992 40672 46998 40724
rect 47581 40715 47639 40721
rect 47581 40681 47593 40715
rect 47627 40712 47639 40715
rect 48038 40712 48044 40724
rect 47627 40684 48044 40712
rect 47627 40681 47639 40684
rect 47581 40675 47639 40681
rect 48038 40672 48044 40684
rect 48096 40672 48102 40724
rect 48038 40372 48044 40384
rect 47999 40344 48044 40372
rect 48038 40332 48044 40344
rect 48096 40332 48102 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 13817 40103 13875 40109
rect 13817 40069 13829 40103
rect 13863 40100 13875 40103
rect 15194 40100 15200 40112
rect 13863 40072 15200 40100
rect 13863 40069 13875 40072
rect 13817 40063 13875 40069
rect 15194 40060 15200 40072
rect 15252 40060 15258 40112
rect 48038 40100 48044 40112
rect 47999 40072 48044 40100
rect 48038 40060 48044 40072
rect 48096 40060 48102 40112
rect 11974 39992 11980 40044
rect 12032 40032 12038 40044
rect 13633 40035 13691 40041
rect 13633 40032 13645 40035
rect 12032 40004 13645 40032
rect 12032 39992 12038 40004
rect 13633 40001 13645 40004
rect 13679 40001 13691 40035
rect 13633 39995 13691 40001
rect 47949 39831 48007 39837
rect 47949 39797 47961 39831
rect 47995 39828 48007 39831
rect 48130 39828 48136 39840
rect 47995 39800 48136 39828
rect 47995 39797 48007 39800
rect 47949 39791 48007 39797
rect 48130 39788 48136 39800
rect 48188 39788 48194 39840
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 47397 39355 47455 39361
rect 47397 39321 47409 39355
rect 47443 39352 47455 39355
rect 48038 39352 48044 39364
rect 47443 39324 48044 39352
rect 47443 39321 47455 39324
rect 47397 39315 47455 39321
rect 48038 39312 48044 39324
rect 48096 39312 48102 39364
rect 45554 39244 45560 39296
rect 45612 39284 45618 39296
rect 47949 39287 48007 39293
rect 47949 39284 47961 39287
rect 45612 39256 47961 39284
rect 45612 39244 45618 39256
rect 47949 39253 47961 39256
rect 47995 39253 48007 39287
rect 47949 39247 48007 39253
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 47029 38947 47087 38953
rect 47029 38913 47041 38947
rect 47075 38944 47087 38947
rect 48038 38944 48044 38956
rect 47075 38916 48044 38944
rect 47075 38913 47087 38916
rect 47029 38907 47087 38913
rect 48038 38904 48044 38916
rect 48096 38904 48102 38956
rect 47762 38768 47768 38820
rect 47820 38808 47826 38820
rect 47857 38811 47915 38817
rect 47857 38808 47869 38811
rect 47820 38780 47869 38808
rect 47820 38768 47826 38780
rect 47857 38777 47869 38780
rect 47903 38777 47915 38811
rect 47857 38771 47915 38777
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 27982 38468 27988 38480
rect 27943 38440 27988 38468
rect 27982 38428 27988 38440
rect 28040 38428 28046 38480
rect 23382 38224 23388 38276
rect 23440 38264 23446 38276
rect 27801 38267 27859 38273
rect 27801 38264 27813 38267
rect 23440 38236 27813 38264
rect 23440 38224 23446 38236
rect 27801 38233 27813 38236
rect 27847 38233 27859 38267
rect 27801 38227 27859 38233
rect 47397 38267 47455 38273
rect 47397 38233 47409 38267
rect 47443 38264 47455 38267
rect 48038 38264 48044 38276
rect 47443 38236 48044 38264
rect 47443 38233 47455 38236
rect 47397 38227 47455 38233
rect 48038 38224 48044 38236
rect 48096 38224 48102 38276
rect 46566 38156 46572 38208
rect 46624 38196 46630 38208
rect 47949 38199 48007 38205
rect 47949 38196 47961 38199
rect 46624 38168 47961 38196
rect 46624 38156 46630 38168
rect 47949 38165 47961 38168
rect 47995 38165 48007 38199
rect 47949 38159 48007 38165
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 48038 37856 48044 37868
rect 47999 37828 48044 37856
rect 48038 37816 48044 37828
rect 48096 37816 48102 37868
rect 47854 37720 47860 37732
rect 47815 37692 47860 37720
rect 47854 37680 47860 37692
rect 47912 37680 47918 37732
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 47581 37451 47639 37457
rect 47581 37417 47593 37451
rect 47627 37448 47639 37451
rect 48038 37448 48044 37460
rect 47627 37420 48044 37448
rect 47627 37417 47639 37420
rect 47581 37411 47639 37417
rect 48038 37408 48044 37420
rect 48096 37408 48102 37460
rect 48038 37108 48044 37120
rect 47999 37080 48044 37108
rect 48038 37068 48044 37080
rect 48096 37068 48102 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 48038 36768 48044 36780
rect 47999 36740 48044 36768
rect 48038 36728 48044 36740
rect 48096 36728 48102 36780
rect 45830 36592 45836 36644
rect 45888 36632 45894 36644
rect 47857 36635 47915 36641
rect 47857 36632 47869 36635
rect 45888 36604 47869 36632
rect 45888 36592 45894 36604
rect 47857 36601 47869 36604
rect 47903 36601 47915 36635
rect 47857 36595 47915 36601
rect 11146 36524 11152 36576
rect 11204 36564 11210 36576
rect 24210 36564 24216 36576
rect 11204 36536 24216 36564
rect 11204 36524 11210 36536
rect 24210 36524 24216 36536
rect 24268 36524 24274 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 9950 36360 9956 36372
rect 9911 36332 9956 36360
rect 9950 36320 9956 36332
rect 10008 36320 10014 36372
rect 2133 36295 2191 36301
rect 2133 36261 2145 36295
rect 2179 36261 2191 36295
rect 2133 36255 2191 36261
rect 1673 36159 1731 36165
rect 1673 36125 1685 36159
rect 1719 36156 1731 36159
rect 2148 36156 2176 36255
rect 1719 36128 2176 36156
rect 2317 36159 2375 36165
rect 1719 36125 1731 36128
rect 1673 36119 1731 36125
rect 2317 36125 2329 36159
rect 2363 36156 2375 36159
rect 2869 36159 2927 36165
rect 2869 36156 2881 36159
rect 2363 36128 2881 36156
rect 2363 36125 2375 36128
rect 2317 36119 2375 36125
rect 2869 36125 2881 36128
rect 2915 36156 2927 36159
rect 11146 36156 11152 36168
rect 2915 36128 11152 36156
rect 2915 36125 2927 36128
rect 2869 36119 2927 36125
rect 11146 36116 11152 36128
rect 11204 36116 11210 36168
rect 10045 36091 10103 36097
rect 10045 36057 10057 36091
rect 10091 36088 10103 36091
rect 15194 36088 15200 36100
rect 10091 36060 15200 36088
rect 10091 36057 10103 36060
rect 10045 36051 10103 36057
rect 15194 36048 15200 36060
rect 15252 36048 15258 36100
rect 47397 36091 47455 36097
rect 47397 36057 47409 36091
rect 47443 36088 47455 36091
rect 48038 36088 48044 36100
rect 47443 36060 48044 36088
rect 47443 36057 47455 36060
rect 47397 36051 47455 36057
rect 48038 36048 48044 36060
rect 48096 36048 48102 36100
rect 1486 36020 1492 36032
rect 1447 35992 1492 36020
rect 1486 35980 1492 35992
rect 1544 35980 1550 36032
rect 47946 36020 47952 36032
rect 47907 35992 47952 36020
rect 47946 35980 47952 35992
rect 48004 35980 48010 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 47029 35683 47087 35689
rect 47029 35649 47041 35683
rect 47075 35680 47087 35683
rect 48038 35680 48044 35692
rect 47075 35652 48044 35680
rect 47075 35649 47087 35652
rect 47029 35643 47087 35649
rect 48038 35640 48044 35652
rect 48096 35640 48102 35692
rect 45922 35504 45928 35556
rect 45980 35544 45986 35556
rect 47857 35547 47915 35553
rect 47857 35544 47869 35547
rect 45980 35516 47869 35544
rect 45980 35504 45986 35516
rect 47857 35513 47869 35516
rect 47903 35513 47915 35547
rect 47857 35507 47915 35513
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 47397 35003 47455 35009
rect 47397 34969 47409 35003
rect 47443 35000 47455 35003
rect 48038 35000 48044 35012
rect 47443 34972 48044 35000
rect 47443 34969 47455 34972
rect 47397 34963 47455 34969
rect 48038 34960 48044 34972
rect 48096 34960 48102 35012
rect 47118 34892 47124 34944
rect 47176 34932 47182 34944
rect 47949 34935 48007 34941
rect 47949 34932 47961 34935
rect 47176 34904 47961 34932
rect 47176 34892 47182 34904
rect 47949 34901 47961 34904
rect 47995 34901 48007 34935
rect 47949 34895 48007 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 48038 34592 48044 34604
rect 47999 34564 48044 34592
rect 48038 34552 48044 34564
rect 48096 34552 48102 34604
rect 47578 34484 47584 34536
rect 47636 34524 47642 34536
rect 47857 34527 47915 34533
rect 47857 34524 47869 34527
rect 47636 34496 47869 34524
rect 47636 34484 47642 34496
rect 47857 34493 47869 34496
rect 47903 34493 47915 34527
rect 47857 34487 47915 34493
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 47581 34187 47639 34193
rect 47581 34153 47593 34187
rect 47627 34184 47639 34187
rect 48038 34184 48044 34196
rect 47627 34156 48044 34184
rect 47627 34153 47639 34156
rect 47581 34147 47639 34153
rect 48038 34144 48044 34156
rect 48096 34144 48102 34196
rect 48038 33844 48044 33856
rect 47999 33816 48044 33844
rect 48038 33804 48044 33816
rect 48096 33804 48102 33856
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 48038 33504 48044 33516
rect 47999 33476 48044 33504
rect 48038 33464 48044 33476
rect 48096 33464 48102 33516
rect 47394 33328 47400 33380
rect 47452 33368 47458 33380
rect 47857 33371 47915 33377
rect 47857 33368 47869 33371
rect 47452 33340 47869 33368
rect 47452 33328 47458 33340
rect 47857 33337 47869 33340
rect 47903 33337 47915 33371
rect 47857 33331 47915 33337
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 47397 32827 47455 32833
rect 47397 32793 47409 32827
rect 47443 32824 47455 32827
rect 48038 32824 48044 32836
rect 47443 32796 48044 32824
rect 47443 32793 47455 32796
rect 47397 32787 47455 32793
rect 48038 32784 48044 32796
rect 48096 32784 48102 32836
rect 47210 32716 47216 32768
rect 47268 32756 47274 32768
rect 47949 32759 48007 32765
rect 47949 32756 47961 32759
rect 47268 32728 47961 32756
rect 47268 32716 47274 32728
rect 47949 32725 47961 32728
rect 47995 32725 48007 32759
rect 47949 32719 48007 32725
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 23382 32484 23388 32496
rect 23343 32456 23388 32484
rect 23382 32444 23388 32456
rect 23440 32444 23446 32496
rect 19886 32376 19892 32428
rect 19944 32416 19950 32428
rect 23201 32419 23259 32425
rect 23201 32416 23213 32419
rect 19944 32388 23213 32416
rect 19944 32376 19950 32388
rect 23201 32385 23213 32388
rect 23247 32385 23259 32419
rect 23201 32379 23259 32385
rect 47029 32419 47087 32425
rect 47029 32385 47041 32419
rect 47075 32416 47087 32419
rect 48038 32416 48044 32428
rect 47075 32388 48044 32416
rect 47075 32385 47087 32388
rect 47029 32379 47087 32385
rect 48038 32376 48044 32388
rect 48096 32376 48102 32428
rect 46014 32240 46020 32292
rect 46072 32280 46078 32292
rect 47857 32283 47915 32289
rect 47857 32280 47869 32283
rect 46072 32252 47869 32280
rect 46072 32240 46078 32252
rect 47857 32249 47869 32252
rect 47903 32249 47915 32283
rect 47857 32243 47915 32249
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 15194 31900 15200 31952
rect 15252 31940 15258 31952
rect 15933 31943 15991 31949
rect 15933 31940 15945 31943
rect 15252 31912 15945 31940
rect 15252 31900 15258 31912
rect 15933 31909 15945 31912
rect 15979 31909 15991 31943
rect 15933 31903 15991 31909
rect 47857 31875 47915 31881
rect 47857 31841 47869 31875
rect 47903 31872 47915 31875
rect 48961 31875 49019 31881
rect 48961 31872 48973 31875
rect 47903 31844 48973 31872
rect 47903 31841 47915 31844
rect 47857 31835 47915 31841
rect 48961 31841 48973 31844
rect 49007 31841 49019 31875
rect 48961 31835 49019 31841
rect 16117 31807 16175 31813
rect 16117 31773 16129 31807
rect 16163 31804 16175 31807
rect 19886 31804 19892 31816
rect 16163 31776 19892 31804
rect 16163 31773 16175 31776
rect 16117 31767 16175 31773
rect 19886 31764 19892 31776
rect 19944 31764 19950 31816
rect 47397 31807 47455 31813
rect 47397 31773 47409 31807
rect 47443 31804 47455 31807
rect 48038 31804 48044 31816
rect 47443 31776 48044 31804
rect 47443 31773 47455 31776
rect 47397 31767 47455 31773
rect 48038 31764 48044 31776
rect 48096 31764 48102 31816
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 48038 31328 48044 31340
rect 47999 31300 48044 31328
rect 48038 31288 48044 31300
rect 48096 31288 48102 31340
rect 45646 31152 45652 31204
rect 45704 31192 45710 31204
rect 47857 31195 47915 31201
rect 47857 31192 47869 31195
rect 45704 31164 47869 31192
rect 45704 31152 45710 31164
rect 47857 31161 47869 31164
rect 47903 31161 47915 31195
rect 47857 31155 47915 31161
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 47581 30923 47639 30929
rect 47581 30889 47593 30923
rect 47627 30920 47639 30923
rect 48038 30920 48044 30932
rect 47627 30892 48044 30920
rect 47627 30889 47639 30892
rect 47581 30883 47639 30889
rect 48038 30880 48044 30892
rect 48096 30880 48102 30932
rect 2133 30855 2191 30861
rect 2133 30821 2145 30855
rect 2179 30821 2191 30855
rect 2133 30815 2191 30821
rect 1673 30719 1731 30725
rect 1673 30685 1685 30719
rect 1719 30716 1731 30719
rect 2148 30716 2176 30815
rect 1719 30688 2176 30716
rect 2317 30719 2375 30725
rect 1719 30685 1731 30688
rect 1673 30679 1731 30685
rect 2317 30685 2329 30719
rect 2363 30716 2375 30719
rect 2363 30688 2912 30716
rect 2363 30685 2375 30688
rect 2317 30679 2375 30685
rect 2884 30592 2912 30688
rect 1486 30580 1492 30592
rect 1447 30552 1492 30580
rect 1486 30540 1492 30552
rect 1544 30540 1550 30592
rect 2866 30580 2872 30592
rect 2827 30552 2872 30580
rect 2866 30540 2872 30552
rect 2924 30580 2930 30592
rect 17218 30580 17224 30592
rect 2924 30552 17224 30580
rect 2924 30540 2930 30552
rect 17218 30540 17224 30552
rect 17276 30540 17282 30592
rect 48038 30580 48044 30592
rect 47999 30552 48044 30580
rect 48038 30540 48044 30552
rect 48096 30540 48102 30592
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 48038 30240 48044 30252
rect 47999 30212 48044 30240
rect 48038 30200 48044 30212
rect 48096 30200 48102 30252
rect 47949 30039 48007 30045
rect 47949 30005 47961 30039
rect 47995 30036 48007 30039
rect 49053 30039 49111 30045
rect 49053 30036 49065 30039
rect 47995 30008 49065 30036
rect 47995 30005 48007 30008
rect 47949 29999 48007 30005
rect 49053 30005 49065 30008
rect 49099 30005 49111 30039
rect 49053 29999 49111 30005
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 47397 29563 47455 29569
rect 47397 29529 47409 29563
rect 47443 29560 47455 29563
rect 48038 29560 48044 29572
rect 47443 29532 48044 29560
rect 47443 29529 47455 29532
rect 47397 29523 47455 29529
rect 48038 29520 48044 29532
rect 48096 29520 48102 29572
rect 45738 29452 45744 29504
rect 45796 29492 45802 29504
rect 47949 29495 48007 29501
rect 47949 29492 47961 29495
rect 45796 29464 47961 29492
rect 45796 29452 45802 29464
rect 47949 29461 47961 29464
rect 47995 29461 48007 29495
rect 47949 29455 48007 29461
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 47029 29155 47087 29161
rect 47029 29121 47041 29155
rect 47075 29152 47087 29155
rect 48038 29152 48044 29164
rect 47075 29124 48044 29152
rect 47075 29121 47087 29124
rect 47029 29115 47087 29121
rect 48038 29112 48044 29124
rect 48096 29112 48102 29164
rect 46658 28976 46664 29028
rect 46716 29016 46722 29028
rect 47857 29019 47915 29025
rect 47857 29016 47869 29019
rect 46716 28988 47869 29016
rect 46716 28976 46722 28988
rect 47857 28985 47869 28988
rect 47903 28985 47915 29019
rect 47857 28979 47915 28985
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 47397 28475 47455 28481
rect 47397 28441 47409 28475
rect 47443 28472 47455 28475
rect 48038 28472 48044 28484
rect 47443 28444 48044 28472
rect 47443 28441 47455 28444
rect 47397 28435 47455 28441
rect 48038 28432 48044 28444
rect 48096 28432 48102 28484
rect 44634 28364 44640 28416
rect 44692 28404 44698 28416
rect 47949 28407 48007 28413
rect 47949 28404 47961 28407
rect 44692 28376 47961 28404
rect 44692 28364 44698 28376
rect 47949 28373 47961 28376
rect 47995 28373 48007 28407
rect 47949 28367 48007 28373
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 48041 28067 48099 28073
rect 48041 28033 48053 28067
rect 48087 28064 48099 28067
rect 48222 28064 48228 28076
rect 48087 28036 48228 28064
rect 48087 28033 48099 28036
rect 48041 28027 48099 28033
rect 48222 28024 48228 28036
rect 48280 28024 48286 28076
rect 47949 27863 48007 27869
rect 47949 27829 47961 27863
rect 47995 27860 48007 27863
rect 48314 27860 48320 27872
rect 47995 27832 48320 27860
rect 47995 27829 48007 27832
rect 47949 27823 48007 27829
rect 48314 27820 48320 27832
rect 48372 27820 48378 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 48133 27591 48191 27597
rect 48133 27557 48145 27591
rect 48179 27588 48191 27591
rect 48222 27588 48228 27600
rect 48179 27560 48228 27588
rect 48179 27557 48191 27560
rect 48133 27551 48191 27557
rect 48222 27548 48228 27560
rect 48280 27548 48286 27600
rect 47581 27319 47639 27325
rect 47581 27285 47593 27319
rect 47627 27316 47639 27319
rect 48038 27316 48044 27328
rect 47627 27288 48044 27316
rect 47627 27285 47639 27288
rect 47581 27279 47639 27285
rect 48038 27276 48044 27288
rect 48096 27276 48102 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 48038 26976 48044 26988
rect 47999 26948 48044 26976
rect 48038 26936 48044 26948
rect 48096 26936 48102 26988
rect 47302 26868 47308 26920
rect 47360 26908 47366 26920
rect 47762 26908 47768 26920
rect 47360 26880 47768 26908
rect 47360 26868 47366 26880
rect 47762 26868 47768 26880
rect 47820 26868 47826 26920
rect 47946 26868 47952 26920
rect 48004 26908 48010 26920
rect 48222 26908 48228 26920
rect 48004 26880 48228 26908
rect 48004 26868 48010 26880
rect 48222 26868 48228 26880
rect 48280 26868 48286 26920
rect 47026 26800 47032 26852
rect 47084 26840 47090 26852
rect 47857 26843 47915 26849
rect 47857 26840 47869 26843
rect 47084 26812 47869 26840
rect 47084 26800 47090 26812
rect 47857 26809 47869 26812
rect 47903 26809 47915 26843
rect 47857 26803 47915 26809
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 47946 26568 47952 26580
rect 47907 26540 47952 26568
rect 47946 26528 47952 26540
rect 48004 26528 48010 26580
rect 47397 26299 47455 26305
rect 47397 26265 47409 26299
rect 47443 26296 47455 26299
rect 48038 26296 48044 26308
rect 47443 26268 48044 26296
rect 47443 26265 47455 26268
rect 47397 26259 47455 26265
rect 48038 26256 48044 26268
rect 48096 26256 48102 26308
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 47029 25891 47087 25897
rect 47029 25857 47041 25891
rect 47075 25888 47087 25891
rect 48038 25888 48044 25900
rect 47075 25860 48044 25888
rect 47075 25857 47087 25860
rect 47029 25851 47087 25857
rect 48038 25848 48044 25860
rect 48096 25848 48102 25900
rect 47670 25712 47676 25764
rect 47728 25752 47734 25764
rect 47857 25755 47915 25761
rect 47857 25752 47869 25755
rect 47728 25724 47869 25752
rect 47728 25712 47734 25724
rect 47857 25721 47869 25724
rect 47903 25721 47915 25755
rect 47857 25715 47915 25721
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 19978 25344 19984 25356
rect 19939 25316 19984 25344
rect 19978 25304 19984 25316
rect 20036 25304 20042 25356
rect 1670 25276 1676 25288
rect 1631 25248 1676 25276
rect 1670 25236 1676 25248
rect 1728 25236 1734 25288
rect 21637 25211 21695 25217
rect 21637 25177 21649 25211
rect 21683 25177 21695 25211
rect 21637 25171 21695 25177
rect 47397 25211 47455 25217
rect 47397 25177 47409 25211
rect 47443 25208 47455 25211
rect 48038 25208 48044 25220
rect 47443 25180 48044 25208
rect 47443 25177 47455 25180
rect 47397 25171 47455 25177
rect 1486 25140 1492 25152
rect 1447 25112 1492 25140
rect 1486 25100 1492 25112
rect 1544 25100 1550 25152
rect 21652 25140 21680 25171
rect 48038 25168 48044 25180
rect 48096 25168 48102 25220
rect 22189 25143 22247 25149
rect 22189 25140 22201 25143
rect 21652 25112 22201 25140
rect 22189 25109 22201 25112
rect 22235 25140 22247 25143
rect 28534 25140 28540 25152
rect 22235 25112 28540 25140
rect 22235 25109 22247 25112
rect 22189 25103 22247 25109
rect 28534 25100 28540 25112
rect 28592 25100 28598 25152
rect 47486 25100 47492 25152
rect 47544 25140 47550 25152
rect 47949 25143 48007 25149
rect 47949 25140 47961 25143
rect 47544 25112 47961 25140
rect 47544 25100 47550 25112
rect 47949 25109 47961 25112
rect 47995 25109 48007 25143
rect 47949 25103 48007 25109
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 1670 24896 1676 24948
rect 1728 24936 1734 24948
rect 1949 24939 2007 24945
rect 1949 24936 1961 24939
rect 1728 24908 1961 24936
rect 1728 24896 1734 24908
rect 1949 24905 1961 24908
rect 1995 24905 2007 24939
rect 1949 24899 2007 24905
rect 2133 24803 2191 24809
rect 2133 24769 2145 24803
rect 2179 24800 2191 24803
rect 2682 24800 2688 24812
rect 2179 24772 2688 24800
rect 2179 24769 2191 24772
rect 2133 24763 2191 24769
rect 2682 24760 2688 24772
rect 2740 24800 2746 24812
rect 8294 24800 8300 24812
rect 2740 24772 8300 24800
rect 2740 24760 2746 24772
rect 8294 24760 8300 24772
rect 8352 24760 8358 24812
rect 47029 24803 47087 24809
rect 47029 24769 47041 24803
rect 47075 24800 47087 24803
rect 48038 24800 48044 24812
rect 47075 24772 48044 24800
rect 47075 24769 47087 24772
rect 47029 24763 47087 24769
rect 48038 24760 48044 24772
rect 48096 24760 48102 24812
rect 47854 24664 47860 24676
rect 47815 24636 47860 24664
rect 47854 24624 47860 24636
rect 47912 24624 47918 24676
rect 2682 24596 2688 24608
rect 2643 24568 2688 24596
rect 2682 24556 2688 24568
rect 2740 24556 2746 24608
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 47397 24123 47455 24129
rect 47397 24089 47409 24123
rect 47443 24120 47455 24123
rect 48038 24120 48044 24132
rect 47443 24092 48044 24120
rect 47443 24089 47455 24092
rect 47397 24083 47455 24089
rect 48038 24080 48044 24092
rect 48096 24080 48102 24132
rect 45370 24012 45376 24064
rect 45428 24052 45434 24064
rect 47949 24055 48007 24061
rect 47949 24052 47961 24055
rect 45428 24024 47961 24052
rect 45428 24012 45434 24024
rect 47949 24021 47961 24024
rect 47995 24021 48007 24055
rect 47949 24015 48007 24021
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 47397 23035 47455 23041
rect 47397 23001 47409 23035
rect 47443 23032 47455 23035
rect 48038 23032 48044 23044
rect 47443 23004 48044 23032
rect 47443 23001 47455 23004
rect 47397 22995 47455 23001
rect 48038 22992 48044 23004
rect 48096 22992 48102 23044
rect 44266 22924 44272 22976
rect 44324 22964 44330 22976
rect 47949 22967 48007 22973
rect 47949 22964 47961 22967
rect 44324 22936 47961 22964
rect 44324 22924 44330 22936
rect 47949 22933 47961 22936
rect 47995 22933 48007 22967
rect 47949 22927 48007 22933
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 47029 22627 47087 22633
rect 47029 22593 47041 22627
rect 47075 22624 47087 22627
rect 48038 22624 48044 22636
rect 47075 22596 48044 22624
rect 47075 22593 47087 22596
rect 47029 22587 47087 22593
rect 48038 22584 48044 22596
rect 48096 22584 48102 22636
rect 47762 22448 47768 22500
rect 47820 22488 47826 22500
rect 47857 22491 47915 22497
rect 47857 22488 47869 22491
rect 47820 22460 47869 22488
rect 47820 22448 47826 22460
rect 47857 22457 47869 22460
rect 47903 22457 47915 22491
rect 47857 22451 47915 22457
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 48222 22108 48228 22160
rect 48280 22148 48286 22160
rect 48406 22148 48412 22160
rect 48280 22120 48412 22148
rect 48280 22108 48286 22120
rect 48406 22108 48412 22120
rect 48464 22108 48470 22160
rect 48038 22040 48044 22092
rect 48096 22080 48102 22092
rect 48096 22052 48268 22080
rect 48096 22040 48102 22052
rect 48240 22024 48268 22052
rect 47397 22015 47455 22021
rect 47397 21981 47409 22015
rect 47443 22012 47455 22015
rect 47946 22012 47952 22024
rect 47443 21984 47952 22012
rect 47443 21981 47455 21984
rect 47397 21975 47455 21981
rect 47946 21972 47952 21984
rect 48004 21972 48010 22024
rect 48222 21972 48228 22024
rect 48280 21972 48286 22024
rect 46845 21947 46903 21953
rect 46845 21913 46857 21947
rect 46891 21944 46903 21947
rect 48038 21944 48044 21956
rect 46891 21916 48044 21944
rect 46891 21913 46903 21916
rect 46845 21907 46903 21913
rect 48038 21904 48044 21916
rect 48096 21904 48102 21956
rect 45462 21836 45468 21888
rect 45520 21876 45526 21888
rect 47949 21879 48007 21885
rect 47949 21876 47961 21879
rect 45520 21848 47961 21876
rect 45520 21836 45526 21848
rect 47949 21845 47961 21848
rect 47995 21845 48007 21879
rect 47949 21839 48007 21845
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 48222 21632 48228 21684
rect 48280 21632 48286 21684
rect 48038 21536 48044 21548
rect 47999 21508 48044 21536
rect 48038 21496 48044 21508
rect 48096 21496 48102 21548
rect 47946 21428 47952 21480
rect 48004 21468 48010 21480
rect 48240 21468 48268 21632
rect 48004 21440 48268 21468
rect 48004 21428 48010 21440
rect 47029 21403 47087 21409
rect 47029 21369 47041 21403
rect 47075 21400 47087 21403
rect 48130 21400 48136 21412
rect 47075 21372 48136 21400
rect 47075 21369 47087 21372
rect 47029 21363 47087 21369
rect 48130 21360 48136 21372
rect 48188 21360 48194 21412
rect 45830 21292 45836 21344
rect 45888 21332 45894 21344
rect 46106 21332 46112 21344
rect 45888 21304 46112 21332
rect 45888 21292 45894 21304
rect 46106 21292 46112 21304
rect 46164 21292 46170 21344
rect 46750 21292 46756 21344
rect 46808 21332 46814 21344
rect 47949 21335 48007 21341
rect 47949 21332 47961 21335
rect 46808 21304 47961 21332
rect 46808 21292 46814 21304
rect 47949 21301 47961 21304
rect 47995 21301 48007 21335
rect 47949 21295 48007 21301
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 45922 21020 45928 21072
rect 45980 21060 45986 21072
rect 47305 21063 47363 21069
rect 47305 21060 47317 21063
rect 45980 21032 47317 21060
rect 45980 21020 45986 21032
rect 47305 21029 47317 21032
rect 47351 21029 47363 21063
rect 47305 21023 47363 21029
rect 46293 20927 46351 20933
rect 46293 20893 46305 20927
rect 46339 20924 46351 20927
rect 47486 20924 47492 20936
rect 46339 20896 47492 20924
rect 46339 20893 46351 20896
rect 46293 20887 46351 20893
rect 47486 20884 47492 20896
rect 47544 20884 47550 20936
rect 48130 20924 48136 20936
rect 48091 20896 48136 20924
rect 48130 20884 48136 20896
rect 48188 20884 48194 20936
rect 46474 20816 46480 20868
rect 46532 20856 46538 20868
rect 46532 20828 47992 20856
rect 46532 20816 46538 20828
rect 46842 20788 46848 20800
rect 46803 20760 46848 20788
rect 46842 20748 46848 20760
rect 46900 20748 46906 20800
rect 47964 20797 47992 20828
rect 47949 20791 48007 20797
rect 47949 20757 47961 20791
rect 47995 20757 48007 20791
rect 47949 20751 48007 20757
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 1210 20544 1216 20596
rect 1268 20584 1274 20596
rect 2590 20584 2596 20596
rect 1268 20556 2596 20584
rect 1268 20544 1274 20556
rect 2590 20544 2596 20556
rect 2648 20544 2654 20596
rect 46290 20544 46296 20596
rect 46348 20584 46354 20596
rect 46385 20587 46443 20593
rect 46385 20584 46397 20587
rect 46348 20556 46397 20584
rect 46348 20544 46354 20556
rect 46385 20553 46397 20556
rect 46431 20553 46443 20587
rect 46385 20547 46443 20553
rect 47029 20587 47087 20593
rect 47029 20553 47041 20587
rect 47075 20584 47087 20587
rect 47946 20584 47952 20596
rect 47075 20556 47952 20584
rect 47075 20553 47087 20556
rect 47029 20547 47087 20553
rect 47946 20544 47952 20556
rect 48004 20584 48010 20596
rect 48222 20584 48228 20596
rect 48004 20556 48228 20584
rect 48004 20544 48010 20556
rect 48222 20544 48228 20556
rect 48280 20544 48286 20596
rect 46842 20408 46848 20460
rect 46900 20448 46906 20460
rect 48133 20451 48191 20457
rect 48133 20448 48145 20451
rect 46900 20420 48145 20448
rect 46900 20408 46906 20420
rect 48133 20417 48145 20420
rect 48179 20448 48191 20451
rect 48222 20448 48228 20460
rect 48179 20420 48228 20448
rect 48179 20417 48191 20420
rect 48133 20411 48191 20417
rect 48222 20408 48228 20420
rect 48280 20408 48286 20460
rect 47578 20204 47584 20256
rect 47636 20244 47642 20256
rect 47949 20247 48007 20253
rect 47949 20244 47961 20247
rect 47636 20216 47961 20244
rect 47636 20204 47642 20216
rect 47949 20213 47961 20216
rect 47995 20213 48007 20247
rect 47949 20207 48007 20213
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 40678 19932 40684 19984
rect 40736 19972 40742 19984
rect 40736 19944 41414 19972
rect 40736 19932 40742 19944
rect 41386 19904 41414 19944
rect 46937 19907 46995 19913
rect 46937 19904 46949 19907
rect 41386 19876 46949 19904
rect 46937 19873 46949 19876
rect 46983 19873 46995 19907
rect 46937 19867 46995 19873
rect 47762 19864 47768 19916
rect 47820 19904 47826 19916
rect 47857 19907 47915 19913
rect 47857 19904 47869 19907
rect 47820 19876 47869 19904
rect 47820 19864 47826 19876
rect 47857 19873 47869 19876
rect 47903 19873 47915 19907
rect 47857 19867 47915 19873
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19836 1731 19839
rect 1946 19836 1952 19848
rect 1719 19808 1952 19836
rect 1719 19805 1731 19808
rect 1673 19799 1731 19805
rect 1946 19796 1952 19808
rect 2004 19796 2010 19848
rect 45741 19839 45799 19845
rect 45741 19805 45753 19839
rect 45787 19805 45799 19839
rect 45922 19836 45928 19848
rect 45883 19808 45928 19836
rect 45741 19799 45799 19805
rect 44818 19728 44824 19780
rect 44876 19768 44882 19780
rect 45281 19771 45339 19777
rect 45281 19768 45293 19771
rect 44876 19740 45293 19768
rect 44876 19728 44882 19740
rect 45281 19737 45293 19740
rect 45327 19737 45339 19771
rect 45756 19768 45784 19799
rect 45922 19796 45928 19808
rect 45980 19796 45986 19848
rect 46290 19836 46296 19848
rect 46251 19808 46296 19836
rect 46290 19796 46296 19808
rect 46348 19796 46354 19848
rect 46382 19796 46388 19848
rect 46440 19836 46446 19848
rect 46440 19808 46485 19836
rect 46440 19796 46446 19808
rect 46842 19796 46848 19848
rect 46900 19836 46906 19848
rect 47397 19839 47455 19845
rect 47397 19836 47409 19839
rect 46900 19808 47409 19836
rect 46900 19796 46906 19808
rect 47397 19805 47409 19808
rect 47443 19805 47455 19839
rect 47578 19836 47584 19848
rect 47539 19808 47584 19836
rect 47397 19799 47455 19805
rect 47578 19796 47584 19808
rect 47636 19796 47642 19848
rect 47946 19836 47952 19848
rect 47907 19808 47952 19836
rect 47946 19796 47952 19808
rect 48004 19796 48010 19848
rect 46198 19768 46204 19780
rect 45756 19740 46204 19768
rect 45281 19731 45339 19737
rect 46198 19728 46204 19740
rect 46256 19728 46262 19780
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 2685 19499 2743 19505
rect 2685 19465 2697 19499
rect 2731 19496 2743 19499
rect 6546 19496 6552 19508
rect 2731 19468 6552 19496
rect 2731 19465 2743 19468
rect 2685 19459 2743 19465
rect 2133 19363 2191 19369
rect 2133 19329 2145 19363
rect 2179 19360 2191 19363
rect 2700 19360 2728 19459
rect 6546 19456 6552 19468
rect 6604 19456 6610 19508
rect 14550 19388 14556 19440
rect 14608 19428 14614 19440
rect 40678 19428 40684 19440
rect 14608 19400 40684 19428
rect 14608 19388 14614 19400
rect 40678 19388 40684 19400
rect 40736 19388 40742 19440
rect 46382 19388 46388 19440
rect 46440 19428 46446 19440
rect 46440 19400 46796 19428
rect 46440 19388 46446 19400
rect 2179 19332 2728 19360
rect 2179 19329 2191 19332
rect 2133 19323 2191 19329
rect 1118 19252 1124 19304
rect 1176 19292 1182 19304
rect 2148 19292 2176 19323
rect 39298 19320 39304 19372
rect 39356 19360 39362 19372
rect 45833 19363 45891 19369
rect 45833 19360 45845 19363
rect 39356 19332 45845 19360
rect 39356 19320 39362 19332
rect 45833 19329 45845 19332
rect 45879 19329 45891 19363
rect 45833 19323 45891 19329
rect 46198 19320 46204 19372
rect 46256 19360 46262 19372
rect 46293 19363 46351 19369
rect 46293 19360 46305 19363
rect 46256 19332 46305 19360
rect 46256 19320 46262 19332
rect 46293 19329 46305 19332
rect 46339 19329 46351 19363
rect 46474 19360 46480 19372
rect 46435 19332 46480 19360
rect 46293 19323 46351 19329
rect 46474 19320 46480 19332
rect 46532 19320 46538 19372
rect 46768 19301 46796 19400
rect 46845 19363 46903 19369
rect 46845 19329 46857 19363
rect 46891 19360 46903 19363
rect 46934 19360 46940 19372
rect 46891 19332 46940 19360
rect 46891 19329 46903 19332
rect 46845 19323 46903 19329
rect 1176 19264 2176 19292
rect 46753 19295 46811 19301
rect 1176 19252 1182 19264
rect 46753 19261 46765 19295
rect 46799 19261 46811 19295
rect 46753 19255 46811 19261
rect 45373 19227 45431 19233
rect 45373 19193 45385 19227
rect 45419 19224 45431 19227
rect 46860 19224 46888 19323
rect 46934 19320 46940 19332
rect 46992 19320 46998 19372
rect 48038 19360 48044 19372
rect 47044 19332 48044 19360
rect 45419 19196 46888 19224
rect 45419 19193 45431 19196
rect 45373 19187 45431 19193
rect 44821 19159 44879 19165
rect 44821 19125 44833 19159
rect 44867 19156 44879 19159
rect 47044 19156 47072 19332
rect 48038 19320 48044 19332
rect 48096 19360 48102 19372
rect 48133 19363 48191 19369
rect 48133 19360 48145 19363
rect 48096 19332 48145 19360
rect 48096 19320 48102 19332
rect 48133 19329 48145 19332
rect 48179 19329 48191 19363
rect 48133 19323 48191 19329
rect 47394 19184 47400 19236
rect 47452 19224 47458 19236
rect 48130 19224 48136 19236
rect 47452 19196 48136 19224
rect 47452 19184 47458 19196
rect 48130 19184 48136 19196
rect 48188 19184 48194 19236
rect 44867 19128 47072 19156
rect 44867 19125 44879 19128
rect 44821 19119 44879 19125
rect 47578 19116 47584 19168
rect 47636 19156 47642 19168
rect 47949 19159 48007 19165
rect 47949 19156 47961 19159
rect 47636 19128 47961 19156
rect 47636 19116 47642 19128
rect 47949 19125 47961 19128
rect 47995 19125 48007 19159
rect 47949 19119 48007 19125
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 47118 18912 47124 18964
rect 47176 18952 47182 18964
rect 47394 18952 47400 18964
rect 47176 18924 47400 18952
rect 47176 18912 47182 18924
rect 47394 18912 47400 18924
rect 47452 18912 47458 18964
rect 45833 18887 45891 18893
rect 45833 18853 45845 18887
rect 45879 18884 45891 18887
rect 47210 18884 47216 18896
rect 45879 18856 47216 18884
rect 45879 18853 45891 18856
rect 45833 18847 45891 18853
rect 47210 18844 47216 18856
rect 47268 18884 47274 18896
rect 47268 18856 47992 18884
rect 47268 18844 47274 18856
rect 45922 18776 45928 18828
rect 45980 18816 45986 18828
rect 46842 18816 46848 18828
rect 45980 18788 46848 18816
rect 45980 18776 45986 18788
rect 46842 18776 46848 18788
rect 46900 18816 46906 18828
rect 47397 18819 47455 18825
rect 47397 18816 47409 18819
rect 46900 18788 47409 18816
rect 46900 18776 46906 18788
rect 47397 18785 47409 18788
rect 47443 18785 47455 18819
rect 47397 18779 47455 18785
rect 47762 18776 47768 18828
rect 47820 18816 47826 18828
rect 47857 18819 47915 18825
rect 47857 18816 47869 18819
rect 47820 18788 47869 18816
rect 47820 18776 47826 18788
rect 47857 18785 47869 18788
rect 47903 18785 47915 18819
rect 47857 18779 47915 18785
rect 45281 18751 45339 18757
rect 45281 18717 45293 18751
rect 45327 18748 45339 18751
rect 46290 18748 46296 18760
rect 45327 18720 46296 18748
rect 45327 18717 45339 18720
rect 45281 18711 45339 18717
rect 46290 18708 46296 18720
rect 46348 18708 46354 18760
rect 47578 18748 47584 18760
rect 47539 18720 47584 18748
rect 47578 18708 47584 18720
rect 47636 18708 47642 18760
rect 47964 18757 47992 18856
rect 47949 18751 48007 18757
rect 47949 18717 47961 18751
rect 47995 18717 48007 18751
rect 47949 18711 48007 18717
rect 46474 18612 46480 18624
rect 46435 18584 46480 18612
rect 46474 18572 46480 18584
rect 46532 18572 46538 18624
rect 47026 18612 47032 18624
rect 46987 18584 47032 18612
rect 47026 18572 47032 18584
rect 47084 18572 47090 18624
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 16114 18368 16120 18420
rect 16172 18408 16178 18420
rect 47026 18408 47032 18420
rect 16172 18380 47032 18408
rect 16172 18368 16178 18380
rect 47026 18368 47032 18380
rect 47084 18368 47090 18420
rect 44821 18343 44879 18349
rect 44821 18309 44833 18343
rect 44867 18340 44879 18343
rect 44867 18312 48176 18340
rect 44867 18309 44879 18312
rect 44821 18303 44879 18309
rect 48148 18284 48176 18312
rect 45373 18275 45431 18281
rect 45373 18241 45385 18275
rect 45419 18272 45431 18275
rect 45554 18272 45560 18284
rect 45419 18244 45560 18272
rect 45419 18241 45431 18244
rect 45373 18235 45431 18241
rect 45554 18232 45560 18244
rect 45612 18232 45618 18284
rect 46106 18232 46112 18284
rect 46164 18272 46170 18284
rect 46290 18272 46296 18284
rect 46164 18244 46296 18272
rect 46164 18232 46170 18244
rect 46290 18232 46296 18244
rect 46348 18232 46354 18284
rect 46474 18272 46480 18284
rect 46435 18244 46480 18272
rect 46474 18232 46480 18244
rect 46532 18232 46538 18284
rect 46845 18275 46903 18281
rect 46845 18241 46857 18275
rect 46891 18241 46903 18275
rect 46845 18235 46903 18241
rect 47029 18275 47087 18281
rect 47029 18241 47041 18275
rect 47075 18272 47087 18275
rect 47762 18272 47768 18284
rect 47075 18244 47768 18272
rect 47075 18241 47087 18244
rect 47029 18235 47087 18241
rect 45572 18136 45600 18232
rect 45922 18164 45928 18216
rect 45980 18204 45986 18216
rect 46385 18207 46443 18213
rect 46385 18204 46397 18207
rect 45980 18176 46397 18204
rect 45980 18164 45986 18176
rect 46385 18173 46397 18176
rect 46431 18173 46443 18207
rect 46385 18167 46443 18173
rect 45572 18108 46428 18136
rect 46106 18068 46112 18080
rect 46067 18040 46112 18068
rect 46106 18028 46112 18040
rect 46164 18028 46170 18080
rect 46400 18068 46428 18108
rect 46860 18068 46888 18235
rect 47762 18232 47768 18244
rect 47820 18232 47826 18284
rect 48130 18272 48136 18284
rect 48091 18244 48136 18272
rect 48130 18232 48136 18244
rect 48188 18232 48194 18284
rect 46400 18040 46888 18068
rect 47578 18028 47584 18080
rect 47636 18068 47642 18080
rect 47949 18071 48007 18077
rect 47949 18068 47961 18071
rect 47636 18040 47961 18068
rect 47636 18028 47642 18040
rect 47949 18037 47961 18040
rect 47995 18037 48007 18071
rect 47949 18031 48007 18037
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 46477 17799 46535 17805
rect 46477 17765 46489 17799
rect 46523 17796 46535 17799
rect 47946 17796 47952 17808
rect 46523 17768 47952 17796
rect 46523 17765 46535 17768
rect 46477 17759 46535 17765
rect 47946 17756 47952 17768
rect 48004 17756 48010 17808
rect 46842 17688 46848 17740
rect 46900 17728 46906 17740
rect 47397 17731 47455 17737
rect 47397 17728 47409 17731
rect 46900 17700 47409 17728
rect 46900 17688 46906 17700
rect 47397 17697 47409 17700
rect 47443 17697 47455 17731
rect 47397 17691 47455 17697
rect 47762 17688 47768 17740
rect 47820 17728 47826 17740
rect 47857 17731 47915 17737
rect 47857 17728 47869 17731
rect 47820 17700 47869 17728
rect 47820 17688 47826 17700
rect 47857 17697 47869 17700
rect 47903 17697 47915 17731
rect 47857 17691 47915 17697
rect 47581 17663 47639 17669
rect 47581 17629 47593 17663
rect 47627 17629 47639 17663
rect 47946 17660 47952 17672
rect 47907 17632 47952 17660
rect 47581 17623 47639 17629
rect 45554 17552 45560 17604
rect 45612 17592 45618 17604
rect 45830 17592 45836 17604
rect 45612 17564 45836 17592
rect 45612 17552 45618 17564
rect 45830 17552 45836 17564
rect 45888 17552 45894 17604
rect 46474 17552 46480 17604
rect 46532 17592 46538 17604
rect 47596 17592 47624 17623
rect 47946 17620 47952 17632
rect 48004 17620 48010 17672
rect 46532 17564 47624 17592
rect 46532 17552 46538 17564
rect 45922 17524 45928 17536
rect 45883 17496 45928 17524
rect 45922 17484 45928 17496
rect 45980 17484 45986 17536
rect 46566 17484 46572 17536
rect 46624 17524 46630 17536
rect 46750 17524 46756 17536
rect 46624 17496 46756 17524
rect 46624 17484 46630 17496
rect 46750 17484 46756 17496
rect 46808 17484 46814 17536
rect 47026 17524 47032 17536
rect 46987 17496 47032 17524
rect 47026 17484 47032 17496
rect 47084 17484 47090 17536
rect 47946 17484 47952 17536
rect 48004 17524 48010 17536
rect 48222 17524 48228 17536
rect 48004 17496 48228 17524
rect 48004 17484 48010 17496
rect 48222 17484 48228 17496
rect 48280 17484 48286 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 45922 17280 45928 17332
rect 45980 17320 45986 17332
rect 45980 17292 48176 17320
rect 45980 17280 45986 17292
rect 13998 17212 14004 17264
rect 14056 17252 14062 17264
rect 47026 17252 47032 17264
rect 14056 17224 47032 17252
rect 14056 17212 14062 17224
rect 47026 17212 47032 17224
rect 47084 17212 47090 17264
rect 47118 17212 47124 17264
rect 47176 17252 47182 17264
rect 47486 17252 47492 17264
rect 47176 17224 47492 17252
rect 47176 17212 47182 17224
rect 47486 17212 47492 17224
rect 47544 17212 47550 17264
rect 46477 17188 46535 17193
rect 46477 17187 46612 17188
rect 46477 17153 46489 17187
rect 46523 17160 46612 17187
rect 46523 17153 46535 17160
rect 46477 17147 46535 17153
rect 45646 17076 45652 17128
rect 45704 17116 45710 17128
rect 45833 17119 45891 17125
rect 45833 17116 45845 17119
rect 45704 17088 45845 17116
rect 45704 17076 45710 17088
rect 45833 17085 45845 17088
rect 45879 17085 45891 17119
rect 45833 17079 45891 17085
rect 45922 17076 45928 17128
rect 45980 17116 45986 17128
rect 46293 17119 46351 17125
rect 46293 17116 46305 17119
rect 45980 17088 46305 17116
rect 45980 17076 45986 17088
rect 46293 17085 46305 17088
rect 46339 17085 46351 17119
rect 46584 17116 46612 17160
rect 46750 17144 46756 17196
rect 46808 17184 46814 17196
rect 46845 17187 46903 17193
rect 46845 17184 46857 17187
rect 46808 17156 46857 17184
rect 46808 17144 46814 17156
rect 46845 17153 46857 17156
rect 46891 17153 46903 17187
rect 46845 17147 46903 17153
rect 46937 17187 46995 17193
rect 46937 17153 46949 17187
rect 46983 17184 46995 17187
rect 47762 17184 47768 17196
rect 46983 17156 47768 17184
rect 46983 17153 46995 17156
rect 46937 17147 46995 17153
rect 47762 17144 47768 17156
rect 47820 17144 47826 17196
rect 48148 17193 48176 17292
rect 48133 17187 48191 17193
rect 48133 17153 48145 17187
rect 48179 17184 48191 17187
rect 48222 17184 48228 17196
rect 48179 17156 48228 17184
rect 48179 17153 48191 17156
rect 48133 17147 48191 17153
rect 48222 17144 48228 17156
rect 48280 17144 48286 17196
rect 47578 17116 47584 17128
rect 46584 17088 47584 17116
rect 46293 17079 46351 17085
rect 47578 17076 47584 17088
rect 47636 17076 47642 17128
rect 45373 17051 45431 17057
rect 45373 17017 45385 17051
rect 45419 17048 45431 17051
rect 46750 17048 46756 17060
rect 45419 17020 46756 17048
rect 45419 17017 45431 17020
rect 45373 17011 45431 17017
rect 46750 17008 46756 17020
rect 46808 17008 46814 17060
rect 46566 16940 46572 16992
rect 46624 16980 46630 16992
rect 47949 16983 48007 16989
rect 47949 16980 47961 16983
rect 46624 16952 47961 16980
rect 46624 16940 46630 16952
rect 47949 16949 47961 16952
rect 47995 16949 48007 16983
rect 47949 16943 48007 16949
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 45833 16779 45891 16785
rect 45833 16745 45845 16779
rect 45879 16776 45891 16779
rect 46290 16776 46296 16788
rect 45879 16748 46296 16776
rect 45879 16745 45891 16748
rect 45833 16739 45891 16745
rect 46290 16736 46296 16748
rect 46348 16736 46354 16788
rect 46474 16776 46480 16788
rect 46435 16748 46480 16776
rect 46474 16736 46480 16748
rect 46532 16736 46538 16788
rect 46308 16708 46336 16736
rect 46308 16680 47992 16708
rect 45281 16643 45339 16649
rect 45281 16609 45293 16643
rect 45327 16640 45339 16643
rect 45327 16612 46336 16640
rect 45327 16609 45339 16612
rect 45281 16603 45339 16609
rect 46308 16584 46336 16612
rect 46290 16572 46296 16584
rect 46251 16544 46296 16572
rect 46290 16532 46296 16544
rect 46348 16532 46354 16584
rect 47394 16572 47400 16584
rect 47355 16544 47400 16572
rect 47394 16532 47400 16544
rect 47452 16532 47458 16584
rect 47578 16572 47584 16584
rect 47539 16544 47584 16572
rect 47578 16532 47584 16544
rect 47636 16532 47642 16584
rect 47964 16581 47992 16680
rect 47949 16575 48007 16581
rect 47949 16541 47961 16575
rect 47995 16541 48007 16575
rect 47949 16535 48007 16541
rect 48038 16532 48044 16584
rect 48096 16572 48102 16584
rect 48096 16544 48141 16572
rect 48096 16532 48102 16544
rect 45922 16464 45928 16516
rect 45980 16504 45986 16516
rect 46842 16504 46848 16516
rect 45980 16476 46848 16504
rect 45980 16464 45986 16476
rect 46842 16464 46848 16476
rect 46900 16464 46906 16516
rect 47026 16436 47032 16448
rect 46987 16408 47032 16436
rect 47026 16396 47032 16408
rect 47084 16396 47090 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 13262 16192 13268 16244
rect 13320 16232 13326 16244
rect 47026 16232 47032 16244
rect 13320 16204 47032 16232
rect 13320 16192 13326 16204
rect 47026 16192 47032 16204
rect 47084 16192 47090 16244
rect 47762 16232 47768 16244
rect 47723 16204 47768 16232
rect 47762 16192 47768 16204
rect 47820 16192 47826 16244
rect 44913 16099 44971 16105
rect 44913 16065 44925 16099
rect 44959 16096 44971 16099
rect 45922 16096 45928 16108
rect 44959 16068 45928 16096
rect 44959 16065 44971 16068
rect 44913 16059 44971 16065
rect 45922 16056 45928 16068
rect 45980 16056 45986 16108
rect 46474 16056 46480 16108
rect 46532 16096 46538 16108
rect 46569 16099 46627 16105
rect 46569 16096 46581 16099
rect 46532 16068 46581 16096
rect 46532 16056 46538 16068
rect 46569 16065 46581 16068
rect 46615 16065 46627 16099
rect 46569 16059 46627 16065
rect 46750 16056 46756 16108
rect 46808 16096 46814 16108
rect 47581 16099 47639 16105
rect 47581 16096 47593 16099
rect 46808 16068 47593 16096
rect 46808 16056 46814 16068
rect 47581 16065 47593 16068
rect 47627 16065 47639 16099
rect 47581 16059 47639 16065
rect 46109 15963 46167 15969
rect 46109 15929 46121 15963
rect 46155 15960 46167 15963
rect 47578 15960 47584 15972
rect 46155 15932 47584 15960
rect 46155 15929 46167 15932
rect 46109 15923 46167 15929
rect 47578 15920 47584 15932
rect 47636 15920 47642 15972
rect 45465 15895 45523 15901
rect 45465 15861 45477 15895
rect 45511 15892 45523 15895
rect 46290 15892 46296 15904
rect 45511 15864 46296 15892
rect 45511 15861 45523 15864
rect 45465 15855 45523 15861
rect 46290 15852 46296 15864
rect 46348 15852 46354 15904
rect 46753 15895 46811 15901
rect 46753 15861 46765 15895
rect 46799 15892 46811 15895
rect 46842 15892 46848 15904
rect 46799 15864 46848 15892
rect 46799 15861 46811 15864
rect 46753 15855 46811 15861
rect 46842 15852 46848 15864
rect 46900 15852 46906 15904
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 45281 15691 45339 15697
rect 45281 15657 45293 15691
rect 45327 15688 45339 15691
rect 48130 15688 48136 15700
rect 45327 15660 48136 15688
rect 45327 15657 45339 15660
rect 45281 15651 45339 15657
rect 48130 15648 48136 15660
rect 48188 15648 48194 15700
rect 46014 15580 46020 15632
rect 46072 15620 46078 15632
rect 46474 15620 46480 15632
rect 46072 15592 46480 15620
rect 46072 15580 46078 15592
rect 46474 15580 46480 15592
rect 46532 15580 46538 15632
rect 33134 15512 33140 15564
rect 33192 15552 33198 15564
rect 46937 15555 46995 15561
rect 46937 15552 46949 15555
rect 33192 15524 46949 15552
rect 33192 15512 33198 15524
rect 46937 15521 46949 15524
rect 46983 15521 46995 15555
rect 47394 15552 47400 15564
rect 47355 15524 47400 15552
rect 46937 15515 46995 15521
rect 47394 15512 47400 15524
rect 47452 15512 47458 15564
rect 47486 15512 47492 15564
rect 47544 15552 47550 15564
rect 47544 15524 47992 15552
rect 47544 15512 47550 15524
rect 46290 15484 46296 15496
rect 46251 15456 46296 15484
rect 46290 15444 46296 15456
rect 46348 15444 46354 15496
rect 47504 15484 47532 15512
rect 47964 15493 47992 15524
rect 46400 15456 47532 15484
rect 47581 15487 47639 15493
rect 45833 15419 45891 15425
rect 45833 15385 45845 15419
rect 45879 15416 45891 15419
rect 46400 15416 46428 15456
rect 47581 15453 47593 15487
rect 47627 15453 47639 15487
rect 47581 15447 47639 15453
rect 47949 15487 48007 15493
rect 47949 15453 47961 15487
rect 47995 15453 48007 15487
rect 47949 15447 48007 15453
rect 47596 15416 47624 15447
rect 48038 15444 48044 15496
rect 48096 15484 48102 15496
rect 48096 15456 48141 15484
rect 48096 15444 48102 15456
rect 45879 15388 46428 15416
rect 46492 15388 47624 15416
rect 45879 15385 45891 15388
rect 45833 15379 45891 15385
rect 46492 15357 46520 15388
rect 46477 15351 46535 15357
rect 46477 15317 46489 15351
rect 46523 15317 46535 15351
rect 46477 15311 46535 15317
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 45554 15104 45560 15156
rect 45612 15144 45618 15156
rect 46842 15144 46848 15156
rect 45612 15116 46848 15144
rect 45612 15104 45618 15116
rect 46842 15104 46848 15116
rect 46900 15104 46906 15156
rect 44729 15079 44787 15085
rect 44729 15045 44741 15079
rect 44775 15076 44787 15079
rect 48406 15076 48412 15088
rect 44775 15048 48412 15076
rect 44775 15045 44787 15048
rect 44729 15039 44787 15045
rect 44177 15011 44235 15017
rect 44177 14977 44189 15011
rect 44223 15008 44235 15011
rect 45189 15011 45247 15017
rect 45189 15008 45201 15011
rect 44223 14980 45201 15008
rect 44223 14977 44235 14980
rect 44177 14971 44235 14977
rect 45189 14977 45201 14980
rect 45235 15008 45247 15011
rect 45554 15008 45560 15020
rect 45235 14980 45560 15008
rect 45235 14977 45247 14980
rect 45189 14971 45247 14977
rect 45554 14968 45560 14980
rect 45612 14968 45618 15020
rect 46477 15011 46535 15017
rect 46477 14977 46489 15011
rect 46523 15008 46535 15011
rect 46566 15008 46572 15020
rect 46523 14980 46572 15008
rect 46523 14977 46535 14980
rect 46477 14971 46535 14977
rect 46566 14968 46572 14980
rect 46624 14968 46630 15020
rect 46860 15017 46888 15048
rect 48406 15036 48412 15048
rect 48464 15036 48470 15088
rect 46845 15011 46903 15017
rect 46845 14977 46857 15011
rect 46891 14977 46903 15011
rect 46845 14971 46903 14977
rect 47026 14968 47032 15020
rect 47084 15008 47090 15020
rect 48038 15008 48044 15020
rect 47084 14980 48044 15008
rect 47084 14968 47090 14980
rect 48038 14968 48044 14980
rect 48096 14968 48102 15020
rect 48130 14968 48136 15020
rect 48188 15008 48194 15020
rect 48188 14980 48233 15008
rect 48188 14968 48194 14980
rect 37918 14900 37924 14952
rect 37976 14940 37982 14952
rect 45833 14943 45891 14949
rect 45833 14940 45845 14943
rect 37976 14912 45845 14940
rect 37976 14900 37982 14912
rect 45833 14909 45845 14912
rect 45879 14909 45891 14943
rect 45833 14903 45891 14909
rect 46385 14943 46443 14949
rect 46385 14909 46397 14943
rect 46431 14940 46443 14943
rect 47394 14940 47400 14952
rect 46431 14912 47400 14940
rect 46431 14909 46443 14912
rect 46385 14903 46443 14909
rect 47394 14900 47400 14912
rect 47452 14900 47458 14952
rect 45373 14807 45431 14813
rect 45373 14773 45385 14807
rect 45419 14804 45431 14807
rect 46474 14804 46480 14816
rect 45419 14776 46480 14804
rect 45419 14773 45431 14776
rect 45373 14767 45431 14773
rect 46474 14764 46480 14776
rect 46532 14764 46538 14816
rect 47578 14764 47584 14816
rect 47636 14804 47642 14816
rect 47949 14807 48007 14813
rect 47949 14804 47961 14807
rect 47636 14776 47961 14804
rect 47636 14764 47642 14776
rect 47949 14773 47961 14776
rect 47995 14773 48007 14807
rect 47949 14767 48007 14773
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 46385 14603 46443 14609
rect 46385 14569 46397 14603
rect 46431 14600 46443 14603
rect 47026 14600 47032 14612
rect 46431 14572 47032 14600
rect 46431 14569 46443 14572
rect 46385 14563 46443 14569
rect 47026 14560 47032 14572
rect 47084 14560 47090 14612
rect 45649 14535 45707 14541
rect 45649 14501 45661 14535
rect 45695 14501 45707 14535
rect 45649 14495 45707 14501
rect 45664 14464 45692 14495
rect 47394 14464 47400 14476
rect 45664 14436 47400 14464
rect 47394 14424 47400 14436
rect 47452 14424 47458 14476
rect 45465 14399 45523 14405
rect 45465 14365 45477 14399
rect 45511 14396 45523 14399
rect 46014 14396 46020 14408
rect 45511 14368 46020 14396
rect 45511 14365 45523 14368
rect 45465 14359 45523 14365
rect 46014 14356 46020 14368
rect 46072 14356 46078 14408
rect 46201 14399 46259 14405
rect 46201 14365 46213 14399
rect 46247 14396 46259 14399
rect 46750 14396 46756 14408
rect 46247 14368 46756 14396
rect 46247 14365 46259 14368
rect 46201 14359 46259 14365
rect 46750 14356 46756 14368
rect 46808 14356 46814 14408
rect 47578 14396 47584 14408
rect 47539 14368 47584 14396
rect 47578 14356 47584 14368
rect 47636 14356 47642 14408
rect 47762 14356 47768 14408
rect 47820 14396 47826 14408
rect 47949 14399 48007 14405
rect 47949 14396 47961 14399
rect 47820 14368 47961 14396
rect 47820 14356 47826 14368
rect 47949 14365 47961 14368
rect 47995 14365 48007 14399
rect 47949 14359 48007 14365
rect 48038 14356 48044 14408
rect 48096 14396 48102 14408
rect 48096 14368 48141 14396
rect 48096 14356 48102 14368
rect 27338 14288 27344 14340
rect 27396 14328 27402 14340
rect 46937 14331 46995 14337
rect 46937 14328 46949 14331
rect 27396 14300 46949 14328
rect 27396 14288 27402 14300
rect 46937 14297 46949 14300
rect 46983 14297 46995 14331
rect 46937 14291 46995 14297
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 2133 14059 2191 14065
rect 2133 14025 2145 14059
rect 2179 14025 2191 14059
rect 2133 14019 2191 14025
rect 45373 14059 45431 14065
rect 45373 14025 45385 14059
rect 45419 14056 45431 14059
rect 47762 14056 47768 14068
rect 45419 14028 47768 14056
rect 45419 14025 45431 14028
rect 45373 14019 45431 14025
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 2148 13920 2176 14019
rect 47762 14016 47768 14028
rect 47820 14016 47826 14068
rect 44821 13991 44879 13997
rect 44821 13957 44833 13991
rect 44867 13988 44879 13991
rect 44867 13960 46888 13988
rect 44867 13957 44879 13960
rect 44821 13951 44879 13957
rect 46860 13932 46888 13960
rect 1719 13892 2176 13920
rect 2317 13923 2375 13929
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 2317 13889 2329 13923
rect 2363 13889 2375 13923
rect 46474 13920 46480 13932
rect 46435 13892 46480 13920
rect 2317 13883 2375 13889
rect 658 13812 664 13864
rect 716 13852 722 13864
rect 2332 13852 2360 13883
rect 46474 13880 46480 13892
rect 46532 13880 46538 13932
rect 46842 13920 46848 13932
rect 46803 13892 46848 13920
rect 46842 13880 46848 13892
rect 46900 13880 46906 13932
rect 47026 13920 47032 13932
rect 46987 13892 47032 13920
rect 47026 13880 47032 13892
rect 47084 13880 47090 13932
rect 48038 13880 48044 13932
rect 48096 13920 48102 13932
rect 48133 13923 48191 13929
rect 48133 13920 48145 13923
rect 48096 13892 48145 13920
rect 48096 13880 48102 13892
rect 48133 13889 48145 13892
rect 48179 13889 48191 13923
rect 48133 13883 48191 13889
rect 2777 13855 2835 13861
rect 2777 13852 2789 13855
rect 716 13824 2789 13852
rect 716 13812 722 13824
rect 2777 13821 2789 13824
rect 2823 13852 2835 13855
rect 4614 13852 4620 13864
rect 2823 13824 4620 13852
rect 2823 13821 2835 13824
rect 2777 13815 2835 13821
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 36630 13812 36636 13864
rect 36688 13852 36694 13864
rect 45833 13855 45891 13861
rect 45833 13852 45845 13855
rect 36688 13824 45845 13852
rect 36688 13812 36694 13824
rect 45833 13821 45845 13824
rect 45879 13821 45891 13855
rect 45833 13815 45891 13821
rect 46569 13855 46627 13861
rect 46569 13821 46581 13855
rect 46615 13852 46627 13855
rect 47394 13852 47400 13864
rect 46615 13824 47400 13852
rect 46615 13821 46627 13824
rect 46569 13815 46627 13821
rect 47394 13812 47400 13824
rect 47452 13812 47458 13864
rect 1486 13784 1492 13796
rect 1447 13756 1492 13784
rect 1486 13744 1492 13756
rect 1544 13744 1550 13796
rect 47578 13676 47584 13728
rect 47636 13716 47642 13728
rect 47949 13719 48007 13725
rect 47949 13716 47961 13719
rect 47636 13688 47961 13716
rect 47636 13676 47642 13688
rect 47949 13685 47961 13688
rect 47995 13685 48007 13719
rect 47949 13679 48007 13685
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 45281 13515 45339 13521
rect 45281 13481 45293 13515
rect 45327 13512 45339 13515
rect 48038 13512 48044 13524
rect 45327 13484 48044 13512
rect 45327 13481 45339 13484
rect 45281 13475 45339 13481
rect 48038 13472 48044 13484
rect 48096 13512 48102 13524
rect 48222 13512 48228 13524
rect 48096 13484 48228 13512
rect 48096 13472 48102 13484
rect 48222 13472 48228 13484
rect 48280 13472 48286 13524
rect 45833 13379 45891 13385
rect 45833 13345 45845 13379
rect 45879 13376 45891 13379
rect 46934 13376 46940 13388
rect 45879 13348 46940 13376
rect 45879 13345 45891 13348
rect 45833 13339 45891 13345
rect 46934 13336 46940 13348
rect 46992 13376 46998 13388
rect 46992 13348 47992 13376
rect 46992 13336 46998 13348
rect 44453 13311 44511 13317
rect 44453 13277 44465 13311
rect 44499 13308 44511 13311
rect 46290 13308 46296 13320
rect 44499 13280 46296 13308
rect 44499 13277 44511 13280
rect 44453 13271 44511 13277
rect 46290 13268 46296 13280
rect 46348 13268 46354 13320
rect 46566 13268 46572 13320
rect 46624 13308 46630 13320
rect 47397 13311 47455 13317
rect 47397 13308 47409 13311
rect 46624 13280 47409 13308
rect 46624 13268 46630 13280
rect 47397 13277 47409 13280
rect 47443 13277 47455 13311
rect 47578 13308 47584 13320
rect 47539 13280 47584 13308
rect 47397 13271 47455 13277
rect 47578 13268 47584 13280
rect 47636 13268 47642 13320
rect 47964 13317 47992 13348
rect 47949 13311 48007 13317
rect 47949 13277 47961 13311
rect 47995 13277 48007 13311
rect 47949 13271 48007 13277
rect 48038 13268 48044 13320
rect 48096 13308 48102 13320
rect 48096 13280 48141 13308
rect 48096 13268 48102 13280
rect 46474 13172 46480 13184
rect 46435 13144 46480 13172
rect 46474 13132 46480 13144
rect 46532 13132 46538 13184
rect 47026 13172 47032 13184
rect 46987 13144 47032 13172
rect 47026 13132 47032 13144
rect 47084 13132 47090 13184
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 47026 12968 47032 12980
rect 8352 12940 47032 12968
rect 8352 12928 8358 12940
rect 47026 12928 47032 12940
rect 47084 12928 47090 12980
rect 45186 12860 45192 12912
rect 45244 12900 45250 12912
rect 45830 12900 45836 12912
rect 45244 12872 45836 12900
rect 45244 12860 45250 12872
rect 45830 12860 45836 12872
rect 45888 12860 45894 12912
rect 47946 12900 47952 12912
rect 46308 12872 47952 12900
rect 45373 12835 45431 12841
rect 45373 12801 45385 12835
rect 45419 12832 45431 12835
rect 46308 12832 46336 12872
rect 46474 12832 46480 12844
rect 45419 12804 46336 12832
rect 46435 12804 46480 12832
rect 45419 12801 45431 12804
rect 45373 12795 45431 12801
rect 46474 12792 46480 12804
rect 46532 12792 46538 12844
rect 46860 12841 46888 12872
rect 47946 12860 47952 12872
rect 48004 12860 48010 12912
rect 46845 12835 46903 12841
rect 46845 12801 46857 12835
rect 46891 12801 46903 12835
rect 46845 12795 46903 12801
rect 46934 12792 46940 12844
rect 46992 12832 46998 12844
rect 47029 12835 47087 12841
rect 47029 12832 47041 12835
rect 46992 12804 47041 12832
rect 46992 12792 46998 12804
rect 47029 12801 47041 12804
rect 47075 12832 47087 12835
rect 48038 12832 48044 12844
rect 47075 12804 48044 12832
rect 47075 12801 47087 12804
rect 47029 12795 47087 12801
rect 48038 12792 48044 12804
rect 48096 12792 48102 12844
rect 48133 12835 48191 12841
rect 48133 12801 48145 12835
rect 48179 12801 48191 12835
rect 48133 12795 48191 12801
rect 45646 12724 45652 12776
rect 45704 12764 45710 12776
rect 45833 12767 45891 12773
rect 45833 12764 45845 12767
rect 45704 12736 45845 12764
rect 45704 12724 45710 12736
rect 45833 12733 45845 12736
rect 45879 12733 45891 12767
rect 46566 12764 46572 12776
rect 46527 12736 46572 12764
rect 45833 12727 45891 12733
rect 46566 12724 46572 12736
rect 46624 12724 46630 12776
rect 48148 12764 48176 12795
rect 47504 12736 48176 12764
rect 44821 12699 44879 12705
rect 44821 12665 44833 12699
rect 44867 12696 44879 12699
rect 46584 12696 46612 12724
rect 46842 12696 46848 12708
rect 44867 12668 46520 12696
rect 46584 12668 46848 12696
rect 44867 12665 44879 12668
rect 44821 12659 44879 12665
rect 46014 12588 46020 12640
rect 46072 12628 46078 12640
rect 46382 12628 46388 12640
rect 46072 12600 46388 12628
rect 46072 12588 46078 12600
rect 46382 12588 46388 12600
rect 46440 12588 46446 12640
rect 46492 12628 46520 12668
rect 46842 12656 46848 12668
rect 46900 12656 46906 12708
rect 46750 12628 46756 12640
rect 46492 12600 46756 12628
rect 46750 12588 46756 12600
rect 46808 12628 46814 12640
rect 47504 12628 47532 12736
rect 46808 12600 47532 12628
rect 46808 12588 46814 12600
rect 47578 12588 47584 12640
rect 47636 12628 47642 12640
rect 47949 12631 48007 12637
rect 47949 12628 47961 12631
rect 47636 12600 47961 12628
rect 47636 12588 47642 12600
rect 47949 12597 47961 12600
rect 47995 12597 48007 12631
rect 47949 12591 48007 12597
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 45278 12384 45284 12436
rect 45336 12424 45342 12436
rect 46477 12427 46535 12433
rect 46477 12424 46489 12427
rect 45336 12396 46489 12424
rect 45336 12384 45342 12396
rect 46477 12393 46489 12396
rect 46523 12393 46535 12427
rect 46477 12387 46535 12393
rect 45833 12359 45891 12365
rect 45833 12325 45845 12359
rect 45879 12356 45891 12359
rect 45879 12328 47716 12356
rect 45879 12325 45891 12328
rect 45833 12319 45891 12325
rect 46014 12248 46020 12300
rect 46072 12288 46078 12300
rect 46566 12288 46572 12300
rect 46072 12260 46572 12288
rect 46072 12248 46078 12260
rect 46566 12248 46572 12260
rect 46624 12248 46630 12300
rect 45281 12223 45339 12229
rect 45281 12189 45293 12223
rect 45327 12220 45339 12223
rect 46290 12220 46296 12232
rect 45327 12192 46296 12220
rect 45327 12189 45339 12192
rect 45281 12183 45339 12189
rect 46290 12180 46296 12192
rect 46348 12180 46354 12232
rect 46474 12220 46480 12232
rect 46400 12192 46480 12220
rect 46400 12152 46428 12192
rect 46474 12180 46480 12192
rect 46532 12180 46538 12232
rect 46842 12180 46848 12232
rect 46900 12220 46906 12232
rect 47397 12223 47455 12229
rect 47397 12220 47409 12223
rect 46900 12192 47409 12220
rect 46900 12180 46906 12192
rect 47397 12189 47409 12192
rect 47443 12189 47455 12223
rect 47578 12220 47584 12232
rect 47539 12192 47584 12220
rect 47397 12183 47455 12189
rect 47578 12180 47584 12192
rect 47636 12180 47642 12232
rect 47688 12220 47716 12328
rect 47857 12291 47915 12297
rect 47857 12257 47869 12291
rect 47903 12288 47915 12291
rect 48038 12288 48044 12300
rect 47903 12260 48044 12288
rect 47903 12257 47915 12260
rect 47857 12251 47915 12257
rect 48038 12248 48044 12260
rect 48096 12248 48102 12300
rect 47949 12223 48007 12229
rect 47949 12220 47961 12223
rect 47688 12192 47961 12220
rect 47949 12189 47961 12192
rect 47995 12220 48007 12223
rect 48961 12223 49019 12229
rect 48961 12220 48973 12223
rect 47995 12192 48973 12220
rect 47995 12189 48007 12192
rect 47949 12183 48007 12189
rect 48961 12189 48973 12192
rect 49007 12189 49019 12223
rect 48961 12183 49019 12189
rect 46124 12124 46428 12152
rect 46124 12096 46152 12124
rect 45554 12044 45560 12096
rect 45612 12084 45618 12096
rect 46014 12084 46020 12096
rect 45612 12056 46020 12084
rect 45612 12044 45618 12056
rect 46014 12044 46020 12056
rect 46072 12044 46078 12096
rect 46106 12044 46112 12096
rect 46164 12044 46170 12096
rect 47026 12084 47032 12096
rect 46987 12056 47032 12084
rect 47026 12044 47032 12056
rect 47084 12044 47090 12096
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 25222 11840 25228 11892
rect 25280 11880 25286 11892
rect 47026 11880 47032 11892
rect 25280 11852 47032 11880
rect 25280 11840 25286 11852
rect 47026 11840 47032 11852
rect 47084 11840 47090 11892
rect 45373 11815 45431 11821
rect 45373 11781 45385 11815
rect 45419 11812 45431 11815
rect 45922 11812 45928 11824
rect 45419 11784 45928 11812
rect 45419 11781 45431 11784
rect 45373 11775 45431 11781
rect 45922 11772 45928 11784
rect 45980 11812 45986 11824
rect 45980 11784 46888 11812
rect 45980 11772 45986 11784
rect 45278 11704 45284 11756
rect 45336 11744 45342 11756
rect 46860 11753 46888 11784
rect 46477 11747 46535 11753
rect 46477 11744 46489 11747
rect 45336 11716 46489 11744
rect 45336 11704 45342 11716
rect 46477 11713 46489 11716
rect 46523 11713 46535 11747
rect 46477 11707 46535 11713
rect 46845 11747 46903 11753
rect 46845 11713 46857 11747
rect 46891 11713 46903 11747
rect 46845 11707 46903 11713
rect 46934 11704 46940 11756
rect 46992 11744 46998 11756
rect 48130 11744 48136 11756
rect 46992 11716 47037 11744
rect 48091 11716 48136 11744
rect 46992 11704 46998 11716
rect 48130 11704 48136 11716
rect 48188 11704 48194 11756
rect 45554 11636 45560 11688
rect 45612 11676 45618 11688
rect 45833 11679 45891 11685
rect 45833 11676 45845 11679
rect 45612 11648 45845 11676
rect 45612 11636 45618 11648
rect 45833 11645 45845 11648
rect 45879 11645 45891 11679
rect 45833 11639 45891 11645
rect 46569 11679 46627 11685
rect 46569 11645 46581 11679
rect 46615 11645 46627 11679
rect 46569 11639 46627 11645
rect 46584 11608 46612 11639
rect 46842 11608 46848 11620
rect 46584 11580 46848 11608
rect 46842 11568 46848 11580
rect 46900 11568 46906 11620
rect 48130 11608 48136 11620
rect 47320 11580 48136 11608
rect 1854 11500 1860 11552
rect 1912 11540 1918 11552
rect 2041 11543 2099 11549
rect 2041 11540 2053 11543
rect 1912 11512 2053 11540
rect 1912 11500 1918 11512
rect 2041 11509 2053 11512
rect 2087 11509 2099 11543
rect 2041 11503 2099 11509
rect 44821 11543 44879 11549
rect 44821 11509 44833 11543
rect 44867 11540 44879 11543
rect 47320 11540 47348 11580
rect 48130 11568 48136 11580
rect 48188 11568 48194 11620
rect 44867 11512 47348 11540
rect 44867 11509 44879 11512
rect 44821 11503 44879 11509
rect 47578 11500 47584 11552
rect 47636 11540 47642 11552
rect 47949 11543 48007 11549
rect 47949 11540 47961 11543
rect 47636 11512 47961 11540
rect 47636 11500 47642 11512
rect 47949 11509 47961 11512
rect 47995 11509 48007 11543
rect 47949 11503 48007 11509
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 46385 11339 46443 11345
rect 46385 11305 46397 11339
rect 46431 11336 46443 11339
rect 46934 11336 46940 11348
rect 46431 11308 46940 11336
rect 46431 11305 46443 11308
rect 46385 11299 46443 11305
rect 46934 11296 46940 11308
rect 46992 11296 46998 11348
rect 45922 11228 45928 11280
rect 45980 11268 45986 11280
rect 46106 11268 46112 11280
rect 45980 11240 46112 11268
rect 45980 11228 45986 11240
rect 46106 11228 46112 11240
rect 46164 11228 46170 11280
rect 45738 11200 45744 11212
rect 45651 11172 45744 11200
rect 45738 11160 45744 11172
rect 45796 11200 45802 11212
rect 45796 11172 46520 11200
rect 45796 11160 45802 11172
rect 45830 11092 45836 11144
rect 45888 11132 45894 11144
rect 46106 11132 46112 11144
rect 45888 11104 46112 11132
rect 45888 11092 45894 11104
rect 46106 11092 46112 11104
rect 46164 11132 46170 11144
rect 46201 11135 46259 11141
rect 46201 11132 46213 11135
rect 46164 11104 46213 11132
rect 46164 11092 46170 11104
rect 46201 11101 46213 11104
rect 46247 11101 46259 11135
rect 46492 11132 46520 11172
rect 46842 11160 46848 11212
rect 46900 11200 46906 11212
rect 47397 11203 47455 11209
rect 47397 11200 47409 11203
rect 46900 11172 47409 11200
rect 46900 11160 46906 11172
rect 47397 11169 47409 11172
rect 47443 11169 47455 11203
rect 47397 11163 47455 11169
rect 47578 11132 47584 11144
rect 46492 11104 47072 11132
rect 47539 11104 47584 11132
rect 46201 11095 46259 11101
rect 1578 11024 1584 11076
rect 1636 11064 1642 11076
rect 1765 11067 1823 11073
rect 1765 11064 1777 11067
rect 1636 11036 1777 11064
rect 1636 11024 1642 11036
rect 1765 11033 1777 11036
rect 1811 11033 1823 11067
rect 2590 11064 2596 11076
rect 2551 11036 2596 11064
rect 1765 11027 1823 11033
rect 2590 11024 2596 11036
rect 2648 11024 2654 11076
rect 3145 11067 3203 11073
rect 3145 11033 3157 11067
rect 3191 11064 3203 11067
rect 3418 11064 3424 11076
rect 3191 11036 3424 11064
rect 3191 11033 3203 11036
rect 3145 11027 3203 11033
rect 3418 11024 3424 11036
rect 3476 11024 3482 11076
rect 3881 11067 3939 11073
rect 3881 11033 3893 11067
rect 3927 11064 3939 11067
rect 3970 11064 3976 11076
rect 3927 11036 3976 11064
rect 3927 11033 3939 11036
rect 3881 11027 3939 11033
rect 3970 11024 3976 11036
rect 4028 11024 4034 11076
rect 4433 11067 4491 11073
rect 4433 11033 4445 11067
rect 4479 11064 4491 11067
rect 4614 11064 4620 11076
rect 4479 11036 4620 11064
rect 4479 11033 4491 11036
rect 4433 11027 4491 11033
rect 4614 11024 4620 11036
rect 4672 11024 4678 11076
rect 4985 11067 5043 11073
rect 4985 11033 4997 11067
rect 5031 11064 5043 11067
rect 5442 11064 5448 11076
rect 5031 11036 5448 11064
rect 5031 11033 5043 11036
rect 4985 11027 5043 11033
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 15286 11024 15292 11076
rect 15344 11064 15350 11076
rect 46937 11067 46995 11073
rect 46937 11064 46949 11067
rect 15344 11036 46949 11064
rect 15344 11024 15350 11036
rect 46937 11033 46949 11036
rect 46983 11033 46995 11067
rect 47044 11064 47072 11104
rect 47578 11092 47584 11104
rect 47636 11092 47642 11144
rect 47949 11135 48007 11141
rect 47949 11101 47961 11135
rect 47995 11101 48007 11135
rect 47949 11095 48007 11101
rect 47964 11064 47992 11095
rect 48038 11092 48044 11144
rect 48096 11132 48102 11144
rect 48096 11104 48141 11132
rect 48096 11092 48102 11104
rect 47044 11036 47992 11064
rect 46937 11027 46995 11033
rect 45186 10956 45192 11008
rect 45244 10996 45250 11008
rect 45738 10996 45744 11008
rect 45244 10968 45744 10996
rect 45244 10956 45250 10968
rect 45738 10956 45744 10968
rect 45796 10956 45802 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 46753 10795 46811 10801
rect 46753 10761 46765 10795
rect 46799 10792 46811 10795
rect 46842 10792 46848 10804
rect 46799 10764 46848 10792
rect 46799 10761 46811 10764
rect 46753 10755 46811 10761
rect 46842 10752 46848 10764
rect 46900 10752 46906 10804
rect 45922 10616 45928 10668
rect 45980 10656 45986 10668
rect 46382 10656 46388 10668
rect 45980 10628 46388 10656
rect 45980 10616 45986 10628
rect 46382 10616 46388 10628
rect 46440 10656 46446 10668
rect 46569 10659 46627 10665
rect 46569 10656 46581 10659
rect 46440 10628 46581 10656
rect 46440 10616 46446 10628
rect 46569 10625 46581 10628
rect 46615 10625 46627 10659
rect 46569 10619 46627 10625
rect 48133 10659 48191 10665
rect 48133 10625 48145 10659
rect 48179 10656 48191 10659
rect 48222 10656 48228 10668
rect 48179 10628 48228 10656
rect 48179 10625 48191 10628
rect 48133 10619 48191 10625
rect 45557 10591 45615 10597
rect 45557 10557 45569 10591
rect 45603 10588 45615 10591
rect 48148 10588 48176 10619
rect 48222 10616 48228 10628
rect 48280 10616 48286 10668
rect 45603 10560 48176 10588
rect 45603 10557 45615 10560
rect 45557 10551 45615 10557
rect 3878 10480 3884 10532
rect 3936 10520 3942 10532
rect 4249 10523 4307 10529
rect 4249 10520 4261 10523
rect 3936 10492 4261 10520
rect 3936 10480 3942 10492
rect 4249 10489 4261 10492
rect 4295 10489 4307 10523
rect 4249 10483 4307 10489
rect 1489 10455 1547 10461
rect 1489 10421 1501 10455
rect 1535 10452 1547 10455
rect 1670 10452 1676 10464
rect 1535 10424 1676 10452
rect 1535 10421 1547 10424
rect 1489 10415 1547 10421
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 2041 10455 2099 10461
rect 2041 10421 2053 10455
rect 2087 10452 2099 10455
rect 2130 10452 2136 10464
rect 2087 10424 2136 10452
rect 2087 10421 2099 10424
rect 2041 10415 2099 10421
rect 2130 10412 2136 10424
rect 2188 10412 2194 10464
rect 2222 10412 2228 10464
rect 2280 10452 2286 10464
rect 2501 10455 2559 10461
rect 2501 10452 2513 10455
rect 2280 10424 2513 10452
rect 2280 10412 2286 10424
rect 2501 10421 2513 10424
rect 2547 10421 2559 10455
rect 2501 10415 2559 10421
rect 3237 10455 3295 10461
rect 3237 10421 3249 10455
rect 3283 10452 3295 10455
rect 3510 10452 3516 10464
rect 3283 10424 3516 10452
rect 3283 10421 3295 10424
rect 3237 10415 3295 10421
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 3789 10455 3847 10461
rect 3789 10421 3801 10455
rect 3835 10452 3847 10455
rect 4062 10452 4068 10464
rect 3835 10424 4068 10452
rect 3835 10421 3847 10424
rect 3789 10415 3847 10421
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4706 10412 4712 10464
rect 4764 10452 4770 10464
rect 4801 10455 4859 10461
rect 4801 10452 4813 10455
rect 4764 10424 4813 10452
rect 4764 10412 4770 10424
rect 4801 10421 4813 10424
rect 4847 10421 4859 10455
rect 5350 10452 5356 10464
rect 5311 10424 5356 10452
rect 4801 10415 4859 10421
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 46109 10455 46167 10461
rect 46109 10421 46121 10455
rect 46155 10452 46167 10455
rect 46934 10452 46940 10464
rect 46155 10424 46940 10452
rect 46155 10421 46167 10424
rect 46109 10415 46167 10421
rect 46934 10412 46940 10424
rect 46992 10412 46998 10464
rect 47578 10412 47584 10464
rect 47636 10452 47642 10464
rect 47949 10455 48007 10461
rect 47949 10452 47961 10455
rect 47636 10424 47961 10452
rect 47636 10412 47642 10424
rect 47949 10421 47961 10424
rect 47995 10421 48007 10455
rect 47949 10415 48007 10421
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 45738 10248 45744 10260
rect 45699 10220 45744 10248
rect 45738 10208 45744 10220
rect 45796 10208 45802 10260
rect 45756 10112 45784 10208
rect 45756 10084 47992 10112
rect 2498 10004 2504 10056
rect 2556 10044 2562 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 2556 10016 3801 10044
rect 2556 10004 2562 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3878 10004 3884 10056
rect 3936 10044 3942 10056
rect 4154 10044 4160 10056
rect 3936 10016 4160 10044
rect 3936 10004 3942 10016
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 45281 10047 45339 10053
rect 45281 10013 45293 10047
rect 45327 10044 45339 10047
rect 46290 10044 46296 10056
rect 45327 10016 46296 10044
rect 45327 10013 45339 10016
rect 45281 10007 45339 10013
rect 46290 10004 46296 10016
rect 46348 10004 46354 10056
rect 47394 10044 47400 10056
rect 47355 10016 47400 10044
rect 47394 10004 47400 10016
rect 47452 10004 47458 10056
rect 47578 10044 47584 10056
rect 47539 10016 47584 10044
rect 47578 10004 47584 10016
rect 47636 10004 47642 10056
rect 47964 10053 47992 10084
rect 47949 10047 48007 10053
rect 47949 10013 47961 10047
rect 47995 10013 48007 10047
rect 47949 10007 48007 10013
rect 48038 10004 48044 10056
rect 48096 10044 48102 10056
rect 48096 10016 48141 10044
rect 48096 10004 48102 10016
rect 934 9936 940 9988
rect 992 9976 998 9988
rect 1949 9979 2007 9985
rect 1949 9976 1961 9979
rect 992 9948 1961 9976
rect 992 9936 998 9948
rect 1949 9945 1961 9948
rect 1995 9945 2007 9979
rect 1949 9939 2007 9945
rect 2038 9936 2044 9988
rect 2096 9976 2102 9988
rect 3053 9979 3111 9985
rect 3053 9976 3065 9979
rect 2096 9948 3065 9976
rect 2096 9936 2102 9948
rect 3053 9945 3065 9948
rect 3099 9945 3111 9979
rect 3053 9939 3111 9945
rect 750 9868 756 9920
rect 808 9908 814 9920
rect 1210 9908 1216 9920
rect 808 9880 1216 9908
rect 808 9868 814 9880
rect 1210 9868 1216 9880
rect 1268 9868 1274 9920
rect 1394 9908 1400 9920
rect 1355 9880 1400 9908
rect 1394 9868 1400 9880
rect 1452 9868 1458 9920
rect 2406 9868 2412 9920
rect 2464 9908 2470 9920
rect 2501 9911 2559 9917
rect 2501 9908 2513 9911
rect 2464 9880 2513 9908
rect 2464 9868 2470 9880
rect 2501 9877 2513 9880
rect 2547 9877 2559 9911
rect 2501 9871 2559 9877
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 4341 9911 4399 9917
rect 4341 9908 4353 9911
rect 2832 9880 4353 9908
rect 2832 9868 2838 9880
rect 4341 9877 4353 9880
rect 4387 9877 4399 9911
rect 5166 9908 5172 9920
rect 5127 9880 5172 9908
rect 4341 9871 4399 9877
rect 5166 9868 5172 9880
rect 5224 9868 5230 9920
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 5813 9911 5871 9917
rect 5813 9908 5825 9911
rect 5592 9880 5825 9908
rect 5592 9868 5598 9880
rect 5813 9877 5825 9880
rect 5859 9877 5871 9911
rect 6454 9908 6460 9920
rect 6415 9880 6460 9908
rect 5813 9871 5871 9877
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 46474 9908 46480 9920
rect 46435 9880 46480 9908
rect 46474 9868 46480 9880
rect 46532 9868 46538 9920
rect 47026 9908 47032 9920
rect 46987 9880 47032 9908
rect 47026 9868 47032 9880
rect 47084 9868 47090 9920
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 1210 9664 1216 9716
rect 1268 9704 1274 9716
rect 2682 9704 2688 9716
rect 1268 9676 2688 9704
rect 1268 9664 1274 9676
rect 2682 9664 2688 9676
rect 2740 9664 2746 9716
rect 6454 9664 6460 9716
rect 6512 9704 6518 9716
rect 47026 9704 47032 9716
rect 6512 9676 47032 9704
rect 6512 9664 6518 9676
rect 47026 9664 47032 9676
rect 47084 9664 47090 9716
rect 1302 9596 1308 9648
rect 1360 9636 1366 9648
rect 6270 9636 6276 9648
rect 1360 9608 6276 9636
rect 1360 9596 1366 9608
rect 6270 9596 6276 9608
rect 6328 9596 6334 9648
rect 7374 9596 7380 9648
rect 7432 9636 7438 9648
rect 8113 9639 8171 9645
rect 8113 9636 8125 9639
rect 7432 9608 8125 9636
rect 7432 9596 7438 9608
rect 8113 9605 8125 9608
rect 8159 9636 8171 9639
rect 8294 9636 8300 9648
rect 8159 9608 8300 9636
rect 8159 9605 8171 9608
rect 8113 9599 8171 9605
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 45373 9639 45431 9645
rect 45373 9605 45385 9639
rect 45419 9636 45431 9639
rect 46658 9636 46664 9648
rect 45419 9608 46664 9636
rect 45419 9605 45431 9608
rect 45373 9599 45431 9605
rect 46658 9596 46664 9608
rect 46716 9596 46722 9648
rect 46934 9596 46940 9648
rect 46992 9636 46998 9648
rect 46992 9608 48176 9636
rect 46992 9596 46998 9608
rect 48148 9580 48176 9608
rect 46474 9568 46480 9580
rect 46435 9540 46480 9568
rect 46474 9528 46480 9540
rect 46532 9528 46538 9580
rect 46845 9571 46903 9577
rect 46845 9537 46857 9571
rect 46891 9537 46903 9571
rect 46845 9531 46903 9537
rect 47029 9571 47087 9577
rect 47029 9537 47041 9571
rect 47075 9568 47087 9571
rect 48038 9568 48044 9580
rect 47075 9540 48044 9568
rect 47075 9537 47087 9540
rect 47029 9531 47087 9537
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 2501 9503 2559 9509
rect 2501 9500 2513 9503
rect 2004 9472 2513 9500
rect 2004 9460 2010 9472
rect 2501 9469 2513 9472
rect 2547 9469 2559 9503
rect 2501 9463 2559 9469
rect 8386 9460 8392 9512
rect 8444 9500 8450 9512
rect 8665 9503 8723 9509
rect 8665 9500 8677 9503
rect 8444 9472 8677 9500
rect 8444 9460 8450 9472
rect 8665 9469 8677 9472
rect 8711 9500 8723 9503
rect 27338 9500 27344 9512
rect 8711 9472 27344 9500
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 27338 9460 27344 9472
rect 27396 9460 27402 9512
rect 45830 9500 45836 9512
rect 45791 9472 45836 9500
rect 45830 9460 45836 9472
rect 45888 9460 45894 9512
rect 46569 9503 46627 9509
rect 46569 9469 46581 9503
rect 46615 9500 46627 9503
rect 46750 9500 46756 9512
rect 46615 9472 46756 9500
rect 46615 9469 46627 9472
rect 46569 9463 46627 9469
rect 46750 9460 46756 9472
rect 46808 9460 46814 9512
rect 46860 9500 46888 9531
rect 48038 9528 48044 9540
rect 48096 9528 48102 9580
rect 48130 9528 48136 9580
rect 48188 9568 48194 9580
rect 48188 9540 48233 9568
rect 48188 9528 48194 9540
rect 49053 9503 49111 9509
rect 49053 9500 49065 9503
rect 46860 9472 49065 9500
rect 4522 9392 4528 9444
rect 4580 9432 4586 9444
rect 5074 9432 5080 9444
rect 4580 9404 5080 9432
rect 4580 9392 4586 9404
rect 5074 9392 5080 9404
rect 5132 9392 5138 9444
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 7561 9435 7619 9441
rect 7561 9432 7573 9435
rect 7064 9404 7573 9432
rect 7064 9392 7070 9404
rect 7561 9401 7573 9404
rect 7607 9432 7619 9435
rect 45554 9432 45560 9444
rect 7607 9404 45560 9432
rect 7607 9401 7619 9404
rect 7561 9395 7619 9401
rect 45554 9392 45560 9404
rect 45612 9392 45618 9444
rect 1486 9364 1492 9376
rect 1447 9336 1492 9364
rect 1486 9324 1492 9336
rect 1544 9324 1550 9376
rect 1762 9324 1768 9376
rect 1820 9364 1826 9376
rect 1949 9367 2007 9373
rect 1949 9364 1961 9367
rect 1820 9336 1961 9364
rect 1820 9324 1826 9336
rect 1949 9333 1961 9336
rect 1995 9333 2007 9367
rect 1949 9327 2007 9333
rect 2866 9324 2872 9376
rect 2924 9364 2930 9376
rect 3053 9367 3111 9373
rect 3053 9364 3065 9367
rect 2924 9336 3065 9364
rect 2924 9324 2930 9336
rect 3053 9333 3065 9336
rect 3099 9333 3111 9367
rect 3694 9364 3700 9376
rect 3655 9336 3700 9364
rect 3053 9327 3111 9333
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 4433 9367 4491 9373
rect 4433 9333 4445 9367
rect 4479 9364 4491 9367
rect 4614 9364 4620 9376
rect 4479 9336 4620 9364
rect 4479 9333 4491 9336
rect 4433 9327 4491 9333
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 4893 9367 4951 9373
rect 4893 9364 4905 9367
rect 4856 9336 4905 9364
rect 4856 9324 4862 9336
rect 4893 9333 4905 9336
rect 4939 9333 4951 9367
rect 4893 9327 4951 9333
rect 5258 9324 5264 9376
rect 5316 9364 5322 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 5316 9336 5549 9364
rect 5316 9324 5322 9336
rect 5537 9333 5549 9336
rect 5583 9333 5595 9367
rect 6362 9364 6368 9376
rect 6323 9336 6368 9364
rect 5537 9327 5595 9333
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 6917 9367 6975 9373
rect 6917 9364 6929 9367
rect 6788 9336 6929 9364
rect 6788 9324 6794 9336
rect 6917 9333 6929 9336
rect 6963 9333 6975 9367
rect 6917 9327 6975 9333
rect 44821 9367 44879 9373
rect 44821 9333 44833 9367
rect 44867 9364 44879 9367
rect 46860 9364 46888 9472
rect 49053 9469 49065 9472
rect 49099 9469 49111 9503
rect 49053 9463 49111 9469
rect 47946 9364 47952 9376
rect 44867 9336 46888 9364
rect 47907 9336 47952 9364
rect 44867 9333 44879 9336
rect 44821 9327 44879 9333
rect 47946 9324 47952 9336
rect 48004 9324 48010 9376
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 5718 9160 5724 9172
rect 1627 9132 5724 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 6730 9120 6736 9172
rect 6788 9160 6794 9172
rect 45830 9160 45836 9172
rect 6788 9132 45836 9160
rect 6788 9120 6794 9132
rect 45830 9120 45836 9132
rect 45888 9120 45894 9172
rect 46382 9160 46388 9172
rect 46295 9132 46388 9160
rect 46382 9120 46388 9132
rect 46440 9160 46446 9172
rect 46750 9160 46756 9172
rect 46440 9132 46756 9160
rect 46440 9120 46446 9132
rect 46750 9120 46756 9132
rect 46808 9160 46814 9172
rect 47394 9160 47400 9172
rect 46808 9132 47400 9160
rect 46808 9120 46814 9132
rect 47394 9120 47400 9132
rect 47452 9120 47458 9172
rect 45646 9092 45652 9104
rect 35866 9064 45652 9092
rect 382 8916 388 8968
rect 440 8956 446 8968
rect 1394 8956 1400 8968
rect 440 8928 1400 8956
rect 440 8916 446 8928
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 7101 8959 7159 8965
rect 7101 8956 7113 8959
rect 5684 8928 7113 8956
rect 5684 8916 5690 8928
rect 7101 8925 7113 8928
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 33134 8956 33140 8968
rect 9732 8928 33140 8956
rect 9732 8916 9738 8928
rect 33134 8916 33140 8928
rect 33192 8916 33198 8968
rect 4982 8888 4988 8900
rect 2746 8860 4988 8888
rect 2314 8780 2320 8832
rect 2372 8820 2378 8832
rect 2409 8823 2467 8829
rect 2409 8820 2421 8823
rect 2372 8792 2421 8820
rect 2372 8780 2378 8792
rect 2409 8789 2421 8792
rect 2455 8820 2467 8823
rect 2746 8820 2774 8860
rect 4982 8848 4988 8860
rect 5040 8848 5046 8900
rect 6641 8891 6699 8897
rect 6641 8857 6653 8891
rect 6687 8888 6699 8891
rect 7282 8888 7288 8900
rect 6687 8860 7288 8888
rect 6687 8857 6699 8860
rect 6641 8851 6699 8857
rect 7282 8848 7288 8860
rect 7340 8848 7346 8900
rect 8110 8848 8116 8900
rect 8168 8888 8174 8900
rect 8938 8888 8944 8900
rect 8168 8860 8944 8888
rect 8168 8848 8174 8860
rect 8938 8848 8944 8860
rect 8996 8848 9002 8900
rect 35866 8888 35894 9064
rect 45646 9052 45652 9064
rect 45704 9052 45710 9104
rect 45741 9095 45799 9101
rect 45741 9061 45753 9095
rect 45787 9092 45799 9095
rect 47210 9092 47216 9104
rect 45787 9064 47216 9092
rect 45787 9061 45799 9064
rect 45741 9055 45799 9061
rect 47210 9052 47216 9064
rect 47268 9052 47274 9104
rect 47394 9024 47400 9036
rect 47355 8996 47400 9024
rect 47394 8984 47400 8996
rect 47452 8984 47458 9036
rect 48314 9024 48320 9036
rect 47964 8996 48320 9024
rect 45186 8916 45192 8968
rect 45244 8956 45250 8968
rect 46198 8956 46204 8968
rect 45244 8928 46204 8956
rect 45244 8916 45250 8928
rect 46198 8916 46204 8928
rect 46256 8916 46262 8968
rect 46290 8916 46296 8968
rect 46348 8956 46354 8968
rect 47964 8965 47992 8996
rect 48314 8984 48320 8996
rect 48372 8984 48378 9036
rect 47581 8959 47639 8965
rect 47581 8956 47593 8959
rect 46348 8928 47593 8956
rect 46348 8916 46354 8928
rect 47581 8925 47593 8928
rect 47627 8925 47639 8959
rect 47581 8919 47639 8925
rect 47949 8959 48007 8965
rect 47949 8925 47961 8959
rect 47995 8925 48007 8959
rect 47949 8919 48007 8925
rect 9508 8860 35894 8888
rect 2958 8820 2964 8832
rect 2455 8792 2774 8820
rect 2919 8792 2964 8820
rect 2455 8789 2467 8792
rect 2409 8783 2467 8789
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 3602 8780 3608 8832
rect 3660 8820 3666 8832
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3660 8792 3801 8820
rect 3660 8780 3666 8792
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 4338 8820 4344 8832
rect 4299 8792 4344 8820
rect 3789 8783 3847 8789
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 4890 8820 4896 8832
rect 4851 8792 4896 8820
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 5537 8823 5595 8829
rect 5537 8789 5549 8823
rect 5583 8820 5595 8823
rect 5902 8820 5908 8832
rect 5583 8792 5908 8820
rect 5583 8789 5595 8792
rect 5537 8783 5595 8789
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 6089 8823 6147 8829
rect 6089 8789 6101 8823
rect 6135 8820 6147 8823
rect 6178 8820 6184 8832
rect 6135 8792 6184 8820
rect 6135 8789 6147 8792
rect 6089 8783 6147 8789
rect 6178 8780 6184 8792
rect 6236 8780 6242 8832
rect 7190 8780 7196 8832
rect 7248 8820 7254 8832
rect 7653 8823 7711 8829
rect 7653 8820 7665 8823
rect 7248 8792 7665 8820
rect 7248 8780 7254 8792
rect 7653 8789 7665 8792
rect 7699 8789 7711 8823
rect 7653 8783 7711 8789
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 8297 8823 8355 8829
rect 8297 8820 8309 8823
rect 7800 8792 8309 8820
rect 7800 8780 7806 8792
rect 8297 8789 8309 8792
rect 8343 8789 8355 8823
rect 8297 8783 8355 8789
rect 9214 8780 9220 8832
rect 9272 8820 9278 8832
rect 9508 8829 9536 8860
rect 37642 8848 37648 8900
rect 37700 8888 37706 8900
rect 46937 8891 46995 8897
rect 46937 8888 46949 8891
rect 37700 8860 46949 8888
rect 37700 8848 37706 8860
rect 46937 8857 46949 8860
rect 46983 8857 46995 8891
rect 46937 8851 46995 8857
rect 9493 8823 9551 8829
rect 9493 8820 9505 8823
rect 9272 8792 9505 8820
rect 9272 8780 9278 8792
rect 9493 8789 9505 8792
rect 9539 8789 9551 8823
rect 9493 8783 9551 8789
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 10045 8823 10103 8829
rect 10045 8820 10057 8823
rect 9732 8792 10057 8820
rect 9732 8780 9738 8792
rect 10045 8789 10057 8792
rect 10091 8789 10103 8823
rect 10045 8783 10103 8789
rect 45189 8823 45247 8829
rect 45189 8789 45201 8823
rect 45235 8820 45247 8823
rect 47964 8820 47992 8919
rect 48038 8916 48044 8968
rect 48096 8956 48102 8968
rect 48096 8928 48141 8956
rect 48096 8916 48102 8928
rect 45235 8792 47992 8820
rect 45235 8789 45247 8792
rect 45189 8783 45247 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8585 2191 8619
rect 5074 8616 5080 8628
rect 2133 8579 2191 8585
rect 4908 8588 5080 8616
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 2148 8480 2176 8579
rect 4908 8560 4936 8588
rect 5074 8576 5080 8588
rect 5132 8576 5138 8628
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 44634 8616 44640 8628
rect 8996 8588 40724 8616
rect 44595 8588 44640 8616
rect 8996 8576 9002 8588
rect 4890 8508 4896 8560
rect 4948 8508 4954 8560
rect 4982 8508 4988 8560
rect 5040 8548 5046 8560
rect 5166 8548 5172 8560
rect 5040 8520 5172 8548
rect 5040 8508 5046 8520
rect 5166 8508 5172 8520
rect 5224 8548 5230 8560
rect 37642 8548 37648 8560
rect 5224 8520 37648 8548
rect 5224 8508 5230 8520
rect 37642 8508 37648 8520
rect 37700 8508 37706 8560
rect 40696 8548 40724 8588
rect 44634 8576 44640 8588
rect 44692 8576 44698 8628
rect 47765 8619 47823 8625
rect 47765 8585 47777 8619
rect 47811 8616 47823 8619
rect 48038 8616 48044 8628
rect 47811 8588 48044 8616
rect 47811 8585 47823 8588
rect 47765 8579 47823 8585
rect 45833 8551 45891 8557
rect 45833 8548 45845 8551
rect 40696 8520 45845 8548
rect 45833 8517 45845 8520
rect 45879 8517 45891 8551
rect 45833 8511 45891 8517
rect 46750 8508 46756 8560
rect 46808 8548 46814 8560
rect 47780 8548 47808 8579
rect 48038 8576 48044 8588
rect 48096 8576 48102 8628
rect 46808 8520 47808 8548
rect 46808 8508 46814 8520
rect 2314 8480 2320 8492
rect 1719 8452 2176 8480
rect 2275 8452 2320 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 3421 8483 3479 8489
rect 3421 8480 3433 8483
rect 3384 8452 3433 8480
rect 3384 8440 3390 8452
rect 3421 8449 3433 8452
rect 3467 8480 3479 8483
rect 4065 8483 4123 8489
rect 4065 8480 4077 8483
rect 3467 8452 4077 8480
rect 3467 8449 3479 8452
rect 3421 8443 3479 8449
rect 4065 8449 4077 8452
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 5074 8480 5080 8492
rect 4764 8452 5080 8480
rect 4764 8440 4770 8452
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 44177 8483 44235 8489
rect 44177 8449 44189 8483
rect 44223 8480 44235 8483
rect 45189 8483 45247 8489
rect 45189 8480 45201 8483
rect 44223 8452 45201 8480
rect 44223 8449 44235 8452
rect 44177 8443 44235 8449
rect 45189 8449 45201 8452
rect 45235 8480 45247 8483
rect 46477 8483 46535 8489
rect 46477 8480 46489 8483
rect 45235 8452 45324 8480
rect 45235 8449 45247 8452
rect 45189 8443 45247 8449
rect 7193 8415 7251 8421
rect 7193 8381 7205 8415
rect 7239 8412 7251 8415
rect 7834 8412 7840 8424
rect 7239 8384 7840 8412
rect 7239 8381 7251 8384
rect 7193 8375 7251 8381
rect 7834 8372 7840 8384
rect 7892 8372 7898 8424
rect 1486 8344 1492 8356
rect 1447 8316 1492 8344
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 4706 8344 4712 8356
rect 4667 8316 4712 8344
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 5166 8344 5172 8356
rect 5127 8316 5172 8344
rect 5166 8304 5172 8316
rect 5224 8304 5230 8356
rect 5810 8344 5816 8356
rect 5771 8316 5816 8344
rect 5810 8304 5816 8316
rect 5868 8304 5874 8356
rect 7650 8344 7656 8356
rect 7611 8316 7656 8344
rect 7650 8304 7656 8316
rect 7708 8304 7714 8356
rect 2869 8279 2927 8285
rect 2869 8245 2881 8279
rect 2915 8276 2927 8279
rect 3234 8276 3240 8288
rect 2915 8248 3240 8276
rect 2915 8245 2927 8248
rect 2869 8239 2927 8245
rect 3234 8236 3240 8248
rect 3292 8236 3298 8288
rect 3605 8279 3663 8285
rect 3605 8245 3617 8279
rect 3651 8276 3663 8279
rect 3878 8276 3884 8288
rect 3651 8248 3884 8276
rect 3651 8245 3663 8248
rect 3605 8239 3663 8245
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 6086 8236 6092 8288
rect 6144 8276 6150 8288
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 6144 8248 6561 8276
rect 6144 8236 6150 8248
rect 6549 8245 6561 8248
rect 6595 8245 6607 8279
rect 8202 8276 8208 8288
rect 8163 8248 8208 8276
rect 6549 8239 6607 8245
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 8662 8236 8668 8288
rect 8720 8276 8726 8288
rect 8757 8279 8815 8285
rect 8757 8276 8769 8279
rect 8720 8248 8769 8276
rect 8720 8236 8726 8248
rect 8757 8245 8769 8248
rect 8803 8245 8815 8279
rect 9306 8276 9312 8288
rect 9267 8248 9312 8276
rect 8757 8239 8815 8245
rect 9306 8236 9312 8248
rect 9364 8236 9370 8288
rect 9858 8276 9864 8288
rect 9819 8248 9864 8276
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 10410 8276 10416 8288
rect 10371 8248 10416 8276
rect 10410 8236 10416 8248
rect 10468 8236 10474 8288
rect 45296 8276 45324 8452
rect 45388 8452 46489 8480
rect 45388 8353 45416 8452
rect 46477 8449 46489 8452
rect 46523 8449 46535 8483
rect 46477 8443 46535 8449
rect 46658 8440 46664 8492
rect 46716 8480 46722 8492
rect 47044 8489 47072 8520
rect 46845 8483 46903 8489
rect 46845 8480 46857 8483
rect 46716 8452 46857 8480
rect 46716 8440 46722 8452
rect 46845 8449 46857 8452
rect 46891 8449 46903 8483
rect 46845 8443 46903 8449
rect 47029 8483 47087 8489
rect 47029 8449 47041 8483
rect 47075 8449 47087 8483
rect 47029 8443 47087 8449
rect 47581 8483 47639 8489
rect 47581 8449 47593 8483
rect 47627 8449 47639 8483
rect 47581 8443 47639 8449
rect 46382 8412 46388 8424
rect 46343 8384 46388 8412
rect 46382 8372 46388 8384
rect 46440 8372 46446 8424
rect 45373 8347 45431 8353
rect 45373 8313 45385 8347
rect 45419 8313 45431 8347
rect 45554 8344 45560 8356
rect 45373 8307 45431 8313
rect 45480 8316 45560 8344
rect 45480 8276 45508 8316
rect 45554 8304 45560 8316
rect 45612 8304 45618 8356
rect 45738 8304 45744 8356
rect 45796 8344 45802 8356
rect 47486 8344 47492 8356
rect 45796 8316 47492 8344
rect 45796 8304 45802 8316
rect 47486 8304 47492 8316
rect 47544 8344 47550 8356
rect 47596 8344 47624 8443
rect 47544 8316 47624 8344
rect 47544 8304 47550 8316
rect 45296 8248 45508 8276
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 2038 8072 2044 8084
rect 1544 8044 2044 8072
rect 1544 8032 1550 8044
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 45738 8032 45744 8084
rect 45796 8072 45802 8084
rect 45833 8075 45891 8081
rect 45833 8072 45845 8075
rect 45796 8044 45845 8072
rect 45796 8032 45802 8044
rect 45833 8041 45845 8044
rect 45879 8041 45891 8075
rect 45833 8035 45891 8041
rect 46477 8075 46535 8081
rect 46477 8041 46489 8075
rect 46523 8072 46535 8075
rect 47118 8072 47124 8084
rect 46523 8044 47124 8072
rect 46523 8041 46535 8044
rect 46477 8035 46535 8041
rect 47118 8032 47124 8044
rect 47176 8032 47182 8084
rect 45189 8007 45247 8013
rect 45189 7973 45201 8007
rect 45235 8004 45247 8007
rect 47670 8004 47676 8016
rect 45235 7976 47676 8004
rect 45235 7973 45247 7976
rect 45189 7967 45247 7973
rect 47670 7964 47676 7976
rect 47728 7964 47734 8016
rect 750 7896 756 7948
rect 808 7936 814 7948
rect 7558 7936 7564 7948
rect 808 7908 7564 7936
rect 808 7896 814 7908
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 14826 7896 14832 7948
rect 14884 7936 14890 7948
rect 30374 7936 30380 7948
rect 14884 7908 30380 7936
rect 14884 7896 14890 7908
rect 30374 7896 30380 7908
rect 30432 7896 30438 7948
rect 47210 7896 47216 7948
rect 47268 7936 47274 7948
rect 47268 7908 47992 7936
rect 47268 7896 47274 7908
rect 290 7828 296 7880
rect 348 7868 354 7880
rect 1394 7868 1400 7880
rect 348 7840 1400 7868
rect 348 7828 354 7840
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7868 2283 7871
rect 2498 7868 2504 7880
rect 2271 7840 2504 7868
rect 2271 7837 2283 7840
rect 2225 7831 2283 7837
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2832 7840 2881 7868
rect 2832 7828 2838 7840
rect 2869 7837 2881 7840
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4062 7868 4068 7880
rect 4019 7840 4068 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 4522 7828 4528 7880
rect 4580 7868 4586 7880
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 4580 7840 4629 7868
rect 4580 7828 4586 7840
rect 4617 7837 4629 7840
rect 4663 7868 4675 7871
rect 5077 7871 5135 7877
rect 5077 7868 5089 7871
rect 4663 7840 5089 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 5077 7837 5089 7840
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 15378 7828 15384 7880
rect 15436 7868 15442 7880
rect 36630 7868 36636 7880
rect 15436 7840 36636 7868
rect 15436 7828 15442 7840
rect 36630 7828 36636 7840
rect 36688 7828 36694 7880
rect 45646 7868 45652 7880
rect 45607 7840 45652 7868
rect 45646 7828 45652 7840
rect 45704 7868 45710 7880
rect 46106 7868 46112 7880
rect 45704 7840 46112 7868
rect 45704 7828 45710 7840
rect 46106 7828 46112 7840
rect 46164 7828 46170 7880
rect 47394 7868 47400 7880
rect 47355 7840 47400 7868
rect 47394 7828 47400 7840
rect 47452 7828 47458 7880
rect 47578 7868 47584 7880
rect 47539 7840 47584 7868
rect 47578 7828 47584 7840
rect 47636 7828 47642 7880
rect 47964 7877 47992 7908
rect 47949 7871 48007 7877
rect 47949 7837 47961 7871
rect 47995 7837 48007 7871
rect 47949 7831 48007 7837
rect 48038 7828 48044 7880
rect 48096 7868 48102 7880
rect 48096 7840 48141 7868
rect 48096 7828 48102 7840
rect 5721 7803 5779 7809
rect 5721 7769 5733 7803
rect 5767 7800 5779 7803
rect 6546 7800 6552 7812
rect 5767 7772 6552 7800
rect 5767 7769 5779 7772
rect 5721 7763 5779 7769
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 15838 7760 15844 7812
rect 15896 7800 15902 7812
rect 39298 7800 39304 7812
rect 15896 7772 39304 7800
rect 15896 7760 15902 7772
rect 39298 7760 39304 7772
rect 39356 7760 39362 7812
rect 43809 7803 43867 7809
rect 43809 7769 43821 7803
rect 43855 7800 43867 7803
rect 44542 7800 44548 7812
rect 43855 7772 44548 7800
rect 43855 7769 43867 7772
rect 43809 7763 43867 7769
rect 44542 7760 44548 7772
rect 44600 7760 44606 7812
rect 44634 7760 44640 7812
rect 44692 7800 44698 7812
rect 45462 7800 45468 7812
rect 44692 7772 45468 7800
rect 44692 7760 44698 7772
rect 45462 7760 45468 7772
rect 45520 7760 45526 7812
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 2038 7732 2044 7744
rect 1627 7704 2044 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 2406 7732 2412 7744
rect 2367 7704 2412 7732
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 3050 7732 3056 7744
rect 3011 7704 3056 7732
rect 3050 7692 3056 7704
rect 3108 7692 3114 7744
rect 3786 7732 3792 7744
rect 3747 7704 3792 7732
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 4430 7732 4436 7744
rect 4391 7704 4436 7732
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 6638 7732 6644 7744
rect 6599 7704 6644 7732
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 7466 7732 7472 7744
rect 7427 7704 7472 7732
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 8018 7732 8024 7744
rect 7979 7704 8024 7732
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 9033 7735 9091 7741
rect 9033 7701 9045 7735
rect 9079 7732 9091 7735
rect 9582 7732 9588 7744
rect 9079 7704 9588 7732
rect 9079 7701 9091 7704
rect 9033 7695 9091 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 9766 7732 9772 7744
rect 9727 7704 9772 7732
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 10134 7692 10140 7744
rect 10192 7732 10198 7744
rect 10229 7735 10287 7741
rect 10229 7732 10241 7735
rect 10192 7704 10241 7732
rect 10192 7692 10198 7704
rect 10229 7701 10241 7704
rect 10275 7701 10287 7735
rect 10778 7732 10784 7744
rect 10739 7704 10784 7732
rect 10229 7695 10287 7701
rect 10778 7692 10784 7704
rect 10836 7692 10842 7744
rect 11330 7732 11336 7744
rect 11291 7704 11336 7732
rect 11330 7692 11336 7704
rect 11388 7692 11394 7744
rect 43070 7692 43076 7744
rect 43128 7732 43134 7744
rect 44266 7732 44272 7744
rect 43128 7704 44272 7732
rect 43128 7692 43134 7704
rect 44266 7692 44272 7704
rect 44324 7692 44330 7744
rect 47026 7732 47032 7744
rect 46987 7704 47032 7732
rect 47026 7692 47032 7704
rect 47084 7692 47090 7744
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 2682 7528 2688 7540
rect 2643 7500 2688 7528
rect 2682 7488 2688 7500
rect 2740 7488 2746 7540
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 6880 7500 9137 7528
rect 6880 7488 6886 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9125 7491 9183 7497
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 47026 7528 47032 7540
rect 11112 7500 47032 7528
rect 11112 7488 11118 7500
rect 47026 7488 47032 7500
rect 47084 7488 47090 7540
rect 2314 7460 2320 7472
rect 1412 7432 2320 7460
rect 1412 7401 1440 7432
rect 2314 7420 2320 7432
rect 2372 7420 2378 7472
rect 44266 7420 44272 7472
rect 44324 7460 44330 7472
rect 44545 7463 44603 7469
rect 44324 7432 44404 7460
rect 44324 7420 44330 7432
rect 661 7395 719 7401
rect 661 7361 673 7395
rect 707 7392 719 7395
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 707 7364 1409 7392
rect 707 7361 719 7364
rect 661 7355 719 7361
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7392 2099 7395
rect 2222 7392 2228 7404
rect 2087 7364 2228 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 937 7327 995 7333
rect 937 7293 949 7327
rect 983 7324 995 7327
rect 2056 7324 2084 7355
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 2869 7395 2927 7401
rect 2869 7392 2881 7395
rect 2746 7364 2881 7392
rect 2746 7324 2774 7364
rect 2869 7361 2881 7364
rect 2915 7361 2927 7395
rect 3510 7392 3516 7404
rect 3471 7364 3516 7392
rect 2869 7355 2927 7361
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 4706 7392 4712 7404
rect 4571 7364 4712 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5258 7392 5264 7404
rect 5215 7364 5264 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5684 7364 5825 7392
rect 5684 7352 5690 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 6362 7392 6368 7404
rect 6052 7364 6368 7392
rect 6052 7352 6058 7364
rect 6362 7352 6368 7364
rect 6420 7392 6426 7404
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 6420 7364 6561 7392
rect 6420 7352 6426 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 7190 7392 7196 7404
rect 7151 7364 7196 7392
rect 6549 7355 6607 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7742 7352 7748 7404
rect 7800 7392 7806 7404
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 7800 7364 7849 7392
rect 7800 7352 7806 7364
rect 7837 7361 7849 7364
rect 7883 7361 7895 7395
rect 8662 7392 8668 7404
rect 8623 7364 8668 7392
rect 7837 7355 7895 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 9306 7392 9312 7404
rect 9219 7364 9312 7392
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 9490 7352 9496 7404
rect 9548 7392 9554 7404
rect 10229 7395 10287 7401
rect 10229 7392 10241 7395
rect 9548 7364 10241 7392
rect 9548 7352 9554 7364
rect 10229 7361 10241 7364
rect 10275 7392 10287 7395
rect 10410 7392 10416 7404
rect 10275 7364 10416 7392
rect 10275 7361 10287 7364
rect 10229 7355 10287 7361
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 12158 7352 12164 7404
rect 12216 7392 12222 7404
rect 43070 7392 43076 7404
rect 12216 7364 43076 7392
rect 12216 7352 12222 7364
rect 43070 7352 43076 7364
rect 43128 7352 43134 7404
rect 43162 7352 43168 7404
rect 43220 7392 43226 7404
rect 43809 7395 43867 7401
rect 43809 7392 43821 7395
rect 43220 7364 43821 7392
rect 43220 7352 43226 7364
rect 43809 7361 43821 7364
rect 43855 7361 43867 7395
rect 43809 7355 43867 7361
rect 43901 7395 43959 7401
rect 43901 7361 43913 7395
rect 43947 7392 43959 7395
rect 44082 7392 44088 7404
rect 43947 7364 44088 7392
rect 43947 7361 43959 7364
rect 43901 7355 43959 7361
rect 44082 7352 44088 7364
rect 44140 7352 44146 7404
rect 44376 7392 44404 7432
rect 44545 7429 44557 7463
rect 44591 7460 44603 7463
rect 45646 7460 45652 7472
rect 44591 7432 45652 7460
rect 44591 7429 44603 7432
rect 44545 7423 44603 7429
rect 45646 7420 45652 7432
rect 45704 7420 45710 7472
rect 47946 7460 47952 7472
rect 46492 7432 47952 7460
rect 44453 7395 44511 7401
rect 44453 7392 44465 7395
rect 44376 7364 44465 7392
rect 44453 7361 44465 7364
rect 44499 7361 44511 7395
rect 45094 7392 45100 7404
rect 45007 7364 45100 7392
rect 44453 7355 44511 7361
rect 45094 7352 45100 7364
rect 45152 7392 45158 7404
rect 45922 7392 45928 7404
rect 45152 7364 45928 7392
rect 45152 7352 45158 7364
rect 45922 7352 45928 7364
rect 45980 7352 45986 7404
rect 46492 7401 46520 7432
rect 47946 7420 47952 7432
rect 48004 7420 48010 7472
rect 46477 7395 46535 7401
rect 46477 7361 46489 7395
rect 46523 7361 46535 7395
rect 46477 7355 46535 7361
rect 46845 7395 46903 7401
rect 46845 7361 46857 7395
rect 46891 7361 46903 7395
rect 46845 7355 46903 7361
rect 983 7296 2084 7324
rect 2240 7296 2774 7324
rect 983 7293 995 7296
rect 937 7287 995 7293
rect 845 7259 903 7265
rect 845 7225 857 7259
rect 891 7256 903 7259
rect 1394 7256 1400 7268
rect 891 7228 1400 7256
rect 891 7225 903 7228
rect 845 7219 903 7225
rect 1394 7216 1400 7228
rect 1452 7256 1458 7268
rect 2240 7256 2268 7296
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 9324 7324 9352 7352
rect 11517 7327 11575 7333
rect 11517 7324 11529 7327
rect 8628 7296 9352 7324
rect 10244 7296 11529 7324
rect 8628 7284 8634 7296
rect 10244 7268 10272 7296
rect 11517 7293 11529 7296
rect 11563 7293 11575 7327
rect 11517 7287 11575 7293
rect 16758 7284 16764 7336
rect 16816 7324 16822 7336
rect 45833 7327 45891 7333
rect 45833 7324 45845 7327
rect 16816 7296 45845 7324
rect 16816 7284 16822 7296
rect 45833 7293 45845 7296
rect 45879 7293 45891 7327
rect 46382 7324 46388 7336
rect 46343 7296 46388 7324
rect 45833 7287 45891 7293
rect 46382 7284 46388 7296
rect 46440 7284 46446 7336
rect 46750 7324 46756 7336
rect 46711 7296 46756 7324
rect 46750 7284 46756 7296
rect 46808 7284 46814 7336
rect 1452 7228 2268 7256
rect 1452 7216 1458 7228
rect 2314 7216 2320 7268
rect 2372 7256 2378 7268
rect 3329 7259 3387 7265
rect 3329 7256 3341 7259
rect 2372 7228 3341 7256
rect 2372 7216 2378 7228
rect 3329 7225 3341 7228
rect 3375 7225 3387 7259
rect 3329 7219 3387 7225
rect 10226 7216 10232 7268
rect 10284 7216 10290 7268
rect 10413 7259 10471 7265
rect 10413 7225 10425 7259
rect 10459 7256 10471 7259
rect 11974 7256 11980 7268
rect 10459 7228 11980 7256
rect 10459 7225 10471 7228
rect 10413 7219 10471 7225
rect 11974 7216 11980 7228
rect 12032 7216 12038 7268
rect 12713 7259 12771 7265
rect 12713 7225 12725 7259
rect 12759 7256 12771 7259
rect 12802 7256 12808 7268
rect 12759 7228 12808 7256
rect 12759 7225 12771 7228
rect 12713 7219 12771 7225
rect 12802 7216 12808 7228
rect 12860 7256 12866 7268
rect 12860 7228 22094 7256
rect 12860 7216 12866 7228
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 2225 7191 2283 7197
rect 2225 7157 2237 7191
rect 2271 7188 2283 7191
rect 2774 7188 2780 7200
rect 2271 7160 2780 7188
rect 2271 7157 2283 7160
rect 2225 7151 2283 7157
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 3970 7148 3976 7200
rect 4028 7188 4034 7200
rect 4341 7191 4399 7197
rect 4341 7188 4353 7191
rect 4028 7160 4353 7188
rect 4028 7148 4034 7160
rect 4341 7157 4353 7160
rect 4387 7157 4399 7191
rect 4982 7188 4988 7200
rect 4943 7160 4988 7188
rect 4341 7151 4399 7157
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 5626 7188 5632 7200
rect 5587 7160 5632 7188
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 6362 7188 6368 7200
rect 6323 7160 6368 7188
rect 6362 7148 6368 7160
rect 6420 7148 6426 7200
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7009 7191 7067 7197
rect 7009 7188 7021 7191
rect 6972 7160 7021 7188
rect 6972 7148 6978 7160
rect 7009 7157 7021 7160
rect 7055 7157 7067 7191
rect 7009 7151 7067 7157
rect 7926 7148 7932 7200
rect 7984 7188 7990 7200
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 7984 7160 8033 7188
rect 7984 7148 7990 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8481 7191 8539 7197
rect 8481 7188 8493 7191
rect 8352 7160 8493 7188
rect 8352 7148 8358 7160
rect 8481 7157 8493 7160
rect 8527 7157 8539 7191
rect 8481 7151 8539 7157
rect 10686 7148 10692 7200
rect 10744 7188 10750 7200
rect 10873 7191 10931 7197
rect 10873 7188 10885 7191
rect 10744 7160 10885 7188
rect 10744 7148 10750 7160
rect 10873 7157 10885 7160
rect 10919 7157 10931 7191
rect 10873 7151 10931 7157
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 12069 7191 12127 7197
rect 12069 7188 12081 7191
rect 11756 7160 12081 7188
rect 11756 7148 11762 7160
rect 12069 7157 12081 7160
rect 12115 7157 12127 7191
rect 22066 7188 22094 7228
rect 41386 7228 44036 7256
rect 41386 7188 41414 7228
rect 42794 7188 42800 7200
rect 22066 7160 41414 7188
rect 42755 7160 42800 7188
rect 12069 7151 12127 7157
rect 42794 7148 42800 7160
rect 42852 7148 42858 7200
rect 43162 7148 43168 7200
rect 43220 7188 43226 7200
rect 43257 7191 43315 7197
rect 43257 7188 43269 7191
rect 43220 7160 43269 7188
rect 43220 7148 43226 7160
rect 43257 7157 43269 7160
rect 43303 7157 43315 7191
rect 44008 7188 44036 7228
rect 44082 7216 44088 7268
rect 44140 7256 44146 7268
rect 45094 7256 45100 7268
rect 44140 7228 45100 7256
rect 44140 7216 44146 7228
rect 45094 7216 45100 7228
rect 45152 7216 45158 7268
rect 45186 7216 45192 7268
rect 45244 7256 45250 7268
rect 45281 7259 45339 7265
rect 45281 7256 45293 7259
rect 45244 7228 45293 7256
rect 45244 7216 45250 7228
rect 45281 7225 45293 7228
rect 45327 7225 45339 7259
rect 45281 7219 45339 7225
rect 45462 7216 45468 7268
rect 45520 7256 45526 7268
rect 46860 7256 46888 7355
rect 45520 7228 46888 7256
rect 45520 7216 45526 7228
rect 46014 7188 46020 7200
rect 44008 7160 46020 7188
rect 43257 7151 43315 7157
rect 46014 7148 46020 7160
rect 46072 7148 46078 7200
rect 47765 7191 47823 7197
rect 47765 7157 47777 7191
rect 47811 7188 47823 7191
rect 47854 7188 47860 7200
rect 47811 7160 47860 7188
rect 47811 7157 47823 7160
rect 47765 7151 47823 7157
rect 47854 7148 47860 7160
rect 47912 7148 47918 7200
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 3418 6944 3424 6996
rect 3476 6984 3482 6996
rect 14366 6984 14372 6996
rect 3476 6956 7880 6984
rect 3476 6944 3482 6956
rect 4172 6928 4200 6956
rect 566 6876 572 6928
rect 624 6916 630 6928
rect 3510 6916 3516 6928
rect 624 6888 3516 6916
rect 624 6876 630 6888
rect 3510 6876 3516 6888
rect 3568 6876 3574 6928
rect 4154 6876 4160 6928
rect 4212 6876 4218 6928
rect 4430 6876 4436 6928
rect 4488 6916 4494 6928
rect 4890 6916 4896 6928
rect 4488 6888 4896 6916
rect 4488 6876 4494 6888
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 2130 6848 2136 6860
rect 1412 6820 2136 6848
rect 474 6740 480 6792
rect 532 6780 538 6792
rect 1412 6789 1440 6820
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 2590 6808 2596 6860
rect 2648 6848 2654 6860
rect 7852 6848 7880 6956
rect 9646 6956 14372 6984
rect 9646 6916 9674 6956
rect 14366 6944 14372 6956
rect 14424 6944 14430 6996
rect 43809 6987 43867 6993
rect 43809 6953 43821 6987
rect 43855 6984 43867 6987
rect 43855 6956 45508 6984
rect 43855 6953 43867 6956
rect 43809 6947 43867 6953
rect 8680 6888 9674 6916
rect 10873 6919 10931 6925
rect 8680 6848 8708 6888
rect 10873 6885 10885 6919
rect 10919 6885 10931 6919
rect 44450 6916 44456 6928
rect 44411 6888 44456 6916
rect 10873 6879 10931 6885
rect 2648 6820 7788 6848
rect 7852 6820 8708 6848
rect 2648 6808 2654 6820
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 532 6752 1409 6780
rect 532 6740 538 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 2038 6780 2044 6792
rect 1999 6752 2044 6780
rect 1397 6743 1455 6749
rect 2038 6740 2044 6752
rect 2096 6740 2102 6792
rect 2314 6740 2320 6792
rect 2372 6780 2378 6792
rect 2685 6783 2743 6789
rect 2685 6780 2697 6783
rect 2372 6752 2697 6780
rect 2372 6740 2378 6752
rect 2685 6749 2697 6752
rect 2731 6782 2743 6783
rect 2731 6780 2820 6782
rect 3234 6780 3240 6792
rect 2731 6754 3240 6780
rect 2731 6749 2743 6754
rect 2792 6752 3240 6754
rect 2685 6743 2743 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 3844 6752 4077 6780
rect 3844 6740 3850 6752
rect 4065 6749 4077 6752
rect 4111 6780 4123 6783
rect 4430 6780 4436 6792
rect 4111 6752 4436 6780
rect 4111 6749 4123 6752
rect 4065 6743 4123 6749
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 4522 6740 4528 6792
rect 4580 6780 4586 6792
rect 4801 6783 4859 6789
rect 4801 6780 4813 6783
rect 4580 6752 4813 6780
rect 4580 6740 4586 6752
rect 4801 6749 4813 6752
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 5350 6740 5356 6792
rect 5408 6780 5414 6792
rect 5629 6783 5687 6789
rect 5408 6752 5580 6780
rect 5408 6740 5414 6752
rect 3418 6672 3424 6724
rect 3476 6712 3482 6724
rect 5552 6712 5580 6752
rect 5629 6749 5641 6783
rect 5675 6780 5687 6783
rect 5902 6780 5908 6792
rect 5675 6752 5908 6780
rect 5675 6749 5687 6752
rect 5629 6743 5687 6749
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 6178 6712 6184 6724
rect 3476 6684 5488 6712
rect 5552 6684 6184 6712
rect 3476 6672 3482 6684
rect 1394 6604 1400 6656
rect 1452 6644 1458 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1452 6616 1593 6644
rect 1452 6604 1458 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 2130 6644 2136 6656
rect 2091 6616 2136 6644
rect 1581 6607 1639 6613
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 2869 6647 2927 6653
rect 2869 6644 2881 6647
rect 2832 6616 2881 6644
rect 2832 6604 2838 6616
rect 2869 6613 2881 6616
rect 2915 6613 2927 6647
rect 2869 6607 2927 6613
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 3881 6647 3939 6653
rect 3881 6644 3893 6647
rect 3568 6616 3893 6644
rect 3568 6604 3574 6616
rect 3881 6613 3893 6616
rect 3927 6613 3939 6647
rect 3881 6607 3939 6613
rect 4617 6647 4675 6653
rect 4617 6613 4629 6647
rect 4663 6644 4675 6647
rect 4890 6644 4896 6656
rect 4663 6616 4896 6644
rect 4663 6613 4675 6616
rect 4617 6607 4675 6613
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 5460 6653 5488 6684
rect 6178 6672 6184 6684
rect 6236 6712 6242 6724
rect 6288 6712 6316 6743
rect 6236 6684 6316 6712
rect 6932 6712 6960 6743
rect 7190 6740 7196 6792
rect 7248 6780 7254 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7248 6752 7573 6780
rect 7248 6740 7254 6752
rect 7561 6749 7573 6752
rect 7607 6780 7619 6783
rect 7650 6780 7656 6792
rect 7607 6752 7656 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 7650 6740 7656 6752
rect 7708 6740 7714 6792
rect 7282 6712 7288 6724
rect 6932 6684 7288 6712
rect 6236 6672 6242 6684
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 7760 6712 7788 6820
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 10888 6848 10916 6879
rect 44450 6876 44456 6888
rect 44508 6876 44514 6928
rect 8812 6820 10916 6848
rect 8812 6808 8818 6820
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 44174 6848 44180 6860
rect 11020 6820 44180 6848
rect 11020 6808 11026 6820
rect 44174 6808 44180 6820
rect 44232 6808 44238 6860
rect 45370 6848 45376 6860
rect 44744 6820 45376 6848
rect 8202 6780 8208 6792
rect 8163 6752 8208 6780
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8904 6752 8953 6780
rect 8904 6740 8910 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6780 9827 6783
rect 9858 6780 9864 6792
rect 9815 6752 9864 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 10284 6752 10425 6780
rect 10284 6740 10290 6752
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10594 6740 10600 6792
rect 10652 6780 10658 6792
rect 11057 6783 11115 6789
rect 11057 6780 11069 6783
rect 10652 6752 11069 6780
rect 10652 6740 10658 6752
rect 11057 6749 11069 6752
rect 11103 6780 11115 6783
rect 11330 6780 11336 6792
rect 11103 6752 11336 6780
rect 11103 6749 11115 6752
rect 11057 6743 11115 6749
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 11606 6740 11612 6792
rect 11664 6780 11670 6792
rect 11701 6783 11759 6789
rect 11701 6780 11713 6783
rect 11664 6752 11713 6780
rect 11664 6740 11670 6752
rect 11701 6749 11713 6752
rect 11747 6780 11759 6783
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 11747 6752 12725 6780
rect 11747 6749 11759 6752
rect 11701 6743 11759 6749
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 13262 6780 13268 6792
rect 13223 6752 13268 6780
rect 12713 6743 12771 6749
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 42794 6740 42800 6792
rect 42852 6780 42858 6792
rect 44269 6783 44327 6789
rect 44269 6780 44281 6783
rect 42852 6752 44281 6780
rect 42852 6740 42858 6752
rect 44269 6749 44281 6752
rect 44315 6776 44327 6783
rect 44744 6780 44772 6820
rect 45370 6808 45376 6820
rect 45428 6808 45434 6860
rect 45480 6848 45508 6956
rect 47210 6848 47216 6860
rect 45480 6820 47216 6848
rect 47210 6808 47216 6820
rect 47268 6808 47274 6860
rect 47394 6848 47400 6860
rect 47355 6820 47400 6848
rect 47394 6808 47400 6820
rect 47452 6808 47458 6860
rect 44376 6776 44772 6780
rect 44315 6752 44772 6776
rect 44315 6749 44404 6752
rect 44269 6748 44404 6749
rect 44269 6743 44327 6748
rect 44818 6740 44824 6792
rect 44876 6780 44882 6792
rect 45005 6783 45063 6789
rect 45005 6780 45017 6783
rect 44876 6752 45017 6780
rect 44876 6740 44882 6752
rect 45005 6749 45017 6752
rect 45051 6749 45063 6783
rect 45646 6780 45652 6792
rect 45607 6752 45652 6780
rect 45005 6743 45063 6749
rect 45646 6740 45652 6752
rect 45704 6740 45710 6792
rect 46477 6783 46535 6789
rect 46477 6749 46489 6783
rect 46523 6749 46535 6783
rect 46477 6743 46535 6749
rect 43254 6712 43260 6724
rect 7760 6684 12434 6712
rect 43215 6684 43260 6712
rect 5445 6647 5503 6653
rect 5445 6613 5457 6647
rect 5491 6613 5503 6647
rect 5445 6607 5503 6613
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 6089 6647 6147 6653
rect 6089 6644 6101 6647
rect 5592 6616 6101 6644
rect 5592 6604 5598 6616
rect 6089 6613 6101 6616
rect 6135 6613 6147 6647
rect 6089 6607 6147 6613
rect 6454 6604 6460 6656
rect 6512 6644 6518 6656
rect 6733 6647 6791 6653
rect 6733 6644 6745 6647
rect 6512 6616 6745 6644
rect 6512 6604 6518 6616
rect 6733 6613 6745 6616
rect 6779 6613 6791 6647
rect 6733 6607 6791 6613
rect 7098 6604 7104 6656
rect 7156 6644 7162 6656
rect 7377 6647 7435 6653
rect 7377 6644 7389 6647
rect 7156 6616 7389 6644
rect 7156 6604 7162 6616
rect 7377 6613 7389 6616
rect 7423 6613 7435 6647
rect 7377 6607 7435 6613
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 8021 6647 8079 6653
rect 8021 6644 8033 6647
rect 7984 6616 8033 6644
rect 7984 6604 7990 6616
rect 8021 6613 8033 6616
rect 8067 6613 8079 6647
rect 9030 6644 9036 6656
rect 8991 6616 9036 6644
rect 8021 6607 8079 6613
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 9122 6604 9128 6656
rect 9180 6644 9186 6656
rect 9585 6647 9643 6653
rect 9585 6644 9597 6647
rect 9180 6616 9597 6644
rect 9180 6604 9186 6616
rect 9585 6613 9597 6616
rect 9631 6613 9643 6647
rect 9585 6607 9643 6613
rect 10229 6647 10287 6653
rect 10229 6613 10241 6647
rect 10275 6644 10287 6647
rect 10410 6644 10416 6656
rect 10275 6616 10416 6644
rect 10275 6613 10287 6616
rect 10229 6607 10287 6613
rect 10410 6604 10416 6616
rect 10468 6604 10474 6656
rect 11514 6644 11520 6656
rect 11475 6616 11520 6644
rect 11514 6604 11520 6616
rect 11572 6604 11578 6656
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 12161 6647 12219 6653
rect 12161 6644 12173 6647
rect 11848 6616 12173 6644
rect 11848 6604 11854 6616
rect 12161 6613 12173 6616
rect 12207 6613 12219 6647
rect 12406 6644 12434 6684
rect 43254 6672 43260 6684
rect 43312 6672 43318 6724
rect 45664 6712 45692 6740
rect 44376 6684 45692 6712
rect 17034 6644 17040 6656
rect 12406 6616 17040 6644
rect 12161 6607 12219 6613
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 42705 6647 42763 6653
rect 42705 6613 42717 6647
rect 42751 6644 42763 6647
rect 44376 6644 44404 6684
rect 42751 6616 44404 6644
rect 45189 6647 45247 6653
rect 42751 6613 42763 6616
rect 42705 6607 42763 6613
rect 45189 6613 45201 6647
rect 45235 6644 45247 6647
rect 45738 6644 45744 6656
rect 45235 6616 45744 6644
rect 45235 6613 45247 6616
rect 45189 6607 45247 6613
rect 45738 6604 45744 6616
rect 45796 6604 45802 6656
rect 45833 6647 45891 6653
rect 45833 6613 45845 6647
rect 45879 6644 45891 6647
rect 46290 6644 46296 6656
rect 45879 6616 46296 6644
rect 45879 6613 45891 6616
rect 45833 6607 45891 6613
rect 46290 6604 46296 6616
rect 46348 6604 46354 6656
rect 46492 6644 46520 6743
rect 46750 6740 46756 6792
rect 46808 6780 46814 6792
rect 47581 6783 47639 6789
rect 47581 6780 47593 6783
rect 46808 6752 47593 6780
rect 46808 6740 46814 6752
rect 47581 6749 47593 6752
rect 47627 6749 47639 6783
rect 47581 6743 47639 6749
rect 47670 6740 47676 6792
rect 47728 6780 47734 6792
rect 47949 6783 48007 6789
rect 47949 6780 47961 6783
rect 47728 6752 47961 6780
rect 47728 6740 47734 6752
rect 47949 6749 47961 6752
rect 47995 6749 48007 6783
rect 47949 6743 48007 6749
rect 48038 6740 48044 6792
rect 48096 6780 48102 6792
rect 48096 6752 48141 6780
rect 48096 6740 48102 6752
rect 46934 6712 46940 6724
rect 46895 6684 46940 6712
rect 46934 6672 46940 6684
rect 46992 6672 46998 6724
rect 48961 6647 49019 6653
rect 48961 6644 48973 6647
rect 46492 6616 48973 6644
rect 48961 6613 48973 6616
rect 49007 6613 49019 6647
rect 48961 6607 49019 6613
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 2038 6400 2044 6452
rect 2096 6440 2102 6452
rect 2406 6440 2412 6452
rect 2096 6412 2412 6440
rect 2096 6400 2102 6412
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 3329 6443 3387 6449
rect 2556 6412 3188 6440
rect 2556 6400 2562 6412
rect 3160 6372 3188 6412
rect 3329 6409 3341 6443
rect 3375 6409 3387 6443
rect 5721 6443 5779 6449
rect 5721 6440 5733 6443
rect 3329 6403 3387 6409
rect 3436 6412 5733 6440
rect 3344 6372 3372 6403
rect 3160 6344 3372 6372
rect 1854 6264 1860 6316
rect 1912 6304 1918 6316
rect 1949 6307 2007 6313
rect 1949 6304 1961 6307
rect 1912 6276 1961 6304
rect 1912 6264 1918 6276
rect 1949 6273 1961 6276
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6273 2835 6307
rect 2777 6267 2835 6273
rect 1578 6196 1584 6248
rect 1636 6236 1642 6248
rect 1636 6208 1900 6236
rect 1636 6196 1642 6208
rect 1872 6180 1900 6208
rect 1854 6128 1860 6180
rect 1912 6128 1918 6180
rect 1964 6168 1992 6267
rect 2792 6236 2820 6267
rect 3234 6264 3240 6316
rect 3292 6304 3298 6316
rect 3436 6304 3464 6412
rect 5721 6409 5733 6412
rect 5767 6409 5779 6443
rect 5721 6403 5779 6409
rect 4338 6372 4344 6384
rect 3528 6344 4344 6372
rect 3528 6313 3556 6344
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 4522 6332 4528 6384
rect 4580 6372 4586 6384
rect 5736 6372 5764 6403
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 9677 6443 9735 6449
rect 9677 6440 9689 6443
rect 8168 6412 9689 6440
rect 8168 6400 8174 6412
rect 9677 6409 9689 6412
rect 9723 6409 9735 6443
rect 9677 6403 9735 6409
rect 11422 6400 11428 6452
rect 11480 6440 11486 6452
rect 23014 6440 23020 6452
rect 11480 6412 23020 6440
rect 11480 6400 11486 6412
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 43257 6443 43315 6449
rect 43257 6409 43269 6443
rect 43303 6440 43315 6443
rect 44082 6440 44088 6452
rect 43303 6412 44088 6440
rect 43303 6409 43315 6412
rect 43257 6403 43315 6409
rect 44082 6400 44088 6412
rect 44140 6400 44146 6452
rect 44266 6400 44272 6452
rect 44324 6440 44330 6452
rect 45462 6440 45468 6452
rect 44324 6412 45468 6440
rect 44324 6400 44330 6412
rect 45462 6400 45468 6412
rect 45520 6400 45526 6452
rect 45922 6440 45928 6452
rect 45883 6412 45928 6440
rect 45922 6400 45928 6412
rect 45980 6400 45986 6452
rect 47765 6443 47823 6449
rect 47765 6409 47777 6443
rect 47811 6440 47823 6443
rect 48038 6440 48044 6452
rect 47811 6412 48044 6440
rect 47811 6409 47823 6412
rect 47765 6403 47823 6409
rect 8478 6372 8484 6384
rect 4580 6344 5212 6372
rect 5736 6344 8484 6372
rect 4580 6332 4586 6344
rect 3292 6276 3464 6304
rect 3513 6307 3571 6313
rect 3292 6264 3298 6276
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 4246 6304 4252 6316
rect 4207 6276 4252 6304
rect 3513 6267 3571 6273
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4798 6264 4804 6316
rect 4856 6304 4862 6316
rect 4985 6307 5043 6313
rect 4985 6304 4997 6307
rect 4856 6276 4997 6304
rect 4856 6264 4862 6276
rect 4985 6273 4997 6276
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 4154 6236 4160 6248
rect 2792 6208 4160 6236
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 5184 6236 5212 6344
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 11054 6372 11060 6384
rect 8588 6344 11060 6372
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 5718 6304 5724 6316
rect 5675 6276 5724 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 7006 6304 7012 6316
rect 6687 6276 7012 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 7374 6304 7380 6316
rect 7335 6276 7380 6304
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6304 8171 6307
rect 8386 6304 8392 6316
rect 8159 6276 8392 6304
rect 8159 6273 8171 6276
rect 8113 6267 8171 6273
rect 8386 6264 8392 6276
rect 8444 6264 8450 6316
rect 5442 6236 5448 6248
rect 5184 6208 5448 6236
rect 5442 6196 5448 6208
rect 5500 6236 5506 6248
rect 8588 6236 8616 6344
rect 11054 6332 11060 6344
rect 11112 6332 11118 6384
rect 13998 6372 14004 6384
rect 13959 6344 14004 6372
rect 13998 6332 14004 6344
rect 14056 6332 14062 6384
rect 14550 6372 14556 6384
rect 14511 6344 14556 6372
rect 14550 6332 14556 6344
rect 14608 6332 14614 6384
rect 44450 6332 44456 6384
rect 44508 6372 44514 6384
rect 47780 6372 47808 6403
rect 48038 6400 48044 6412
rect 48096 6400 48102 6452
rect 44508 6344 46520 6372
rect 44508 6332 44514 6344
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6304 9275 6307
rect 9674 6304 9680 6316
rect 9263 6276 9680 6304
rect 9263 6273 9275 6276
rect 9217 6267 9275 6273
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 9861 6307 9919 6313
rect 9861 6273 9873 6307
rect 9907 6304 9919 6307
rect 10134 6304 10140 6316
rect 9907 6276 10140 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10505 6307 10563 6313
rect 10505 6273 10517 6307
rect 10551 6304 10563 6307
rect 10778 6304 10784 6316
rect 10551 6276 10784 6304
rect 10551 6273 10563 6276
rect 10505 6267 10563 6273
rect 5500 6208 8616 6236
rect 5500 6196 5506 6208
rect 9398 6196 9404 6248
rect 9456 6236 9462 6248
rect 10520 6236 10548 6267
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 11238 6264 11244 6316
rect 11296 6304 11302 6316
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 11296 6276 11989 6304
rect 11296 6264 11302 6276
rect 11977 6273 11989 6276
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 17218 6264 17224 6316
rect 17276 6304 17282 6316
rect 23658 6304 23664 6316
rect 17276 6276 23664 6304
rect 17276 6264 17282 6276
rect 23658 6264 23664 6276
rect 23716 6264 23722 6316
rect 41877 6307 41935 6313
rect 41877 6273 41889 6307
rect 41923 6304 41935 6307
rect 43717 6307 43775 6313
rect 43717 6304 43729 6307
rect 41923 6276 43729 6304
rect 41923 6273 41935 6276
rect 41877 6267 41935 6273
rect 43717 6273 43729 6276
rect 43763 6273 43775 6307
rect 43717 6267 43775 6273
rect 44361 6307 44419 6313
rect 44361 6273 44373 6307
rect 44407 6304 44419 6307
rect 44542 6304 44548 6316
rect 44407 6276 44548 6304
rect 44407 6273 44419 6276
rect 44361 6267 44419 6273
rect 12250 6236 12256 6248
rect 9456 6208 10548 6236
rect 12211 6208 12256 6236
rect 9456 6196 9462 6208
rect 12250 6196 12256 6208
rect 12308 6196 12314 6248
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 39298 6236 39304 6248
rect 14424 6208 39304 6236
rect 14424 6196 14430 6208
rect 39298 6196 39304 6208
rect 39356 6196 39362 6248
rect 43162 6236 43168 6248
rect 41386 6208 43168 6236
rect 10962 6168 10968 6180
rect 1964 6140 10968 6168
rect 10962 6128 10968 6140
rect 11020 6128 11026 6180
rect 11330 6128 11336 6180
rect 11388 6168 11394 6180
rect 41386 6168 41414 6208
rect 43162 6196 43168 6208
rect 43220 6196 43226 6248
rect 43732 6236 43760 6267
rect 44542 6264 44548 6276
rect 44600 6304 44606 6316
rect 44910 6304 44916 6316
rect 44600 6276 44916 6304
rect 44600 6264 44606 6276
rect 44910 6264 44916 6276
rect 44968 6264 44974 6316
rect 45186 6304 45192 6316
rect 45147 6276 45192 6304
rect 45186 6264 45192 6276
rect 45244 6264 45250 6316
rect 46492 6313 46520 6344
rect 47044 6344 47808 6372
rect 46477 6307 46535 6313
rect 46477 6273 46489 6307
rect 46523 6273 46535 6307
rect 46842 6304 46848 6316
rect 46803 6276 46848 6304
rect 46477 6267 46535 6273
rect 46842 6264 46848 6276
rect 46900 6264 46906 6316
rect 47044 6313 47072 6344
rect 47029 6307 47087 6313
rect 47029 6273 47041 6307
rect 47075 6273 47087 6307
rect 47029 6267 47087 6273
rect 47486 6264 47492 6316
rect 47544 6304 47550 6316
rect 47581 6307 47639 6313
rect 47581 6304 47593 6307
rect 47544 6276 47593 6304
rect 47544 6264 47550 6276
rect 47581 6273 47593 6276
rect 47627 6273 47639 6307
rect 47581 6267 47639 6273
rect 45554 6236 45560 6248
rect 43732 6208 45560 6236
rect 45554 6196 45560 6208
rect 45612 6196 45618 6248
rect 46569 6239 46627 6245
rect 46569 6205 46581 6239
rect 46615 6205 46627 6239
rect 46569 6199 46627 6205
rect 11388 6140 41414 6168
rect 42705 6171 42763 6177
rect 11388 6128 11394 6140
rect 42705 6137 42717 6171
rect 42751 6168 42763 6171
rect 43254 6168 43260 6180
rect 42751 6140 43260 6168
rect 42751 6137 42763 6140
rect 42705 6131 42763 6137
rect 43254 6128 43260 6140
rect 43312 6128 43318 6180
rect 43901 6171 43959 6177
rect 43901 6137 43913 6171
rect 43947 6168 43959 6171
rect 46584 6168 46612 6199
rect 47394 6168 47400 6180
rect 43947 6140 45784 6168
rect 46584 6140 47400 6168
rect 43947 6137 43959 6140
rect 43901 6131 43959 6137
rect 753 6103 811 6109
rect 753 6069 765 6103
rect 799 6100 811 6103
rect 1118 6100 1124 6112
rect 799 6072 1124 6100
rect 799 6069 811 6072
rect 753 6063 811 6069
rect 1118 6060 1124 6072
rect 1176 6060 1182 6112
rect 1578 6060 1584 6112
rect 1636 6100 1642 6112
rect 1765 6103 1823 6109
rect 1765 6100 1777 6103
rect 1636 6072 1777 6100
rect 1636 6060 1642 6072
rect 1765 6069 1777 6072
rect 1811 6069 1823 6103
rect 1765 6063 1823 6069
rect 2406 6060 2412 6112
rect 2464 6100 2470 6112
rect 2593 6103 2651 6109
rect 2593 6100 2605 6103
rect 2464 6072 2605 6100
rect 2464 6060 2470 6072
rect 2593 6069 2605 6072
rect 2639 6069 2651 6103
rect 2593 6063 2651 6069
rect 3786 6060 3792 6112
rect 3844 6100 3850 6112
rect 4065 6103 4123 6109
rect 4065 6100 4077 6103
rect 3844 6072 4077 6100
rect 3844 6060 3850 6072
rect 4065 6069 4077 6072
rect 4111 6069 4123 6103
rect 4065 6063 4123 6069
rect 4801 6103 4859 6109
rect 4801 6069 4813 6103
rect 4847 6100 4859 6103
rect 5074 6100 5080 6112
rect 4847 6072 5080 6100
rect 4847 6069 4859 6072
rect 4801 6063 4859 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 6178 6100 6184 6112
rect 5776 6072 6184 6100
rect 5776 6060 5782 6072
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 6270 6060 6276 6112
rect 6328 6100 6334 6112
rect 6457 6103 6515 6109
rect 6457 6100 6469 6103
rect 6328 6072 6469 6100
rect 6328 6060 6334 6072
rect 6457 6069 6469 6072
rect 6503 6069 6515 6103
rect 6457 6063 6515 6069
rect 7006 6060 7012 6112
rect 7064 6100 7070 6112
rect 7193 6103 7251 6109
rect 7193 6100 7205 6103
rect 7064 6072 7205 6100
rect 7064 6060 7070 6072
rect 7193 6069 7205 6072
rect 7239 6069 7251 6103
rect 7193 6063 7251 6069
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 7929 6103 7987 6109
rect 7929 6100 7941 6103
rect 7616 6072 7941 6100
rect 7616 6060 7622 6072
rect 7929 6069 7941 6072
rect 7975 6069 7987 6103
rect 7929 6063 7987 6069
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 8386 6100 8392 6112
rect 8260 6072 8392 6100
rect 8260 6060 8266 6072
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 9030 6100 9036 6112
rect 8991 6072 9036 6100
rect 9030 6060 9036 6072
rect 9088 6060 9094 6112
rect 10318 6100 10324 6112
rect 10279 6072 10324 6100
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 12526 6060 12532 6112
rect 12584 6100 12590 6112
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 12584 6072 12909 6100
rect 12584 6060 12590 6072
rect 12897 6069 12909 6072
rect 12943 6069 12955 6103
rect 12897 6063 12955 6069
rect 13078 6060 13084 6112
rect 13136 6100 13142 6112
rect 13449 6103 13507 6109
rect 13449 6100 13461 6103
rect 13136 6072 13461 6100
rect 13136 6060 13142 6072
rect 13449 6069 13461 6072
rect 13495 6069 13507 6103
rect 15194 6100 15200 6112
rect 15155 6072 15200 6100
rect 13449 6063 13507 6069
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 44542 6100 44548 6112
rect 44503 6072 44548 6100
rect 44542 6060 44548 6072
rect 44600 6060 44606 6112
rect 45094 6100 45100 6112
rect 45055 6072 45100 6100
rect 45094 6060 45100 6072
rect 45152 6060 45158 6112
rect 45756 6100 45784 6140
rect 47394 6128 47400 6140
rect 47452 6128 47458 6180
rect 47578 6100 47584 6112
rect 45756 6072 47584 6100
rect 47578 6060 47584 6072
rect 47636 6060 47642 6112
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 1026 5856 1032 5908
rect 1084 5896 1090 5908
rect 2130 5896 2136 5908
rect 1084 5868 2136 5896
rect 1084 5856 1090 5868
rect 2130 5856 2136 5868
rect 2188 5896 2194 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 2188 5868 4077 5896
rect 2188 5856 2194 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 7374 5896 7380 5908
rect 4065 5859 4123 5865
rect 6472 5868 6868 5896
rect 7335 5868 7380 5896
rect 1118 5788 1124 5840
rect 1176 5828 1182 5840
rect 2225 5831 2283 5837
rect 2225 5828 2237 5831
rect 1176 5800 2237 5828
rect 1176 5788 1182 5800
rect 2225 5797 2237 5800
rect 2271 5797 2283 5831
rect 2225 5791 2283 5797
rect 2332 5800 6224 5828
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1673 5695 1731 5701
rect 1673 5692 1685 5695
rect 1544 5664 1685 5692
rect 1544 5652 1550 5664
rect 1673 5661 1685 5664
rect 1719 5692 1731 5695
rect 2332 5692 2360 5800
rect 4154 5760 4160 5772
rect 4115 5732 4160 5760
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 5442 5720 5448 5772
rect 5500 5720 5506 5772
rect 6196 5760 6224 5800
rect 6472 5760 6500 5868
rect 6730 5788 6736 5840
rect 6788 5788 6794 5840
rect 6840 5828 6868 5868
rect 7374 5856 7380 5868
rect 7432 5896 7438 5908
rect 8110 5896 8116 5908
rect 7432 5868 8116 5896
rect 7432 5856 7438 5868
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8260 5868 9045 5896
rect 8260 5856 8266 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 9306 5856 9312 5908
rect 9364 5896 9370 5908
rect 10226 5896 10232 5908
rect 9364 5868 10232 5896
rect 9364 5856 9370 5868
rect 10226 5856 10232 5868
rect 10284 5856 10290 5908
rect 12250 5856 12256 5908
rect 12308 5896 12314 5908
rect 14737 5899 14795 5905
rect 14737 5896 14749 5899
rect 12308 5868 14749 5896
rect 12308 5856 12314 5868
rect 14737 5865 14749 5868
rect 14783 5896 14795 5899
rect 15286 5896 15292 5908
rect 14783 5868 15292 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 15838 5896 15844 5908
rect 15799 5868 15844 5896
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 43809 5899 43867 5905
rect 43809 5865 43821 5899
rect 43855 5896 43867 5899
rect 46385 5899 46443 5905
rect 43855 5868 46244 5896
rect 43855 5865 43867 5868
rect 43809 5859 43867 5865
rect 45002 5828 45008 5840
rect 6840 5800 45008 5828
rect 45002 5788 45008 5800
rect 45060 5788 45066 5840
rect 45186 5788 45192 5840
rect 45244 5828 45250 5840
rect 46109 5831 46167 5837
rect 46109 5828 46121 5831
rect 45244 5800 46121 5828
rect 45244 5788 45250 5800
rect 46109 5797 46121 5800
rect 46155 5797 46167 5831
rect 46216 5828 46244 5868
rect 46385 5865 46397 5899
rect 46431 5896 46443 5899
rect 47394 5896 47400 5908
rect 46431 5868 47400 5896
rect 46431 5865 46443 5868
rect 46385 5859 46443 5865
rect 47394 5856 47400 5868
rect 47452 5856 47458 5908
rect 46750 5828 46756 5840
rect 46216 5800 46756 5828
rect 46109 5791 46167 5797
rect 46750 5788 46756 5800
rect 46808 5788 46814 5840
rect 47210 5828 47216 5840
rect 47171 5800 47216 5828
rect 47210 5788 47216 5800
rect 47268 5788 47274 5840
rect 47302 5788 47308 5840
rect 47360 5828 47366 5840
rect 47360 5800 47992 5828
rect 47360 5788 47366 5800
rect 6196 5732 6500 5760
rect 1719 5664 2360 5692
rect 2409 5695 2467 5701
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 2409 5661 2421 5695
rect 2455 5692 2467 5695
rect 2590 5692 2596 5704
rect 2455 5664 2596 5692
rect 2455 5661 2467 5664
rect 2409 5655 2467 5661
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5692 3203 5695
rect 4246 5692 4252 5704
rect 3191 5664 4252 5692
rect 3191 5661 3203 5664
rect 3145 5655 3203 5661
rect 4246 5652 4252 5664
rect 4304 5652 4310 5704
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5692 5135 5695
rect 5460 5692 5488 5720
rect 5123 5664 5488 5692
rect 5123 5661 5135 5664
rect 5077 5655 5135 5661
rect 5718 5652 5724 5704
rect 5776 5692 5782 5704
rect 5813 5695 5871 5701
rect 5813 5692 5825 5695
rect 5776 5664 5825 5692
rect 5776 5652 5782 5664
rect 5813 5661 5825 5664
rect 5859 5661 5871 5695
rect 5813 5655 5871 5661
rect 6178 5652 6184 5704
rect 6236 5692 6242 5704
rect 6561 5695 6619 5701
rect 6236 5664 6500 5692
rect 6236 5652 6242 5664
rect 2130 5584 2136 5636
rect 2188 5624 2194 5636
rect 2188 5596 3188 5624
rect 2188 5584 2194 5596
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2958 5556 2964 5568
rect 2919 5528 2964 5556
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 3160 5556 3188 5596
rect 3234 5584 3240 5636
rect 3292 5624 3298 5636
rect 3973 5627 4031 5633
rect 3973 5624 3985 5627
rect 3292 5596 3985 5624
rect 3292 5584 3298 5596
rect 3973 5593 3985 5596
rect 4019 5593 4031 5627
rect 4341 5627 4399 5633
rect 4341 5624 4353 5627
rect 3973 5587 4031 5593
rect 4172 5596 4353 5624
rect 4172 5568 4200 5596
rect 4341 5593 4353 5596
rect 4387 5593 4399 5627
rect 4341 5587 4399 5593
rect 5442 5584 5448 5636
rect 5500 5624 5506 5636
rect 6472 5624 6500 5664
rect 6561 5661 6573 5695
rect 6607 5692 6619 5695
rect 6748 5692 6776 5788
rect 10962 5760 10968 5772
rect 8404 5732 10968 5760
rect 6607 5664 6776 5692
rect 6607 5661 6619 5664
rect 6561 5655 6619 5661
rect 6822 5652 6828 5704
rect 6880 5692 6886 5704
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 6880 5664 7297 5692
rect 6880 5652 6886 5664
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 7469 5695 7527 5701
rect 7469 5692 7481 5695
rect 7432 5664 7481 5692
rect 7432 5652 7438 5664
rect 7469 5661 7481 5664
rect 7515 5692 7527 5695
rect 8110 5692 8116 5704
rect 7515 5664 8116 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 8404 5701 8432 5732
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 12434 5760 12440 5772
rect 11348 5732 12440 5760
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5661 8447 5695
rect 9214 5692 9220 5704
rect 9175 5664 9220 5692
rect 8389 5655 8447 5661
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9674 5692 9680 5704
rect 9635 5664 9680 5692
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5692 10011 5695
rect 10042 5692 10048 5704
rect 9999 5664 10048 5692
rect 9999 5661 10011 5664
rect 9953 5655 10011 5661
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10873 5695 10931 5701
rect 10873 5692 10885 5695
rect 10284 5664 10885 5692
rect 10284 5652 10290 5664
rect 10873 5661 10885 5664
rect 10919 5692 10931 5695
rect 11348 5692 11376 5732
rect 12434 5720 12440 5732
rect 12492 5720 12498 5772
rect 14274 5720 14280 5772
rect 14332 5760 14338 5772
rect 15194 5760 15200 5772
rect 14332 5732 15200 5760
rect 14332 5720 14338 5732
rect 15194 5720 15200 5732
rect 15252 5760 15258 5772
rect 44450 5760 44456 5772
rect 15252 5732 44456 5760
rect 15252 5720 15258 5732
rect 44450 5720 44456 5732
rect 44508 5720 44514 5772
rect 44542 5720 44548 5772
rect 44600 5760 44606 5772
rect 44600 5732 47624 5760
rect 44600 5720 44606 5732
rect 11698 5692 11704 5704
rect 10919 5664 11376 5692
rect 11659 5664 11704 5692
rect 10919 5661 10931 5664
rect 10873 5655 10931 5661
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 17218 5692 17224 5704
rect 12032 5664 17224 5692
rect 12032 5652 12038 5664
rect 17218 5652 17224 5664
rect 17276 5652 17282 5704
rect 41509 5695 41567 5701
rect 41509 5661 41521 5695
rect 41555 5692 41567 5695
rect 43622 5692 43628 5704
rect 41555 5664 43628 5692
rect 41555 5661 41567 5664
rect 41509 5655 41567 5661
rect 43622 5652 43628 5664
rect 43680 5692 43686 5704
rect 43680 5664 43725 5692
rect 43680 5652 43686 5664
rect 44082 5652 44088 5704
rect 44140 5692 44146 5704
rect 44269 5695 44327 5701
rect 44269 5692 44281 5695
rect 44140 5664 44281 5692
rect 44140 5652 44146 5664
rect 44269 5661 44281 5664
rect 44315 5661 44327 5695
rect 44269 5655 44327 5661
rect 45373 5695 45431 5701
rect 45373 5661 45385 5695
rect 45419 5692 45431 5695
rect 45830 5692 45836 5704
rect 45419 5664 45836 5692
rect 45419 5661 45431 5664
rect 45373 5655 45431 5661
rect 45830 5652 45836 5664
rect 45888 5652 45894 5704
rect 46109 5695 46167 5701
rect 46109 5661 46121 5695
rect 46155 5692 46167 5695
rect 46201 5695 46259 5701
rect 46201 5692 46213 5695
rect 46155 5664 46213 5692
rect 46155 5661 46167 5664
rect 46109 5655 46167 5661
rect 46201 5661 46213 5664
rect 46247 5661 46259 5695
rect 47394 5692 47400 5704
rect 47355 5664 47400 5692
rect 46201 5655 46259 5661
rect 47394 5652 47400 5664
rect 47452 5652 47458 5704
rect 47596 5701 47624 5732
rect 47964 5701 47992 5800
rect 47581 5695 47639 5701
rect 47581 5661 47593 5695
rect 47627 5661 47639 5695
rect 47581 5655 47639 5661
rect 47949 5695 48007 5701
rect 47949 5661 47961 5695
rect 47995 5661 48007 5695
rect 47949 5655 48007 5661
rect 48038 5652 48044 5704
rect 48096 5692 48102 5704
rect 48096 5664 48141 5692
rect 48096 5652 48102 5664
rect 5500 5596 5856 5624
rect 6472 5596 9674 5624
rect 5500 5584 5506 5596
rect 4154 5556 4160 5568
rect 3160 5528 4160 5556
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 4249 5559 4307 5565
rect 4249 5525 4261 5559
rect 4295 5556 4307 5559
rect 4614 5556 4620 5568
rect 4295 5528 4620 5556
rect 4295 5525 4307 5528
rect 4249 5519 4307 5525
rect 4614 5516 4620 5528
rect 4672 5516 4678 5568
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 4893 5559 4951 5565
rect 4893 5556 4905 5559
rect 4856 5528 4905 5556
rect 4856 5516 4862 5528
rect 4893 5525 4905 5528
rect 4939 5525 4951 5559
rect 4893 5519 4951 5525
rect 5629 5559 5687 5565
rect 5629 5525 5641 5559
rect 5675 5556 5687 5559
rect 5718 5556 5724 5568
rect 5675 5528 5724 5556
rect 5675 5525 5687 5528
rect 5629 5519 5687 5525
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 5828 5556 5856 5596
rect 6365 5559 6423 5565
rect 6365 5556 6377 5559
rect 5828 5528 6377 5556
rect 6365 5525 6377 5528
rect 6411 5525 6423 5559
rect 6365 5519 6423 5525
rect 7653 5559 7711 5565
rect 7653 5525 7665 5559
rect 7699 5556 7711 5559
rect 8110 5556 8116 5568
rect 7699 5528 8116 5556
rect 7699 5525 7711 5528
rect 7653 5519 7711 5525
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 8205 5559 8263 5565
rect 8205 5525 8217 5559
rect 8251 5556 8263 5559
rect 8294 5556 8300 5568
rect 8251 5528 8300 5556
rect 8251 5525 8263 5528
rect 8205 5519 8263 5525
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 9646 5556 9674 5596
rect 10594 5584 10600 5636
rect 10652 5624 10658 5636
rect 11057 5627 11115 5633
rect 11057 5624 11069 5627
rect 10652 5596 11069 5624
rect 10652 5584 10658 5596
rect 11057 5593 11069 5596
rect 11103 5593 11115 5627
rect 11238 5624 11244 5636
rect 11199 5596 11244 5624
rect 11057 5587 11115 5593
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 14366 5624 14372 5636
rect 11348 5596 14372 5624
rect 11348 5556 11376 5596
rect 14366 5584 14372 5596
rect 14424 5584 14430 5636
rect 45593 5627 45651 5633
rect 45593 5593 45605 5627
rect 45639 5624 45651 5627
rect 47486 5624 47492 5636
rect 45639 5596 47492 5624
rect 45639 5593 45651 5596
rect 45593 5587 45651 5593
rect 47486 5584 47492 5596
rect 47544 5584 47550 5636
rect 9646 5528 11376 5556
rect 11885 5559 11943 5565
rect 11885 5525 11897 5559
rect 11931 5556 11943 5559
rect 12250 5556 12256 5568
rect 11931 5528 12256 5556
rect 11931 5525 11943 5528
rect 11885 5519 11943 5525
rect 12250 5516 12256 5528
rect 12308 5516 12314 5568
rect 12894 5556 12900 5568
rect 12855 5528 12900 5556
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 12986 5516 12992 5568
rect 13044 5556 13050 5568
rect 13449 5559 13507 5565
rect 13449 5556 13461 5559
rect 13044 5528 13461 5556
rect 13044 5516 13050 5528
rect 13449 5525 13461 5528
rect 13495 5525 13507 5559
rect 13449 5519 13507 5525
rect 13630 5516 13636 5568
rect 13688 5556 13694 5568
rect 14093 5559 14151 5565
rect 14093 5556 14105 5559
rect 13688 5528 14105 5556
rect 13688 5516 13694 5528
rect 14093 5525 14105 5528
rect 14139 5525 14151 5559
rect 14093 5519 14151 5525
rect 15197 5559 15255 5565
rect 15197 5525 15209 5559
rect 15243 5556 15255 5559
rect 15378 5556 15384 5568
rect 15243 5528 15384 5556
rect 15243 5525 15255 5528
rect 15197 5519 15255 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 42058 5556 42064 5568
rect 42019 5528 42064 5556
rect 42058 5516 42064 5528
rect 42116 5516 42122 5568
rect 42610 5556 42616 5568
rect 42571 5528 42616 5556
rect 42610 5516 42616 5528
rect 42668 5516 42674 5568
rect 43165 5559 43223 5565
rect 43165 5525 43177 5559
rect 43211 5556 43223 5559
rect 44266 5556 44272 5568
rect 43211 5528 44272 5556
rect 43211 5525 43223 5528
rect 43165 5519 43223 5525
rect 44266 5516 44272 5528
rect 44324 5516 44330 5568
rect 44453 5559 44511 5565
rect 44453 5525 44465 5559
rect 44499 5556 44511 5559
rect 45186 5556 45192 5568
rect 44499 5528 45192 5556
rect 44499 5525 44511 5528
rect 44453 5519 44511 5525
rect 45186 5516 45192 5528
rect 45244 5516 45250 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 2869 5355 2927 5361
rect 2869 5352 2881 5355
rect 2746 5324 2881 5352
rect 1302 5244 1308 5296
rect 1360 5284 1366 5296
rect 2746 5284 2774 5324
rect 2869 5321 2881 5324
rect 2915 5321 2927 5355
rect 2869 5315 2927 5321
rect 3234 5312 3240 5364
rect 3292 5352 3298 5364
rect 3602 5352 3608 5364
rect 3292 5324 3608 5352
rect 3292 5312 3298 5324
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 6914 5352 6920 5364
rect 6104 5324 6920 5352
rect 3694 5284 3700 5296
rect 1360 5256 2774 5284
rect 3655 5256 3700 5284
rect 1360 5244 1366 5256
rect 3694 5244 3700 5256
rect 3752 5244 3758 5296
rect 4154 5244 4160 5296
rect 4212 5284 4218 5296
rect 4522 5284 4528 5296
rect 4212 5256 4528 5284
rect 4212 5244 4218 5256
rect 4522 5244 4528 5256
rect 4580 5284 4586 5296
rect 4617 5287 4675 5293
rect 4617 5284 4629 5287
rect 4580 5256 4629 5284
rect 4580 5244 4586 5256
rect 4617 5253 4629 5256
rect 4663 5253 4675 5287
rect 4617 5247 4675 5253
rect 1210 5176 1216 5228
rect 1268 5176 1274 5228
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 2130 5216 2136 5228
rect 1719 5188 2136 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5216 2835 5219
rect 2866 5216 2872 5228
rect 2823 5188 2872 5216
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 5721 5219 5779 5225
rect 5721 5185 5733 5219
rect 5767 5216 5779 5219
rect 6104 5216 6132 5324
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 7650 5352 7656 5364
rect 7576 5324 7656 5352
rect 7282 5284 7288 5296
rect 6748 5256 7288 5284
rect 6748 5225 6776 5256
rect 7282 5244 7288 5256
rect 7340 5244 7346 5296
rect 5767 5188 6132 5216
rect 6733 5219 6791 5225
rect 5767 5185 5779 5188
rect 5721 5179 5779 5185
rect 6733 5185 6745 5219
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 1228 5080 1256 5176
rect 3694 5108 3700 5160
rect 3752 5148 3758 5160
rect 4062 5148 4068 5160
rect 3752 5120 4068 5148
rect 3752 5108 3758 5120
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 6178 5108 6184 5160
rect 6236 5148 6242 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6236 5120 6837 5148
rect 6236 5108 6242 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 7576 5148 7604 5324
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 8478 5312 8484 5364
rect 8536 5352 8542 5364
rect 9214 5352 9220 5364
rect 8536 5324 9220 5352
rect 8536 5312 8542 5324
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 10134 5352 10140 5364
rect 9646 5324 10140 5352
rect 9646 5284 9674 5324
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10870 5312 10876 5364
rect 10928 5352 10934 5364
rect 10928 5324 15332 5352
rect 10928 5312 10934 5324
rect 10226 5284 10232 5296
rect 8128 5256 9674 5284
rect 10187 5256 10232 5284
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 7745 5219 7803 5225
rect 7745 5216 7757 5219
rect 7708 5188 7757 5216
rect 7708 5176 7714 5188
rect 7745 5185 7757 5188
rect 7791 5216 7803 5219
rect 8018 5216 8024 5228
rect 7791 5188 8024 5216
rect 7791 5185 7803 5188
rect 7745 5179 7803 5185
rect 8018 5176 8024 5188
rect 8076 5176 8082 5228
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 7576 5120 7941 5148
rect 6825 5111 6883 5117
rect 7929 5117 7941 5120
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 3881 5083 3939 5089
rect 3881 5080 3893 5083
rect 1228 5052 3893 5080
rect 3881 5049 3893 5052
rect 3927 5049 3939 5083
rect 3881 5043 3939 5049
rect 4893 5083 4951 5089
rect 4893 5049 4905 5083
rect 4939 5080 4951 5083
rect 4939 5052 7972 5080
rect 4939 5049 4951 5052
rect 4893 5043 4951 5049
rect 198 4972 204 5024
rect 256 5012 262 5024
rect 1489 5015 1547 5021
rect 1489 5012 1501 5015
rect 256 4984 1501 5012
rect 256 4972 262 4984
rect 1489 4981 1501 4984
rect 1535 4981 1547 5015
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 1489 4975 1547 4981
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 5350 4972 5356 5024
rect 5408 5012 5414 5024
rect 5537 5015 5595 5021
rect 5537 5012 5549 5015
rect 5408 4984 5549 5012
rect 5408 4972 5414 4984
rect 5537 4981 5549 4984
rect 5583 4981 5595 5015
rect 5537 4975 5595 4981
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 7101 5015 7159 5021
rect 6880 4984 6925 5012
rect 6880 4972 6886 4984
rect 7101 4981 7113 5015
rect 7147 5012 7159 5015
rect 7374 5012 7380 5024
rect 7147 4984 7380 5012
rect 7147 4981 7159 4984
rect 7101 4975 7159 4981
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 7944 5012 7972 5052
rect 8018 5040 8024 5092
rect 8076 5080 8082 5092
rect 8128 5080 8156 5256
rect 10226 5244 10232 5256
rect 10284 5244 10290 5296
rect 10594 5244 10600 5296
rect 10652 5284 10658 5296
rect 10965 5287 11023 5293
rect 10965 5284 10977 5287
rect 10652 5256 10977 5284
rect 10652 5244 10658 5256
rect 10965 5253 10977 5256
rect 11011 5284 11023 5287
rect 11330 5284 11336 5296
rect 11011 5256 11336 5284
rect 11011 5253 11023 5256
rect 10965 5247 11023 5253
rect 11330 5244 11336 5256
rect 11388 5244 11394 5296
rect 14550 5284 14556 5296
rect 12406 5256 14556 5284
rect 8849 5219 8907 5225
rect 8849 5185 8861 5219
rect 8895 5216 8907 5219
rect 9861 5219 9919 5225
rect 8895 5188 9812 5216
rect 8895 5185 8907 5188
rect 8849 5179 8907 5185
rect 8294 5108 8300 5160
rect 8352 5108 8358 5160
rect 8478 5108 8484 5160
rect 8536 5148 8542 5160
rect 8941 5151 8999 5157
rect 8941 5148 8953 5151
rect 8536 5120 8953 5148
rect 8536 5108 8542 5120
rect 8941 5117 8953 5120
rect 8987 5117 8999 5151
rect 9784 5148 9812 5188
rect 9861 5185 9873 5219
rect 9907 5216 9919 5219
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 9907 5188 9965 5216
rect 9907 5185 9919 5188
rect 9861 5179 9919 5185
rect 9953 5185 9965 5188
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 12406 5216 12434 5256
rect 14550 5244 14556 5256
rect 14608 5244 14614 5296
rect 11839 5188 12434 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 13078 5176 13084 5228
rect 13136 5216 13142 5228
rect 15304 5225 15332 5324
rect 15654 5312 15660 5364
rect 15712 5352 15718 5364
rect 15841 5355 15899 5361
rect 15841 5352 15853 5355
rect 15712 5324 15853 5352
rect 15712 5312 15718 5324
rect 15841 5321 15853 5324
rect 15887 5352 15899 5355
rect 16114 5352 16120 5364
rect 15887 5324 16120 5352
rect 15887 5321 15899 5324
rect 15841 5315 15899 5321
rect 16114 5312 16120 5324
rect 16172 5312 16178 5364
rect 42797 5355 42855 5361
rect 42797 5321 42809 5355
rect 42843 5352 42855 5355
rect 44634 5352 44640 5364
rect 42843 5324 44640 5352
rect 42843 5321 42855 5324
rect 42797 5315 42855 5321
rect 44634 5312 44640 5324
rect 44692 5312 44698 5364
rect 42610 5244 42616 5296
rect 42668 5284 42674 5296
rect 44082 5284 44088 5296
rect 42668 5256 44088 5284
rect 42668 5244 42674 5256
rect 44082 5244 44088 5256
rect 44140 5244 44146 5296
rect 44174 5244 44180 5296
rect 44232 5284 44238 5296
rect 44545 5287 44603 5293
rect 44545 5284 44557 5287
rect 44232 5256 44557 5284
rect 44232 5244 44238 5256
rect 44545 5253 44557 5256
rect 44591 5253 44603 5287
rect 44545 5247 44603 5253
rect 15289 5219 15347 5225
rect 13136 5188 13181 5216
rect 13136 5176 13142 5188
rect 15289 5185 15301 5219
rect 15335 5216 15347 5219
rect 25222 5216 25228 5228
rect 15335 5188 25228 5216
rect 15335 5185 15347 5188
rect 15289 5179 15347 5185
rect 25222 5176 25228 5188
rect 25280 5176 25286 5228
rect 43254 5216 43260 5228
rect 43215 5188 43260 5216
rect 43254 5176 43260 5188
rect 43312 5176 43318 5228
rect 43901 5219 43959 5225
rect 43901 5185 43913 5219
rect 43947 5216 43959 5219
rect 44450 5216 44456 5228
rect 43947 5188 44456 5216
rect 43947 5185 43959 5188
rect 43901 5179 43959 5185
rect 10594 5148 10600 5160
rect 9784 5120 10600 5148
rect 8941 5111 8999 5117
rect 10594 5108 10600 5120
rect 10652 5108 10658 5160
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 21358 5148 21364 5160
rect 11112 5120 21364 5148
rect 11112 5108 11118 5120
rect 21358 5108 21364 5120
rect 21416 5108 21422 5160
rect 41877 5151 41935 5157
rect 41877 5117 41889 5151
rect 41923 5148 41935 5151
rect 43916 5148 43944 5179
rect 44450 5176 44456 5188
rect 44508 5176 44514 5228
rect 45189 5219 45247 5225
rect 45189 5185 45201 5219
rect 45235 5185 45247 5219
rect 45189 5179 45247 5185
rect 45557 5219 45615 5225
rect 45557 5185 45569 5219
rect 45603 5216 45615 5219
rect 47118 5216 47124 5228
rect 45603 5188 47124 5216
rect 45603 5185 45615 5188
rect 45557 5179 45615 5185
rect 45094 5148 45100 5160
rect 41923 5120 43944 5148
rect 45055 5120 45100 5148
rect 41923 5117 41935 5120
rect 41877 5111 41935 5117
rect 45094 5108 45100 5120
rect 45152 5108 45158 5160
rect 8076 5052 8156 5080
rect 8312 5080 8340 5108
rect 9217 5083 9275 5089
rect 8312 5052 9168 5080
rect 8076 5040 8082 5052
rect 8294 5012 8300 5024
rect 7944 4984 8300 5012
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 8478 4972 8484 5024
rect 8536 5012 8542 5024
rect 8849 5015 8907 5021
rect 8849 5012 8861 5015
rect 8536 4984 8861 5012
rect 8536 4972 8542 4984
rect 8849 4981 8861 4984
rect 8895 5012 8907 5015
rect 8938 5012 8944 5024
rect 8895 4984 8944 5012
rect 8895 4981 8907 4984
rect 8849 4975 8907 4981
rect 8938 4972 8944 4984
rect 8996 4972 9002 5024
rect 9140 5012 9168 5052
rect 9217 5049 9229 5083
rect 9263 5080 9275 5083
rect 9861 5083 9919 5089
rect 9861 5080 9873 5083
rect 9263 5052 9873 5080
rect 9263 5049 9275 5052
rect 9217 5043 9275 5049
rect 9861 5049 9873 5052
rect 9907 5049 9919 5083
rect 9861 5043 9919 5049
rect 10502 5040 10508 5092
rect 10560 5080 10566 5092
rect 11609 5083 11667 5089
rect 11609 5080 11621 5083
rect 10560 5052 11621 5080
rect 10560 5040 10566 5052
rect 11609 5049 11621 5052
rect 11655 5049 11667 5083
rect 14645 5083 14703 5089
rect 14645 5080 14657 5083
rect 11609 5043 11667 5049
rect 11716 5052 14657 5080
rect 9490 5012 9496 5024
rect 9140 4984 9496 5012
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 11330 4972 11336 5024
rect 11388 5012 11394 5024
rect 11716 5012 11744 5052
rect 14645 5049 14657 5052
rect 14691 5049 14703 5083
rect 14645 5043 14703 5049
rect 43441 5083 43499 5089
rect 43441 5049 43453 5083
rect 43487 5080 43499 5083
rect 45204 5080 45232 5179
rect 47118 5176 47124 5188
rect 47176 5176 47182 5228
rect 45370 5108 45376 5160
rect 45428 5148 45434 5160
rect 45465 5151 45523 5157
rect 45465 5148 45477 5151
rect 45428 5120 45477 5148
rect 45428 5108 45434 5120
rect 45465 5117 45477 5120
rect 45511 5148 45523 5151
rect 45830 5148 45836 5160
rect 45511 5120 45836 5148
rect 45511 5117 45523 5120
rect 45465 5111 45523 5117
rect 45830 5108 45836 5120
rect 45888 5108 45894 5160
rect 43487 5052 45232 5080
rect 43487 5049 43499 5052
rect 43441 5043 43499 5049
rect 11388 4984 11744 5012
rect 11388 4972 11394 4984
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 11940 4984 12265 5012
rect 11940 4972 11946 4984
rect 12253 4981 12265 4984
rect 12299 4981 12311 5015
rect 12253 4975 12311 4981
rect 12342 4972 12348 5024
rect 12400 5012 12406 5024
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 12400 4984 12909 5012
rect 12400 4972 12406 4984
rect 12897 4981 12909 4984
rect 12943 4981 12955 5015
rect 12897 4975 12955 4981
rect 13170 4972 13176 5024
rect 13228 5012 13234 5024
rect 13541 5015 13599 5021
rect 13541 5012 13553 5015
rect 13228 4984 13553 5012
rect 13228 4972 13234 4984
rect 13541 4981 13553 4984
rect 13587 4981 13599 5015
rect 14090 5012 14096 5024
rect 14051 4984 14096 5012
rect 13541 4975 13599 4981
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 29086 5012 29092 5024
rect 29047 4984 29092 5012
rect 29086 4972 29092 4984
rect 29144 4972 29150 5024
rect 30006 5012 30012 5024
rect 29967 4984 30012 5012
rect 30006 4972 30012 4984
rect 30064 4972 30070 5024
rect 41322 5012 41328 5024
rect 41283 4984 41328 5012
rect 41322 4972 41328 4984
rect 41380 4972 41386 5024
rect 44085 5015 44143 5021
rect 44085 4981 44097 5015
rect 44131 5012 44143 5015
rect 45646 5012 45652 5024
rect 44131 4984 45652 5012
rect 44131 4981 44143 4984
rect 44085 4975 44143 4981
rect 45646 4972 45652 4984
rect 45704 4972 45710 5024
rect 46201 5015 46259 5021
rect 46201 4981 46213 5015
rect 46247 5012 46259 5015
rect 46290 5012 46296 5024
rect 46247 4984 46296 5012
rect 46247 4981 46259 4984
rect 46201 4975 46259 4981
rect 46290 4972 46296 4984
rect 46348 4972 46354 5024
rect 46658 4972 46664 5024
rect 46716 5012 46722 5024
rect 46845 5015 46903 5021
rect 46845 5012 46857 5015
rect 46716 4984 46857 5012
rect 46716 4972 46722 4984
rect 46845 4981 46857 4984
rect 46891 4981 46903 5015
rect 46845 4975 46903 4981
rect 47026 4972 47032 5024
rect 47084 5012 47090 5024
rect 47581 5015 47639 5021
rect 47581 5012 47593 5015
rect 47084 4984 47593 5012
rect 47084 4972 47090 4984
rect 47581 4981 47593 4984
rect 47627 4981 47639 5015
rect 47581 4975 47639 4981
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 2314 4808 2320 4820
rect 1627 4780 2320 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 2314 4768 2320 4780
rect 2372 4768 2378 4820
rect 2590 4768 2596 4820
rect 2648 4808 2654 4820
rect 2866 4808 2872 4820
rect 2648 4780 2872 4808
rect 2648 4768 2654 4780
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 8478 4808 8484 4820
rect 4080 4780 8484 4808
rect 658 4700 664 4752
rect 716 4740 722 4752
rect 2409 4743 2467 4749
rect 2409 4740 2421 4743
rect 716 4712 2421 4740
rect 716 4700 722 4712
rect 2409 4709 2421 4712
rect 2455 4709 2467 4743
rect 2409 4703 2467 4709
rect 4080 4684 4108 4780
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 8938 4808 8944 4820
rect 8588 4780 8708 4808
rect 8899 4780 8944 4808
rect 8588 4752 8616 4780
rect 8202 4740 8208 4752
rect 6564 4712 8208 4740
rect 753 4675 811 4681
rect 753 4641 765 4675
rect 799 4672 811 4675
rect 799 4644 1900 4672
rect 799 4641 811 4644
rect 753 4635 811 4641
rect 1026 4564 1032 4616
rect 1084 4604 1090 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 1084 4576 1409 4604
rect 1084 4564 1090 4576
rect 1397 4573 1409 4576
rect 1443 4604 1455 4607
rect 1762 4604 1768 4616
rect 1443 4576 1768 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 1762 4564 1768 4576
rect 1820 4564 1826 4616
rect 1872 4468 1900 4644
rect 4062 4632 4068 4684
rect 4120 4632 4126 4684
rect 6564 4681 6592 4712
rect 8202 4700 8208 4712
rect 8260 4700 8266 4752
rect 8570 4700 8576 4752
rect 8628 4700 8634 4752
rect 8680 4740 8708 4780
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9030 4768 9036 4820
rect 9088 4808 9094 4820
rect 9401 4811 9459 4817
rect 9088 4780 9352 4808
rect 9088 4768 9094 4780
rect 8846 4740 8852 4752
rect 8680 4712 8852 4740
rect 8846 4700 8852 4712
rect 8904 4740 8910 4752
rect 8904 4712 9168 4740
rect 8904 4700 8910 4712
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4641 6607 4675
rect 8018 4672 8024 4684
rect 6549 4635 6607 4641
rect 6840 4644 8024 4672
rect 4338 4564 4344 4616
rect 4396 4604 4402 4616
rect 5169 4607 5227 4613
rect 5169 4604 5181 4607
rect 4396 4576 5181 4604
rect 4396 4564 4402 4576
rect 5169 4573 5181 4576
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 5810 4564 5816 4616
rect 5868 4604 5874 4616
rect 6086 4604 6092 4616
rect 5868 4576 6092 4604
rect 5868 4564 5874 4576
rect 6086 4564 6092 4576
rect 6144 4604 6150 4616
rect 6273 4607 6331 4613
rect 6273 4604 6285 4607
rect 6144 4576 6285 4604
rect 6144 4564 6150 4576
rect 6273 4573 6285 4576
rect 6319 4573 6331 4607
rect 6273 4567 6331 4573
rect 2038 4496 2044 4548
rect 2096 4536 2102 4548
rect 2685 4539 2743 4545
rect 2685 4536 2697 4539
rect 2096 4508 2697 4536
rect 2096 4496 2102 4508
rect 2685 4505 2697 4508
rect 2731 4536 2743 4539
rect 3234 4536 3240 4548
rect 2731 4508 3240 4536
rect 2731 4505 2743 4508
rect 2685 4499 2743 4505
rect 3234 4496 3240 4508
rect 3292 4496 3298 4548
rect 4249 4539 4307 4545
rect 4249 4505 4261 4539
rect 4295 4536 4307 4539
rect 4430 4536 4436 4548
rect 4295 4508 4436 4536
rect 4295 4505 4307 4508
rect 4249 4499 4307 4505
rect 4430 4496 4436 4508
rect 4488 4496 4494 4548
rect 5537 4539 5595 4545
rect 5537 4505 5549 4539
rect 5583 4536 5595 4539
rect 6840 4536 6868 4644
rect 8018 4632 8024 4644
rect 8076 4632 8082 4684
rect 8294 4632 8300 4684
rect 8352 4672 8358 4684
rect 9140 4681 9168 4712
rect 9214 4700 9220 4752
rect 9272 4700 9278 4752
rect 9125 4675 9183 4681
rect 8352 4644 8432 4672
rect 8352 4632 8358 4644
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 6972 4576 7205 4604
rect 6972 4564 6978 4576
rect 7193 4573 7205 4576
rect 7239 4604 7251 4607
rect 7834 4604 7840 4616
rect 7239 4576 7840 4604
rect 7239 4573 7251 4576
rect 7193 4567 7251 4573
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 8404 4613 8432 4644
rect 9125 4641 9137 4675
rect 9171 4641 9183 4675
rect 9125 4635 9183 4641
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 8846 4564 8852 4616
rect 8904 4604 8910 4616
rect 9232 4613 9260 4700
rect 9324 4672 9352 4780
rect 9401 4777 9413 4811
rect 9447 4808 9459 4811
rect 9674 4808 9680 4820
rect 9447 4780 9680 4808
rect 9447 4777 9459 4780
rect 9401 4771 9459 4777
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 17126 4808 17132 4820
rect 9784 4780 17132 4808
rect 9490 4700 9496 4752
rect 9548 4740 9554 4752
rect 9784 4740 9812 4780
rect 17126 4768 17132 4780
rect 17184 4768 17190 4820
rect 43349 4811 43407 4817
rect 43349 4777 43361 4811
rect 43395 4808 43407 4811
rect 46382 4808 46388 4820
rect 43395 4780 46388 4808
rect 43395 4777 43407 4780
rect 43349 4771 43407 4777
rect 46382 4768 46388 4780
rect 46440 4768 46446 4820
rect 11422 4740 11428 4752
rect 9548 4712 9812 4740
rect 9968 4712 11428 4740
rect 9548 4700 9554 4712
rect 9324 4644 9674 4672
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8904 4576 8953 4604
rect 8904 4564 8910 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4573 9275 4607
rect 9646 4604 9674 4644
rect 9766 4604 9772 4616
rect 9646 4576 9772 4604
rect 9217 4567 9275 4573
rect 9766 4564 9772 4576
rect 9824 4604 9830 4616
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 9824 4576 9873 4604
rect 9824 4564 9830 4576
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 5583 4508 6868 4536
rect 7469 4539 7527 4545
rect 5583 4505 5595 4508
rect 5537 4499 5595 4505
rect 7469 4505 7481 4539
rect 7515 4536 7527 4539
rect 9968 4536 9996 4712
rect 11422 4700 11428 4712
rect 11480 4700 11486 4752
rect 11606 4700 11612 4752
rect 11664 4740 11670 4752
rect 13081 4743 13139 4749
rect 13081 4740 13093 4743
rect 11664 4712 13093 4740
rect 11664 4700 11670 4712
rect 13081 4709 13093 4712
rect 13127 4709 13139 4743
rect 13081 4703 13139 4709
rect 14366 4700 14372 4752
rect 14424 4740 14430 4752
rect 43901 4743 43959 4749
rect 43901 4740 43913 4743
rect 14424 4712 43913 4740
rect 14424 4700 14430 4712
rect 43901 4709 43913 4712
rect 43947 4709 43959 4743
rect 45370 4740 45376 4752
rect 43901 4703 43959 4709
rect 44095 4712 45376 4740
rect 11054 4672 11060 4684
rect 11015 4644 11060 4672
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 11238 4632 11244 4684
rect 11296 4672 11302 4684
rect 11790 4672 11796 4684
rect 11296 4644 11796 4672
rect 11296 4632 11302 4644
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 12802 4672 12808 4684
rect 11992 4644 12808 4672
rect 10778 4604 10784 4616
rect 10739 4576 10784 4604
rect 10778 4564 10784 4576
rect 10836 4604 10842 4616
rect 11992 4613 12020 4644
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 16942 4672 16948 4684
rect 16903 4644 16948 4672
rect 16942 4632 16948 4644
rect 17000 4632 17006 4684
rect 11977 4607 12035 4613
rect 10836 4576 11284 4604
rect 10836 4564 10842 4576
rect 7515 4508 9996 4536
rect 10137 4539 10195 4545
rect 7515 4505 7527 4508
rect 7469 4499 7527 4505
rect 10137 4505 10149 4539
rect 10183 4536 10195 4539
rect 10962 4536 10968 4548
rect 10183 4508 10968 4536
rect 10183 4505 10195 4508
rect 10137 4499 10195 4505
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 11256 4536 11284 4576
rect 11977 4573 11989 4607
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12492 4576 12537 4604
rect 12492 4564 12498 4576
rect 13814 4564 13820 4616
rect 13872 4604 13878 4616
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13872 4576 14105 4604
rect 13872 4564 13878 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 15194 4564 15200 4616
rect 15252 4604 15258 4616
rect 15657 4607 15715 4613
rect 15657 4604 15669 4607
rect 15252 4576 15669 4604
rect 15252 4564 15258 4576
rect 15657 4573 15669 4576
rect 15703 4573 15715 4607
rect 15657 4567 15715 4573
rect 28997 4607 29055 4613
rect 28997 4573 29009 4607
rect 29043 4604 29055 4607
rect 29086 4604 29092 4616
rect 29043 4576 29092 4604
rect 29043 4573 29055 4576
rect 28997 4567 29055 4573
rect 29086 4564 29092 4576
rect 29144 4604 29150 4616
rect 29914 4604 29920 4616
rect 29144 4576 29920 4604
rect 29144 4564 29150 4576
rect 29914 4564 29920 4576
rect 29972 4564 29978 4616
rect 30006 4564 30012 4616
rect 30064 4604 30070 4616
rect 30101 4607 30159 4613
rect 30101 4604 30113 4607
rect 30064 4576 30113 4604
rect 30064 4564 30070 4576
rect 30101 4573 30113 4576
rect 30147 4573 30159 4607
rect 37918 4604 37924 4616
rect 30101 4567 30159 4573
rect 35866 4576 37924 4604
rect 13630 4536 13636 4548
rect 11256 4508 13636 4536
rect 13630 4496 13636 4508
rect 13688 4496 13694 4548
rect 35866 4536 35894 4576
rect 37918 4564 37924 4576
rect 37976 4564 37982 4616
rect 42058 4564 42064 4616
rect 42116 4604 42122 4616
rect 42518 4604 42524 4616
rect 42116 4576 42524 4604
rect 42116 4564 42122 4576
rect 42518 4564 42524 4576
rect 42576 4564 42582 4616
rect 44095 4613 44123 4712
rect 45370 4700 45376 4712
rect 45428 4700 45434 4752
rect 45738 4700 45744 4752
rect 45796 4740 45802 4752
rect 45796 4712 47624 4740
rect 45796 4700 45802 4712
rect 45094 4672 45100 4684
rect 44468 4644 45100 4672
rect 44468 4613 44496 4644
rect 45094 4632 45100 4644
rect 45152 4672 45158 4684
rect 45465 4675 45523 4681
rect 45465 4672 45477 4675
rect 45152 4644 45477 4672
rect 45152 4632 45158 4644
rect 45465 4641 45477 4644
rect 45511 4641 45523 4675
rect 45465 4635 45523 4641
rect 45830 4632 45836 4684
rect 45888 4672 45894 4684
rect 45925 4675 45983 4681
rect 45925 4672 45937 4675
rect 45888 4644 45937 4672
rect 45888 4632 45894 4644
rect 45925 4641 45937 4644
rect 45971 4641 45983 4675
rect 47394 4672 47400 4684
rect 47355 4644 47400 4672
rect 45925 4635 45983 4641
rect 47394 4632 47400 4644
rect 47452 4632 47458 4684
rect 44080 4607 44138 4613
rect 44080 4573 44092 4607
rect 44126 4573 44138 4607
rect 44080 4567 44138 4573
rect 44453 4607 44511 4613
rect 44453 4573 44465 4607
rect 44499 4573 44511 4607
rect 45002 4604 45008 4616
rect 44963 4576 45008 4604
rect 44453 4567 44511 4573
rect 45002 4564 45008 4576
rect 45060 4564 45066 4616
rect 45646 4604 45652 4616
rect 45607 4576 45652 4604
rect 45646 4564 45652 4576
rect 45704 4564 45710 4616
rect 46017 4607 46075 4613
rect 46017 4573 46029 4607
rect 46063 4604 46075 4607
rect 46566 4604 46572 4616
rect 46063 4576 46572 4604
rect 46063 4573 46075 4576
rect 46017 4567 46075 4573
rect 19306 4508 35894 4536
rect 41969 4539 42027 4545
rect 4341 4471 4399 4477
rect 4341 4468 4353 4471
rect 1872 4440 4353 4468
rect 4341 4437 4353 4440
rect 4387 4437 4399 4471
rect 4341 4431 4399 4437
rect 7834 4428 7840 4480
rect 7892 4468 7898 4480
rect 8205 4471 8263 4477
rect 8205 4468 8217 4471
rect 7892 4440 8217 4468
rect 7892 4428 7898 4440
rect 8205 4437 8217 4440
rect 8251 4437 8263 4471
rect 8205 4431 8263 4437
rect 9030 4428 9036 4480
rect 9088 4468 9094 4480
rect 9582 4468 9588 4480
rect 9088 4440 9588 4468
rect 9088 4428 9094 4440
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 10594 4468 10600 4480
rect 9732 4440 10600 4468
rect 9732 4428 9738 4440
rect 10594 4428 10600 4440
rect 10652 4428 10658 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11793 4471 11851 4477
rect 11793 4468 11805 4471
rect 11112 4440 11805 4468
rect 11112 4428 11118 4440
rect 11793 4437 11805 4440
rect 11839 4437 11851 4471
rect 11793 4431 11851 4437
rect 12158 4428 12164 4480
rect 12216 4468 12222 4480
rect 14737 4471 14795 4477
rect 14737 4468 14749 4471
rect 12216 4440 14749 4468
rect 12216 4428 12222 4440
rect 14737 4437 14749 4440
rect 14783 4437 14795 4471
rect 16298 4468 16304 4480
rect 16259 4440 16304 4468
rect 14737 4431 14795 4437
rect 16298 4428 16304 4440
rect 16356 4468 16362 4480
rect 19306 4468 19334 4508
rect 41969 4505 41981 4539
rect 42015 4536 42027 4539
rect 44174 4536 44180 4548
rect 42015 4508 44180 4536
rect 42015 4505 42027 4508
rect 41969 4499 42027 4505
rect 44174 4496 44180 4508
rect 44232 4496 44238 4548
rect 44269 4539 44327 4545
rect 44269 4505 44281 4539
rect 44315 4505 44327 4539
rect 44269 4499 44327 4505
rect 28810 4468 28816 4480
rect 16356 4440 19334 4468
rect 28771 4440 28816 4468
rect 16356 4428 16362 4440
rect 28810 4428 28816 4440
rect 28868 4428 28874 4480
rect 29454 4428 29460 4480
rect 29512 4468 29518 4480
rect 29549 4471 29607 4477
rect 29549 4468 29561 4471
rect 29512 4440 29561 4468
rect 29512 4428 29518 4440
rect 29549 4437 29561 4440
rect 29595 4437 29607 4471
rect 29549 4431 29607 4437
rect 30285 4471 30343 4477
rect 30285 4437 30297 4471
rect 30331 4468 30343 4471
rect 30558 4468 30564 4480
rect 30331 4440 30564 4468
rect 30331 4437 30343 4440
rect 30285 4431 30343 4437
rect 30558 4428 30564 4440
rect 30616 4428 30622 4480
rect 30742 4468 30748 4480
rect 30703 4440 30748 4468
rect 30742 4428 30748 4440
rect 30800 4428 30806 4480
rect 31386 4468 31392 4480
rect 31347 4440 31392 4468
rect 31386 4428 31392 4440
rect 31444 4428 31450 4480
rect 40402 4468 40408 4480
rect 40363 4440 40408 4468
rect 40402 4428 40408 4440
rect 40460 4428 40466 4480
rect 40862 4468 40868 4480
rect 40823 4440 40868 4468
rect 40862 4428 40868 4440
rect 40920 4428 40926 4480
rect 41506 4468 41512 4480
rect 41467 4440 41512 4468
rect 41506 4428 41512 4440
rect 41564 4428 41570 4480
rect 42705 4471 42763 4477
rect 42705 4437 42717 4471
rect 42751 4468 42763 4471
rect 44284 4468 44312 4499
rect 44634 4496 44640 4548
rect 44692 4536 44698 4548
rect 46032 4536 46060 4567
rect 46566 4564 46572 4576
rect 46624 4564 46630 4616
rect 47596 4613 47624 4712
rect 47581 4607 47639 4613
rect 47581 4573 47593 4607
rect 47627 4573 47639 4607
rect 47581 4567 47639 4573
rect 47762 4564 47768 4616
rect 47820 4604 47826 4616
rect 47949 4607 48007 4613
rect 47949 4604 47961 4607
rect 47820 4576 47961 4604
rect 47820 4564 47826 4576
rect 47949 4573 47961 4576
rect 47995 4573 48007 4607
rect 47949 4567 48007 4573
rect 48038 4564 48044 4616
rect 48096 4604 48102 4616
rect 48096 4576 48141 4604
rect 48096 4564 48102 4576
rect 46934 4536 46940 4548
rect 44692 4508 46060 4536
rect 46895 4508 46940 4536
rect 44692 4496 44698 4508
rect 46934 4496 46940 4508
rect 46992 4496 46998 4548
rect 42751 4440 44312 4468
rect 42751 4437 42763 4440
rect 42705 4431 42763 4437
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 1854 4224 1860 4276
rect 1912 4264 1918 4276
rect 1912 4236 3004 4264
rect 1912 4224 1918 4236
rect 1946 4196 1952 4208
rect 1907 4168 1952 4196
rect 1946 4156 1952 4168
rect 2004 4156 2010 4208
rect 750 4088 756 4140
rect 808 4128 814 4140
rect 1486 4128 1492 4140
rect 808 4100 1492 4128
rect 808 4088 814 4100
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 2314 4128 2320 4140
rect 2275 4100 2320 4128
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4126 2835 4131
rect 2976 4128 3004 4236
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3108 4236 3740 4264
rect 3108 4224 3114 4236
rect 3712 4208 3740 4236
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 5629 4267 5687 4273
rect 5629 4264 5641 4267
rect 4488 4236 5641 4264
rect 4488 4224 4494 4236
rect 5629 4233 5641 4236
rect 5675 4233 5687 4267
rect 5629 4227 5687 4233
rect 5902 4224 5908 4276
rect 5960 4264 5966 4276
rect 5960 4236 6868 4264
rect 5960 4224 5966 4236
rect 3694 4156 3700 4208
rect 3752 4156 3758 4208
rect 4338 4196 4344 4208
rect 3988 4168 4344 4196
rect 2884 4126 3004 4128
rect 2823 4100 3004 4126
rect 3053 4131 3111 4137
rect 2823 4098 2912 4100
rect 2823 4097 2835 4098
rect 2777 4091 2835 4097
rect 3053 4097 3065 4131
rect 3099 4128 3111 4131
rect 3234 4128 3240 4140
rect 3099 4100 3240 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3789 4131 3847 4137
rect 3789 4097 3801 4131
rect 3835 4128 3847 4131
rect 3988 4128 4016 4168
rect 4338 4156 4344 4168
rect 4396 4156 4402 4208
rect 6546 4156 6552 4208
rect 6604 4156 6610 4208
rect 6840 4205 6868 4236
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 8573 4267 8631 4273
rect 8573 4264 8585 4267
rect 8536 4236 8585 4264
rect 8536 4224 8542 4236
rect 8573 4233 8585 4236
rect 8619 4233 8631 4267
rect 8573 4227 8631 4233
rect 8846 4224 8852 4276
rect 8904 4224 8910 4276
rect 9582 4224 9588 4276
rect 9640 4264 9646 4276
rect 9766 4264 9772 4276
rect 9640 4236 9772 4264
rect 9640 4224 9646 4236
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 10336 4236 10548 4264
rect 6825 4199 6883 4205
rect 6825 4165 6837 4199
rect 6871 4165 6883 4199
rect 7006 4196 7012 4208
rect 6825 4159 6883 4165
rect 6932 4168 7012 4196
rect 3835 4100 4016 4128
rect 3835 4097 3847 4100
rect 3789 4091 3847 4097
rect 4062 4088 4068 4140
rect 4120 4088 4126 4140
rect 4522 4137 4528 4140
rect 4516 4128 4528 4137
rect 4483 4100 4528 4128
rect 4516 4091 4528 4100
rect 4522 4088 4528 4091
rect 4580 4088 4586 4140
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 6564 4128 6592 4156
rect 5960 4100 6592 4128
rect 5960 4088 5966 4100
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4060 2927 4063
rect 4080 4060 4108 4088
rect 2915 4032 3004 4060
rect 2915 4029 2927 4032
rect 2869 4023 2927 4029
rect 2976 4004 3004 4032
rect 3068 4032 4108 4060
rect 4249 4063 4307 4069
rect 937 3995 995 4001
rect 937 3961 949 3995
rect 983 3992 995 3995
rect 1486 3992 1492 4004
rect 983 3964 1492 3992
rect 983 3961 995 3964
rect 937 3955 995 3961
rect 1486 3952 1492 3964
rect 1544 3952 1550 4004
rect 2958 3952 2964 4004
rect 3016 3952 3022 4004
rect 1118 3884 1124 3936
rect 1176 3924 1182 3936
rect 2777 3927 2835 3933
rect 2777 3924 2789 3927
rect 1176 3896 2789 3924
rect 1176 3884 1182 3896
rect 2777 3893 2789 3896
rect 2823 3924 2835 3927
rect 3068 3924 3096 4032
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 3234 3924 3240 3936
rect 2823 3896 3096 3924
rect 3195 3896 3240 3924
rect 2823 3893 2835 3896
rect 2777 3887 2835 3893
rect 3234 3884 3240 3896
rect 3292 3884 3298 3936
rect 4264 3924 4292 4023
rect 6546 4020 6552 4072
rect 6604 4060 6610 4072
rect 6932 4060 6960 4168
rect 7006 4156 7012 4168
rect 7064 4156 7070 4208
rect 8864 4196 8892 4224
rect 7116 4168 8892 4196
rect 7116 4128 7144 4168
rect 6604 4032 6960 4060
rect 7024 4100 7144 4128
rect 6604 4020 6610 4032
rect 7024 3924 7052 4100
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 8205 4131 8263 4137
rect 8205 4128 8217 4131
rect 8168 4100 8217 4128
rect 8168 4088 8174 4100
rect 8205 4097 8217 4100
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 8220 3992 8248 4091
rect 8478 4088 8484 4140
rect 8536 4128 8542 4140
rect 8757 4131 8815 4137
rect 8757 4128 8769 4131
rect 8536 4100 8769 4128
rect 8536 4088 8542 4100
rect 8757 4097 8769 4100
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4128 9275 4131
rect 9398 4128 9404 4140
rect 9263 4100 9404 4128
rect 9263 4097 9275 4100
rect 9217 4091 9275 4097
rect 8297 4063 8355 4069
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 8386 4060 8392 4072
rect 8343 4032 8392 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8772 4060 8800 4091
rect 9398 4088 9404 4100
rect 9456 4088 9462 4140
rect 9493 4131 9551 4137
rect 9493 4097 9505 4131
rect 9539 4097 9551 4131
rect 9493 4091 9551 4097
rect 9508 4060 9536 4091
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 10336 4128 10364 4236
rect 10520 4196 10548 4236
rect 10594 4224 10600 4276
rect 10652 4264 10658 4276
rect 13078 4264 13084 4276
rect 10652 4236 13084 4264
rect 10652 4224 10658 4236
rect 13078 4224 13084 4236
rect 13136 4224 13142 4276
rect 41506 4224 41512 4276
rect 41564 4264 41570 4276
rect 47762 4264 47768 4276
rect 41564 4236 47768 4264
rect 41564 4224 41570 4236
rect 47762 4224 47768 4236
rect 47820 4224 47826 4276
rect 10686 4196 10692 4208
rect 10520 4168 10692 4196
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 13998 4196 14004 4208
rect 13188 4168 14004 4196
rect 10413 4131 10471 4137
rect 10413 4128 10425 4131
rect 9640 4100 9996 4128
rect 10336 4100 10425 4128
rect 9640 4088 9646 4100
rect 9968 4072 9996 4100
rect 10413 4097 10425 4100
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 13188 4128 13216 4168
rect 13998 4156 14004 4168
rect 14056 4156 14062 4208
rect 41322 4196 41328 4208
rect 30668 4168 31524 4196
rect 12575 4100 13216 4128
rect 13265 4131 13323 4137
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 16942 4128 16948 4140
rect 13311 4100 16948 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 8772 4032 9536 4060
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 9732 4032 9777 4060
rect 9732 4020 9738 4032
rect 9950 4020 9956 4072
rect 10008 4020 10014 4072
rect 10686 4060 10692 4072
rect 10647 4032 10692 4060
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 11808 4060 11836 4091
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4128 20131 4131
rect 20162 4128 20168 4140
rect 20119 4100 20168 4128
rect 20119 4097 20131 4100
rect 20073 4091 20131 4097
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 20346 4088 20352 4140
rect 20404 4128 20410 4140
rect 30668 4128 30696 4168
rect 20404 4100 30696 4128
rect 20404 4088 20410 4100
rect 30742 4088 30748 4140
rect 30800 4128 30806 4140
rect 31386 4128 31392 4140
rect 30800 4100 30845 4128
rect 31347 4100 31392 4128
rect 30800 4088 30806 4100
rect 31386 4088 31392 4100
rect 31444 4088 31450 4140
rect 31496 4128 31524 4168
rect 40880 4168 41328 4196
rect 40880 4128 40908 4168
rect 41322 4156 41328 4168
rect 41380 4156 41386 4208
rect 45830 4196 45836 4208
rect 45020 4168 45836 4196
rect 31496 4100 40908 4128
rect 41233 4131 41291 4137
rect 41233 4097 41245 4131
rect 41279 4128 41291 4131
rect 41690 4128 41696 4140
rect 41279 4100 41696 4128
rect 41279 4097 41291 4100
rect 41233 4091 41291 4097
rect 41690 4088 41696 4100
rect 41748 4088 41754 4140
rect 43441 4131 43499 4137
rect 43441 4097 43453 4131
rect 43487 4128 43499 4131
rect 45020 4128 45048 4168
rect 45830 4156 45836 4168
rect 45888 4156 45894 4208
rect 45186 4128 45192 4140
rect 43487 4100 45048 4128
rect 45147 4100 45192 4128
rect 43487 4097 43499 4100
rect 43441 4091 43499 4097
rect 45186 4088 45192 4100
rect 45244 4088 45250 4140
rect 45554 4128 45560 4140
rect 45515 4100 45560 4128
rect 45554 4088 45560 4100
rect 45612 4088 45618 4140
rect 45646 4088 45652 4140
rect 45704 4128 45710 4140
rect 47857 4131 47915 4137
rect 47857 4128 47869 4131
rect 45704 4100 47869 4128
rect 45704 4088 45710 4100
rect 47857 4097 47869 4100
rect 47903 4097 47915 4131
rect 47857 4091 47915 4097
rect 48682 4088 48688 4140
rect 48740 4128 48746 4140
rect 48961 4131 49019 4137
rect 48961 4128 48973 4131
rect 48740 4100 48973 4128
rect 48740 4088 48746 4100
rect 48961 4097 48973 4100
rect 49007 4097 49019 4131
rect 48961 4091 49019 4097
rect 16298 4060 16304 4072
rect 11808 4032 16304 4060
rect 16298 4020 16304 4032
rect 16356 4020 16362 4072
rect 17034 4020 17040 4072
rect 17092 4060 17098 4072
rect 44545 4063 44603 4069
rect 44545 4060 44557 4063
rect 17092 4032 44557 4060
rect 17092 4020 17098 4032
rect 44545 4029 44557 4032
rect 44591 4029 44603 4063
rect 45094 4060 45100 4072
rect 45055 4032 45100 4060
rect 44545 4023 44603 4029
rect 45094 4020 45100 4032
rect 45152 4020 45158 4072
rect 45370 4020 45376 4072
rect 45428 4060 45434 4072
rect 45465 4063 45523 4069
rect 45465 4060 45477 4063
rect 45428 4032 45477 4060
rect 45428 4020 45434 4032
rect 45465 4029 45477 4032
rect 45511 4029 45523 4063
rect 47210 4060 47216 4072
rect 45465 4023 45523 4029
rect 45664 4032 47216 4060
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 8220 3964 9321 3992
rect 9309 3961 9321 3964
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 9398 3952 9404 4004
rect 9456 3952 9462 4004
rect 9784 3964 10640 3992
rect 4264 3896 7052 3924
rect 7101 3927 7159 3933
rect 7101 3893 7113 3927
rect 7147 3924 7159 3927
rect 7834 3924 7840 3936
rect 7147 3896 7840 3924
rect 7147 3893 7159 3896
rect 7101 3887 7159 3893
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 8386 3884 8392 3936
rect 8444 3924 8450 3936
rect 9416 3924 9444 3952
rect 8444 3896 9444 3924
rect 8444 3884 8450 3896
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 9784 3924 9812 3964
rect 9548 3896 9812 3924
rect 9548 3884 9554 3896
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 10502 3924 10508 3936
rect 10376 3896 10508 3924
rect 10376 3884 10382 3896
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 10612 3924 10640 3964
rect 10962 3952 10968 4004
rect 11020 3992 11026 4004
rect 13725 3995 13783 4001
rect 13725 3992 13737 3995
rect 11020 3964 13737 3992
rect 11020 3952 11026 3964
rect 13725 3961 13737 3964
rect 13771 3961 13783 3995
rect 13725 3955 13783 3961
rect 13832 3964 14504 3992
rect 11609 3927 11667 3933
rect 11609 3924 11621 3927
rect 10612 3896 11621 3924
rect 11609 3893 11621 3896
rect 11655 3893 11667 3927
rect 11609 3887 11667 3893
rect 11790 3884 11796 3936
rect 11848 3924 11854 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 11848 3896 12357 3924
rect 11848 3884 11854 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12345 3887 12403 3893
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 13081 3927 13139 3933
rect 13081 3924 13093 3927
rect 12768 3896 13093 3924
rect 12768 3884 12774 3896
rect 13081 3893 13093 3896
rect 13127 3893 13139 3927
rect 13081 3887 13139 3893
rect 13446 3884 13452 3936
rect 13504 3924 13510 3936
rect 13832 3924 13860 3964
rect 14366 3924 14372 3936
rect 13504 3896 13860 3924
rect 14327 3896 14372 3924
rect 13504 3884 13510 3896
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 14476 3924 14504 3964
rect 14550 3952 14556 4004
rect 14608 3992 14614 4004
rect 15657 3995 15715 4001
rect 15657 3992 15669 3995
rect 14608 3964 15669 3992
rect 14608 3952 14614 3964
rect 15657 3961 15669 3964
rect 15703 3961 15715 3995
rect 15657 3955 15715 3961
rect 17126 3952 17132 4004
rect 17184 3992 17190 4004
rect 22097 3995 22155 4001
rect 22097 3992 22109 3995
rect 17184 3964 22109 3992
rect 17184 3952 17190 3964
rect 22097 3961 22109 3964
rect 22143 3992 22155 3995
rect 22278 3992 22284 4004
rect 22143 3964 22284 3992
rect 22143 3961 22155 3964
rect 22097 3955 22155 3961
rect 22278 3952 22284 3964
rect 22336 3952 22342 4004
rect 29730 3952 29736 4004
rect 29788 3992 29794 4004
rect 30742 3992 30748 4004
rect 29788 3964 30748 3992
rect 29788 3952 29794 3964
rect 30742 3952 30748 3964
rect 30800 3952 30806 4004
rect 40129 3995 40187 4001
rect 40129 3992 40141 3995
rect 30852 3964 40141 3992
rect 15013 3927 15071 3933
rect 15013 3924 15025 3927
rect 14476 3896 15025 3924
rect 15013 3893 15025 3896
rect 15059 3893 15071 3927
rect 15013 3887 15071 3893
rect 16390 3884 16396 3936
rect 16448 3924 16454 3936
rect 16669 3927 16727 3933
rect 16669 3924 16681 3927
rect 16448 3896 16681 3924
rect 16448 3884 16454 3896
rect 16669 3893 16681 3896
rect 16715 3893 16727 3927
rect 16669 3887 16727 3893
rect 17218 3884 17224 3936
rect 17276 3924 17282 3936
rect 17313 3927 17371 3933
rect 17313 3924 17325 3927
rect 17276 3896 17325 3924
rect 17276 3884 17282 3896
rect 17313 3893 17325 3896
rect 17359 3893 17371 3927
rect 18414 3924 18420 3936
rect 18375 3896 18420 3924
rect 17313 3887 17371 3893
rect 18414 3884 18420 3896
rect 18472 3884 18478 3936
rect 27982 3924 27988 3936
rect 27943 3896 27988 3924
rect 27982 3884 27988 3896
rect 28040 3884 28046 3936
rect 28626 3924 28632 3936
rect 28587 3896 28632 3924
rect 28626 3884 28632 3896
rect 28684 3884 28690 3936
rect 28902 3884 28908 3936
rect 28960 3924 28966 3936
rect 29089 3927 29147 3933
rect 29089 3924 29101 3927
rect 28960 3896 29101 3924
rect 28960 3884 28966 3896
rect 29089 3893 29101 3896
rect 29135 3893 29147 3927
rect 30098 3924 30104 3936
rect 30059 3896 30104 3924
rect 29089 3887 29147 3893
rect 30098 3884 30104 3896
rect 30156 3884 30162 3936
rect 30190 3884 30196 3936
rect 30248 3924 30254 3936
rect 30561 3927 30619 3933
rect 30561 3924 30573 3927
rect 30248 3896 30573 3924
rect 30248 3884 30254 3896
rect 30561 3893 30573 3896
rect 30607 3893 30619 3927
rect 30561 3887 30619 3893
rect 30650 3884 30656 3936
rect 30708 3924 30714 3936
rect 30852 3924 30880 3964
rect 40129 3961 40141 3964
rect 40175 3992 40187 3995
rect 45554 3992 45560 4004
rect 40175 3964 45560 3992
rect 40175 3961 40187 3964
rect 40129 3955 40187 3961
rect 45554 3952 45560 3964
rect 45612 3952 45618 4004
rect 31202 3924 31208 3936
rect 30708 3896 30880 3924
rect 31163 3896 31208 3924
rect 30708 3884 30714 3896
rect 31202 3884 31208 3896
rect 31260 3884 31266 3936
rect 40678 3924 40684 3936
rect 40639 3896 40684 3924
rect 40678 3884 40684 3896
rect 40736 3884 40742 3936
rect 41874 3924 41880 3936
rect 41835 3896 41880 3924
rect 41874 3884 41880 3896
rect 41932 3884 41938 3936
rect 42794 3924 42800 3936
rect 42755 3896 42800 3924
rect 42794 3884 42800 3896
rect 42852 3884 42858 3936
rect 44085 3927 44143 3933
rect 44085 3893 44097 3927
rect 44131 3924 44143 3927
rect 45664 3924 45692 4032
rect 47210 4020 47216 4032
rect 47268 4020 47274 4072
rect 46014 3952 46020 4004
rect 46072 3992 46078 4004
rect 46845 3995 46903 4001
rect 46845 3992 46857 3995
rect 46072 3964 46857 3992
rect 46072 3952 46078 3964
rect 46845 3961 46857 3964
rect 46891 3961 46903 3995
rect 48130 3992 48136 4004
rect 46845 3955 46903 3961
rect 47964 3964 48136 3992
rect 44131 3896 45692 3924
rect 44131 3893 44143 3896
rect 44085 3887 44143 3893
rect 45738 3884 45744 3936
rect 45796 3924 45802 3936
rect 46201 3927 46259 3933
rect 46201 3924 46213 3927
rect 45796 3896 46213 3924
rect 45796 3884 45802 3896
rect 46201 3893 46213 3896
rect 46247 3893 46259 3927
rect 46201 3887 46259 3893
rect 46382 3884 46388 3936
rect 46440 3924 46446 3936
rect 47964 3924 47992 3964
rect 48130 3952 48136 3964
rect 48188 3952 48194 4004
rect 46440 3896 47992 3924
rect 48041 3927 48099 3933
rect 46440 3884 46446 3896
rect 48041 3893 48053 3927
rect 48087 3924 48099 3927
rect 49786 3924 49792 3936
rect 48087 3896 49792 3924
rect 48087 3893 48099 3896
rect 48041 3887 48099 3893
rect 49786 3884 49792 3896
rect 49844 3884 49850 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 842 3680 848 3732
rect 900 3720 906 3732
rect 1857 3723 1915 3729
rect 1857 3720 1869 3723
rect 900 3692 1869 3720
rect 900 3680 906 3692
rect 1857 3689 1869 3692
rect 1903 3689 1915 3723
rect 1857 3683 1915 3689
rect 3053 3723 3111 3729
rect 3053 3689 3065 3723
rect 3099 3720 3111 3723
rect 3142 3720 3148 3732
rect 3099 3692 3148 3720
rect 3099 3689 3111 3692
rect 3053 3683 3111 3689
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 3789 3723 3847 3729
rect 3789 3720 3801 3723
rect 3292 3692 3801 3720
rect 3292 3680 3298 3692
rect 3789 3689 3801 3692
rect 3835 3689 3847 3723
rect 4890 3720 4896 3732
rect 3789 3683 3847 3689
rect 4172 3692 4896 3720
rect 1946 3612 1952 3664
rect 2004 3652 2010 3664
rect 2866 3652 2872 3664
rect 2004 3624 2872 3652
rect 2004 3612 2010 3624
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 3694 3652 3700 3664
rect 3344 3624 3700 3652
rect 658 3476 664 3528
rect 716 3516 722 3528
rect 2130 3516 2136 3528
rect 716 3488 2136 3516
rect 716 3476 722 3488
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 3344 3516 3372 3624
rect 3694 3612 3700 3624
rect 3752 3612 3758 3664
rect 2240 3488 3372 3516
rect 937 3451 995 3457
rect 937 3417 949 3451
rect 983 3448 995 3451
rect 2240 3448 2268 3488
rect 983 3420 2268 3448
rect 2777 3451 2835 3457
rect 983 3417 995 3420
rect 937 3411 995 3417
rect 2777 3417 2789 3451
rect 2823 3448 2835 3451
rect 2884 3448 2912 3488
rect 3694 3476 3700 3528
rect 3752 3516 3758 3528
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 3752 3488 3985 3516
rect 3752 3476 3758 3488
rect 3973 3485 3985 3488
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4172 3516 4200 3692
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 6178 3680 6184 3732
rect 6236 3720 6242 3732
rect 6273 3723 6331 3729
rect 6273 3720 6285 3723
rect 6236 3692 6285 3720
rect 6236 3680 6242 3692
rect 6273 3689 6285 3692
rect 6319 3689 6331 3723
rect 6273 3683 6331 3689
rect 6733 3723 6791 3729
rect 6733 3689 6745 3723
rect 6779 3720 6791 3723
rect 6822 3720 6828 3732
rect 6779 3692 6828 3720
rect 6779 3689 6791 3692
rect 6733 3683 6791 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 9306 3720 9312 3732
rect 8352 3692 9312 3720
rect 8352 3680 8358 3692
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 11790 3720 11796 3732
rect 9646 3692 11796 3720
rect 4249 3655 4307 3661
rect 4249 3621 4261 3655
rect 4295 3652 4307 3655
rect 7469 3655 7527 3661
rect 7469 3652 7481 3655
rect 4295 3624 7481 3652
rect 4295 3621 4307 3624
rect 4249 3615 4307 3621
rect 7469 3621 7481 3624
rect 7515 3621 7527 3655
rect 7469 3615 7527 3621
rect 8386 3612 8392 3664
rect 8444 3652 8450 3664
rect 8754 3652 8760 3664
rect 8444 3624 8760 3652
rect 8444 3612 8450 3624
rect 8754 3612 8760 3624
rect 8812 3612 8818 3664
rect 8846 3612 8852 3664
rect 8904 3652 8910 3664
rect 9646 3652 9674 3692
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 11974 3680 11980 3732
rect 12032 3680 12038 3732
rect 12158 3680 12164 3732
rect 12216 3720 12222 3732
rect 14366 3720 14372 3732
rect 12216 3692 14372 3720
rect 12216 3680 12222 3692
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 14642 3680 14648 3732
rect 14700 3720 14706 3732
rect 40678 3720 40684 3732
rect 14700 3692 40684 3720
rect 14700 3680 14706 3692
rect 40678 3680 40684 3692
rect 40736 3680 40742 3732
rect 41877 3723 41935 3729
rect 41877 3689 41889 3723
rect 41923 3720 41935 3723
rect 44910 3720 44916 3732
rect 41923 3692 44916 3720
rect 41923 3689 41935 3692
rect 41877 3683 41935 3689
rect 44910 3680 44916 3692
rect 44968 3680 44974 3732
rect 45097 3723 45155 3729
rect 45097 3720 45109 3723
rect 45020 3692 45109 3720
rect 8904 3624 9674 3652
rect 8904 3612 8910 3624
rect 9858 3612 9864 3664
rect 9916 3652 9922 3664
rect 10410 3652 10416 3664
rect 9916 3624 10416 3652
rect 9916 3612 9922 3624
rect 10410 3612 10416 3624
rect 10468 3612 10474 3664
rect 11992 3652 12020 3680
rect 12713 3655 12771 3661
rect 12713 3652 12725 3655
rect 11992 3624 12725 3652
rect 12713 3621 12725 3624
rect 12759 3621 12771 3655
rect 12713 3615 12771 3621
rect 14826 3612 14832 3664
rect 14884 3652 14890 3664
rect 16117 3655 16175 3661
rect 16117 3652 16129 3655
rect 14884 3624 16129 3652
rect 14884 3612 14890 3624
rect 16117 3621 16129 3624
rect 16163 3621 16175 3655
rect 23750 3652 23756 3664
rect 23711 3624 23756 3652
rect 16117 3615 16175 3621
rect 23750 3612 23756 3624
rect 23808 3612 23814 3664
rect 29546 3612 29552 3664
rect 29604 3652 29610 3664
rect 30193 3655 30251 3661
rect 30193 3652 30205 3655
rect 29604 3624 30205 3652
rect 29604 3612 29610 3624
rect 30193 3621 30205 3624
rect 30239 3621 30251 3655
rect 30193 3615 30251 3621
rect 30282 3612 30288 3664
rect 30340 3652 30346 3664
rect 31386 3652 31392 3664
rect 30340 3624 31392 3652
rect 30340 3612 30346 3624
rect 31386 3612 31392 3624
rect 31444 3612 31450 3664
rect 39298 3612 39304 3664
rect 39356 3652 39362 3664
rect 45020 3652 45048 3692
rect 45097 3689 45109 3692
rect 45143 3689 45155 3723
rect 45462 3720 45468 3732
rect 45097 3683 45155 3689
rect 45388 3692 45468 3720
rect 39356 3624 45048 3652
rect 39356 3612 39362 3624
rect 6549 3587 6607 3593
rect 6549 3584 6561 3587
rect 6380 3556 6561 3584
rect 4338 3516 4344 3528
rect 4172 3488 4344 3516
rect 4065 3479 4123 3485
rect 2823 3420 2912 3448
rect 2823 3417 2835 3420
rect 2777 3411 2835 3417
rect 2958 3408 2964 3460
rect 3016 3448 3022 3460
rect 3789 3451 3847 3457
rect 3789 3448 3801 3451
rect 3016 3420 3801 3448
rect 3016 3408 3022 3420
rect 3789 3417 3801 3420
rect 3835 3417 3847 3451
rect 3789 3411 3847 3417
rect 3142 3340 3148 3392
rect 3200 3380 3206 3392
rect 4080 3380 4108 3479
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 4982 3476 4988 3528
rect 5040 3516 5046 3528
rect 5166 3516 5172 3528
rect 5040 3488 5172 3516
rect 5040 3476 5046 3488
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 4614 3408 4620 3460
rect 4672 3448 4678 3460
rect 5350 3448 5356 3460
rect 4672 3420 5356 3448
rect 4672 3408 4678 3420
rect 5350 3408 5356 3420
rect 5408 3408 5414 3460
rect 3200 3352 4108 3380
rect 3200 3340 3206 3352
rect 4522 3340 4528 3392
rect 4580 3380 4586 3392
rect 5261 3383 5319 3389
rect 5261 3380 5273 3383
rect 4580 3352 5273 3380
rect 4580 3340 4586 3352
rect 5261 3349 5273 3352
rect 5307 3349 5319 3383
rect 6380 3380 6408 3556
rect 6549 3553 6561 3556
rect 6595 3553 6607 3587
rect 6549 3547 6607 3553
rect 6638 3544 6644 3596
rect 6696 3584 6702 3596
rect 6822 3584 6828 3596
rect 6696 3556 6828 3584
rect 6696 3544 6702 3556
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 7926 3584 7932 3596
rect 7887 3556 7932 3584
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 9030 3544 9036 3596
rect 9088 3584 9094 3596
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 9088 3556 9137 3584
rect 9088 3544 9094 3556
rect 9125 3553 9137 3556
rect 9171 3553 9183 3587
rect 9950 3584 9956 3596
rect 9125 3547 9183 3553
rect 9220 3556 9956 3584
rect 6457 3519 6515 3525
rect 6457 3485 6469 3519
rect 6503 3485 6515 3519
rect 7098 3516 7104 3528
rect 6457 3479 6515 3485
rect 6656 3488 7104 3516
rect 6472 3448 6500 3479
rect 6656 3448 6684 3488
rect 7098 3476 7104 3488
rect 7156 3476 7162 3528
rect 7374 3516 7380 3528
rect 7335 3488 7380 3516
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 7653 3519 7711 3525
rect 7653 3485 7665 3519
rect 7699 3485 7711 3519
rect 7653 3479 7711 3485
rect 6472 3420 6684 3448
rect 6733 3451 6791 3457
rect 6733 3417 6745 3451
rect 6779 3448 6791 3451
rect 7466 3448 7472 3460
rect 6779 3420 7472 3448
rect 6779 3417 6791 3420
rect 6733 3411 6791 3417
rect 7466 3408 7472 3420
rect 7524 3408 7530 3460
rect 7668 3448 7696 3479
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 8938 3516 8944 3528
rect 8352 3488 8944 3516
rect 8352 3476 8358 3488
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 9220 3448 9248 3556
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 10502 3544 10508 3596
rect 10560 3544 10566 3596
rect 11422 3584 11428 3596
rect 10796 3556 11428 3584
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9824 3488 9873 3516
rect 9824 3476 9830 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 10137 3519 10195 3525
rect 10137 3485 10149 3519
rect 10183 3516 10195 3519
rect 10520 3516 10548 3544
rect 10796 3525 10824 3556
rect 11422 3544 11428 3556
rect 11480 3544 11486 3596
rect 11885 3587 11943 3593
rect 11885 3553 11897 3587
rect 11931 3553 11943 3587
rect 11885 3547 11943 3553
rect 10183 3488 10548 3516
rect 10781 3519 10839 3525
rect 10183 3485 10195 3488
rect 10137 3479 10195 3485
rect 10781 3485 10793 3519
rect 10827 3485 10839 3519
rect 10781 3479 10839 3485
rect 10796 3448 10824 3479
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11296 3488 11713 3516
rect 11296 3476 11302 3488
rect 11701 3485 11713 3488
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 11054 3448 11060 3460
rect 7668 3420 9248 3448
rect 9508 3420 10824 3448
rect 11015 3420 11060 3448
rect 9508 3392 9536 3420
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 11900 3448 11928 3547
rect 12618 3544 12624 3596
rect 12676 3584 12682 3596
rect 13357 3587 13415 3593
rect 13357 3584 13369 3587
rect 12676 3556 13369 3584
rect 12676 3544 12682 3556
rect 13357 3553 13369 3556
rect 13403 3553 13415 3587
rect 13357 3547 13415 3553
rect 14274 3544 14280 3596
rect 14332 3584 14338 3596
rect 14332 3556 14412 3584
rect 14332 3544 14338 3556
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3516 12955 3519
rect 13262 3516 13268 3528
rect 12943 3488 13268 3516
rect 12943 3485 12955 3488
rect 12897 3479 12955 3485
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 14384 3525 14412 3556
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 16761 3587 16819 3593
rect 16761 3584 16773 3587
rect 16080 3556 16773 3584
rect 16080 3544 16086 3556
rect 16761 3553 16773 3556
rect 16807 3553 16819 3587
rect 16761 3547 16819 3553
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3485 14427 3519
rect 14369 3479 14427 3485
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 14829 3519 14887 3525
rect 14829 3516 14841 3519
rect 14792 3488 14841 3516
rect 14792 3476 14798 3488
rect 14829 3485 14841 3488
rect 14875 3485 14887 3519
rect 14829 3479 14887 3485
rect 15010 3476 15016 3528
rect 15068 3516 15074 3528
rect 15473 3519 15531 3525
rect 15473 3516 15485 3519
rect 15068 3488 15485 3516
rect 15068 3476 15074 3488
rect 15473 3485 15485 3488
rect 15519 3485 15531 3519
rect 15473 3479 15531 3485
rect 16942 3476 16948 3528
rect 17000 3516 17006 3528
rect 17405 3519 17463 3525
rect 17405 3516 17417 3519
rect 17000 3488 17417 3516
rect 17000 3476 17006 3488
rect 17405 3485 17417 3488
rect 17451 3485 17463 3519
rect 17405 3479 17463 3485
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 18049 3519 18107 3525
rect 18049 3516 18061 3519
rect 17920 3488 18061 3516
rect 17920 3476 17926 3488
rect 18049 3485 18061 3488
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 19058 3476 19064 3528
rect 19116 3516 19122 3528
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 19116 3488 19257 3516
rect 19116 3476 19122 3488
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 19889 3519 19947 3525
rect 19889 3516 19901 3519
rect 19484 3488 19901 3516
rect 19484 3476 19490 3488
rect 19889 3485 19901 3488
rect 19935 3485 19947 3519
rect 20530 3516 20536 3528
rect 20491 3488 20536 3516
rect 19889 3479 19947 3485
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20806 3476 20812 3528
rect 20864 3516 20870 3528
rect 21177 3519 21235 3525
rect 21177 3516 21189 3519
rect 20864 3488 21189 3516
rect 20864 3476 20870 3488
rect 21177 3485 21189 3488
rect 21223 3485 21235 3519
rect 21177 3479 21235 3485
rect 21450 3476 21456 3528
rect 21508 3516 21514 3528
rect 21821 3519 21879 3525
rect 21821 3516 21833 3519
rect 21508 3488 21833 3516
rect 21508 3476 21514 3488
rect 21821 3485 21833 3488
rect 21867 3485 21879 3519
rect 21821 3479 21879 3485
rect 22370 3476 22376 3528
rect 22428 3516 22434 3528
rect 22465 3519 22523 3525
rect 22465 3516 22477 3519
rect 22428 3488 22477 3516
rect 22428 3476 22434 3488
rect 22465 3485 22477 3488
rect 22511 3485 22523 3519
rect 23290 3516 23296 3528
rect 23251 3488 23296 3516
rect 22465 3479 22523 3485
rect 23290 3476 23296 3488
rect 23348 3476 23354 3528
rect 24118 3476 24124 3528
rect 24176 3516 24182 3528
rect 24397 3519 24455 3525
rect 24397 3516 24409 3519
rect 24176 3488 24409 3516
rect 24176 3476 24182 3488
rect 24397 3485 24409 3488
rect 24443 3485 24455 3519
rect 25038 3516 25044 3528
rect 24999 3488 25044 3516
rect 24397 3479 24455 3485
rect 25038 3476 25044 3488
rect 25096 3476 25102 3528
rect 25958 3516 25964 3528
rect 25919 3488 25964 3516
rect 25958 3476 25964 3488
rect 26016 3476 26022 3528
rect 26234 3476 26240 3528
rect 26292 3516 26298 3528
rect 26421 3519 26479 3525
rect 26421 3516 26433 3519
rect 26292 3488 26433 3516
rect 26292 3476 26298 3488
rect 26421 3485 26433 3488
rect 26467 3485 26479 3519
rect 26421 3479 26479 3485
rect 27341 3519 27399 3525
rect 27341 3485 27353 3519
rect 27387 3516 27399 3519
rect 27430 3516 27436 3528
rect 27387 3488 27436 3516
rect 27387 3485 27399 3488
rect 27341 3479 27399 3485
rect 27430 3476 27436 3488
rect 27488 3476 27494 3528
rect 27985 3519 28043 3525
rect 27985 3485 27997 3519
rect 28031 3516 28043 3519
rect 28074 3516 28080 3528
rect 28031 3488 28080 3516
rect 28031 3485 28043 3488
rect 27985 3479 28043 3485
rect 28074 3476 28080 3488
rect 28132 3476 28138 3528
rect 28350 3476 28356 3528
rect 28408 3516 28414 3528
rect 28445 3519 28503 3525
rect 28445 3516 28457 3519
rect 28408 3488 28457 3516
rect 28408 3476 28414 3488
rect 28445 3485 28457 3488
rect 28491 3485 28503 3519
rect 28445 3479 28503 3485
rect 29270 3476 29276 3528
rect 29328 3516 29334 3528
rect 29549 3519 29607 3525
rect 29549 3516 29561 3519
rect 29328 3488 29561 3516
rect 29328 3476 29334 3488
rect 29549 3485 29561 3488
rect 29595 3485 29607 3519
rect 29549 3479 29607 3485
rect 30466 3476 30472 3528
rect 30524 3516 30530 3528
rect 30837 3519 30895 3525
rect 30837 3516 30849 3519
rect 30524 3488 30849 3516
rect 30524 3476 30530 3488
rect 30837 3485 30849 3488
rect 30883 3485 30895 3519
rect 30837 3479 30895 3485
rect 31018 3476 31024 3528
rect 31076 3516 31082 3528
rect 31481 3519 31539 3525
rect 31481 3516 31493 3519
rect 31076 3488 31493 3516
rect 31076 3476 31082 3488
rect 31481 3485 31493 3488
rect 31527 3485 31539 3519
rect 31481 3479 31539 3485
rect 31938 3476 31944 3528
rect 31996 3516 32002 3528
rect 32125 3519 32183 3525
rect 32125 3516 32137 3519
rect 31996 3488 32137 3516
rect 31996 3476 32002 3488
rect 32125 3485 32137 3488
rect 32171 3485 32183 3519
rect 32125 3479 32183 3485
rect 33045 3519 33103 3525
rect 33045 3485 33057 3519
rect 33091 3516 33103 3519
rect 33134 3516 33140 3528
rect 33091 3488 33140 3516
rect 33091 3485 33103 3488
rect 33045 3479 33103 3485
rect 33134 3476 33140 3488
rect 33192 3476 33198 3528
rect 34606 3476 34612 3528
rect 34664 3516 34670 3528
rect 34701 3519 34759 3525
rect 34701 3516 34713 3519
rect 34664 3488 34713 3516
rect 34664 3476 34670 3488
rect 34701 3485 34713 3488
rect 34747 3485 34759 3519
rect 35342 3516 35348 3528
rect 35303 3488 35348 3516
rect 34701 3479 34759 3485
rect 35342 3476 35348 3488
rect 35400 3476 35406 3528
rect 35802 3476 35808 3528
rect 35860 3516 35866 3528
rect 35989 3519 36047 3525
rect 35989 3516 36001 3519
rect 35860 3488 36001 3516
rect 35860 3476 35866 3488
rect 35989 3485 36001 3488
rect 36035 3485 36047 3519
rect 35989 3479 36047 3485
rect 36170 3476 36176 3528
rect 36228 3516 36234 3528
rect 36633 3519 36691 3525
rect 36633 3516 36645 3519
rect 36228 3488 36645 3516
rect 36228 3476 36234 3488
rect 36633 3485 36645 3488
rect 36679 3485 36691 3519
rect 36633 3479 36691 3485
rect 36998 3476 37004 3528
rect 37056 3516 37062 3528
rect 37277 3519 37335 3525
rect 37277 3516 37289 3519
rect 37056 3488 37289 3516
rect 37056 3476 37062 3488
rect 37277 3485 37289 3488
rect 37323 3485 37335 3519
rect 38194 3516 38200 3528
rect 38155 3488 38200 3516
rect 37277 3479 37335 3485
rect 38194 3476 38200 3488
rect 38252 3476 38258 3528
rect 39114 3516 39120 3528
rect 39075 3488 39120 3516
rect 39114 3476 39120 3488
rect 39172 3476 39178 3528
rect 40310 3516 40316 3528
rect 40271 3488 40316 3516
rect 40310 3476 40316 3488
rect 40368 3476 40374 3528
rect 41230 3516 41236 3528
rect 41191 3488 41236 3516
rect 41230 3476 41236 3488
rect 41288 3476 41294 3528
rect 41877 3519 41935 3525
rect 41877 3516 41889 3519
rect 41386 3488 41889 3516
rect 35250 3448 35256 3460
rect 11900 3420 35256 3448
rect 35250 3408 35256 3420
rect 35308 3408 35314 3460
rect 35894 3408 35900 3460
rect 35952 3448 35958 3460
rect 40402 3448 40408 3460
rect 35952 3420 40408 3448
rect 35952 3408 35958 3420
rect 40402 3408 40408 3420
rect 40460 3408 40466 3460
rect 8018 3380 8024 3392
rect 6380 3352 8024 3380
rect 5261 3343 5319 3349
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 9490 3340 9496 3392
rect 9548 3340 9554 3392
rect 9766 3340 9772 3392
rect 9824 3380 9830 3392
rect 10134 3380 10140 3392
rect 9824 3352 10140 3380
rect 9824 3340 9830 3352
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 10502 3340 10508 3392
rect 10560 3380 10566 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 10560 3352 14197 3380
rect 10560 3340 10566 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 14185 3343 14243 3349
rect 24210 3340 24216 3392
rect 24268 3380 24274 3392
rect 31110 3380 31116 3392
rect 24268 3352 31116 3380
rect 24268 3340 24274 3352
rect 31110 3340 31116 3352
rect 31168 3340 31174 3392
rect 36078 3340 36084 3392
rect 36136 3380 36142 3392
rect 41386 3380 41414 3488
rect 41877 3485 41889 3488
rect 41923 3485 41935 3519
rect 42150 3516 42156 3528
rect 42111 3488 42156 3516
rect 41877 3479 41935 3485
rect 42150 3476 42156 3488
rect 42208 3476 42214 3528
rect 42981 3519 43039 3525
rect 42981 3485 42993 3519
rect 43027 3516 43039 3519
rect 43070 3516 43076 3528
rect 43027 3488 43076 3516
rect 43027 3485 43039 3488
rect 42981 3479 43039 3485
rect 43070 3476 43076 3488
rect 43128 3476 43134 3528
rect 43809 3519 43867 3525
rect 43809 3485 43821 3519
rect 43855 3485 43867 3519
rect 43809 3479 43867 3485
rect 44453 3519 44511 3525
rect 44453 3485 44465 3519
rect 44499 3516 44511 3519
rect 45002 3516 45008 3528
rect 44499 3488 45008 3516
rect 44499 3485 44511 3488
rect 44453 3479 44511 3485
rect 36136 3352 41414 3380
rect 43824 3380 43852 3479
rect 45002 3476 45008 3488
rect 45060 3476 45066 3528
rect 45278 3525 45284 3528
rect 45276 3516 45284 3525
rect 45239 3488 45284 3516
rect 45276 3479 45284 3488
rect 45278 3476 45284 3479
rect 45336 3476 45342 3528
rect 45388 3525 45416 3692
rect 45462 3680 45468 3692
rect 45520 3680 45526 3732
rect 45830 3680 45836 3732
rect 45888 3720 45894 3732
rect 47486 3720 47492 3732
rect 45888 3692 47492 3720
rect 45888 3680 45894 3692
rect 47486 3680 47492 3692
rect 47544 3680 47550 3732
rect 46753 3655 46811 3661
rect 46753 3621 46765 3655
rect 46799 3652 46811 3655
rect 49142 3652 49148 3664
rect 46799 3624 49148 3652
rect 46799 3621 46811 3624
rect 46753 3615 46811 3621
rect 49142 3612 49148 3624
rect 49200 3612 49206 3664
rect 47397 3587 47455 3593
rect 47397 3553 47409 3587
rect 47443 3584 47455 3587
rect 48958 3584 48964 3596
rect 47443 3556 48964 3584
rect 47443 3553 47455 3556
rect 47397 3547 47455 3553
rect 48958 3544 48964 3556
rect 49016 3544 49022 3596
rect 45373 3519 45431 3525
rect 45373 3485 45385 3519
rect 45419 3485 45431 3519
rect 45646 3516 45652 3528
rect 45607 3488 45652 3516
rect 45373 3479 45431 3485
rect 45646 3476 45652 3488
rect 45704 3476 45710 3528
rect 47857 3519 47915 3525
rect 47857 3485 47869 3519
rect 47903 3485 47915 3519
rect 47857 3479 47915 3485
rect 45465 3451 45523 3457
rect 45465 3417 45477 3451
rect 45511 3448 45523 3451
rect 45830 3448 45836 3460
rect 45511 3420 45836 3448
rect 45511 3417 45523 3420
rect 45465 3411 45523 3417
rect 45830 3408 45836 3420
rect 45888 3408 45894 3460
rect 45370 3380 45376 3392
rect 43824 3352 45376 3380
rect 36136 3340 36142 3352
rect 45370 3340 45376 3352
rect 45428 3340 45434 3392
rect 45554 3340 45560 3392
rect 45612 3380 45618 3392
rect 47872 3380 47900 3479
rect 45612 3352 47900 3380
rect 48041 3383 48099 3389
rect 45612 3340 45618 3352
rect 48041 3349 48053 3383
rect 48087 3380 48099 3383
rect 49510 3380 49516 3392
rect 48087 3352 49516 3380
rect 48087 3349 48099 3352
rect 48041 3343 48099 3349
rect 49510 3340 49516 3352
rect 49568 3340 49574 3392
rect 661 3315 719 3321
rect 661 3281 673 3315
rect 707 3312 719 3315
rect 934 3312 940 3324
rect 707 3284 940 3312
rect 707 3281 719 3284
rect 661 3275 719 3281
rect 934 3272 940 3284
rect 992 3272 998 3324
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 1394 3136 1400 3188
rect 1452 3176 1458 3188
rect 2774 3176 2780 3188
rect 1452 3148 2780 3176
rect 1452 3136 1458 3148
rect 2774 3136 2780 3148
rect 2832 3136 2838 3188
rect 2866 3136 2872 3188
rect 2924 3136 2930 3188
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3142 3176 3148 3188
rect 3099 3148 3148 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 3694 3176 3700 3188
rect 3655 3148 3700 3176
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 3878 3136 3884 3188
rect 3936 3136 3942 3188
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 4801 3179 4859 3185
rect 4801 3176 4813 3179
rect 4488 3148 4813 3176
rect 4488 3136 4494 3148
rect 4801 3145 4813 3148
rect 4847 3145 4859 3179
rect 4801 3139 4859 3145
rect 5353 3179 5411 3185
rect 5353 3145 5365 3179
rect 5399 3176 5411 3179
rect 6730 3176 6736 3188
rect 5399 3148 6736 3176
rect 5399 3145 5411 3148
rect 5353 3139 5411 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 7282 3176 7288 3188
rect 7243 3148 7288 3176
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 9582 3176 9588 3188
rect 7883 3148 9588 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 9674 3136 9680 3188
rect 9732 3136 9738 3188
rect 10042 3136 10048 3188
rect 10100 3176 10106 3188
rect 12342 3176 12348 3188
rect 10100 3148 12348 3176
rect 10100 3136 10106 3148
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12986 3176 12992 3188
rect 12636 3148 12992 3176
rect 1762 3068 1768 3120
rect 1820 3108 1826 3120
rect 2130 3108 2136 3120
rect 1820 3080 2136 3108
rect 1820 3068 1826 3080
rect 2130 3068 2136 3080
rect 2188 3068 2194 3120
rect 2222 3068 2228 3120
rect 2280 3108 2286 3120
rect 2593 3111 2651 3117
rect 2593 3108 2605 3111
rect 2280 3080 2605 3108
rect 2280 3068 2286 3080
rect 2593 3077 2605 3080
rect 2639 3077 2651 3111
rect 2884 3108 2912 3136
rect 2593 3071 2651 3077
rect 2792 3080 2912 3108
rect 106 3000 112 3052
rect 164 3040 170 3052
rect 1489 3043 1547 3049
rect 1489 3040 1501 3043
rect 164 3012 1501 3040
rect 164 3000 170 3012
rect 1489 3009 1501 3012
rect 1535 3040 1547 3043
rect 1670 3040 1676 3052
rect 1535 3012 1676 3040
rect 1535 3009 1547 3012
rect 1489 3003 1547 3009
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 2792 3049 2820 3080
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 2777 3003 2835 3009
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 3896 3049 3924 3136
rect 4157 3111 4215 3117
rect 4157 3077 4169 3111
rect 4203 3108 4215 3111
rect 4890 3108 4896 3120
rect 4203 3080 4896 3108
rect 4203 3077 4215 3080
rect 4157 3071 4215 3077
rect 4890 3068 4896 3080
rect 4948 3068 4954 3120
rect 5813 3111 5871 3117
rect 5813 3077 5825 3111
rect 5859 3108 5871 3111
rect 6362 3108 6368 3120
rect 5859 3080 6368 3108
rect 5859 3077 5871 3080
rect 5813 3071 5871 3077
rect 6362 3068 6368 3080
rect 6420 3068 6426 3120
rect 8757 3111 8815 3117
rect 8757 3077 8769 3111
rect 8803 3108 8815 3111
rect 9692 3108 9720 3136
rect 8803 3080 9720 3108
rect 8803 3077 8815 3080
rect 8757 3071 8815 3077
rect 3864 3043 3924 3049
rect 2924 3012 2969 3040
rect 2924 3000 2930 3012
rect 3864 3009 3876 3043
rect 3910 3012 3924 3043
rect 3910 3009 3922 3012
rect 3864 3003 3922 3009
rect 4246 3000 4252 3052
rect 4304 3040 4310 3052
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 4304 3012 4629 3040
rect 4304 3000 4310 3012
rect 4617 3009 4629 3012
rect 4663 3009 4675 3043
rect 5534 3040 5540 3052
rect 5495 3012 5540 3040
rect 4617 3003 4675 3009
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 6273 3043 6331 3049
rect 6273 3040 6285 3043
rect 5960 3012 6285 3040
rect 5960 3000 5966 3012
rect 6273 3009 6285 3012
rect 6319 3009 6331 3043
rect 6638 3040 6644 3052
rect 6599 3012 6644 3040
rect 6273 3003 6331 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3040 6791 3043
rect 7101 3043 7159 3049
rect 6779 3012 7052 3040
rect 6779 3009 6791 3012
rect 6733 3003 6791 3009
rect 845 2975 903 2981
rect 845 2941 857 2975
rect 891 2972 903 2975
rect 1762 2972 1768 2984
rect 891 2944 1768 2972
rect 891 2941 903 2944
rect 845 2935 903 2941
rect 1762 2932 1768 2944
rect 1820 2932 1826 2984
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2972 2099 2975
rect 2087 2944 3372 2972
rect 2087 2941 2099 2944
rect 2041 2935 2099 2941
rect 566 2864 572 2916
rect 624 2904 630 2916
rect 3344 2904 3372 2944
rect 3418 2932 3424 2984
rect 3476 2972 3482 2984
rect 3973 2975 4031 2981
rect 3973 2972 3985 2975
rect 3476 2944 3985 2972
rect 3476 2932 3482 2944
rect 3973 2941 3985 2944
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 4338 2972 4344 2984
rect 4212 2944 4344 2972
rect 4212 2932 4218 2944
rect 4338 2932 4344 2944
rect 4396 2932 4402 2984
rect 4890 2932 4896 2984
rect 4948 2972 4954 2984
rect 5258 2972 5264 2984
rect 4948 2944 5264 2972
rect 4948 2932 4954 2944
rect 5258 2932 5264 2944
rect 5316 2932 5322 2984
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 6454 2972 6460 2984
rect 5767 2944 6460 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 6454 2932 6460 2944
rect 6512 2932 6518 2984
rect 6914 2932 6920 2984
rect 6972 2932 6978 2984
rect 3694 2904 3700 2916
rect 624 2876 2084 2904
rect 3344 2876 3700 2904
rect 624 2864 630 2876
rect 2056 2848 2084 2876
rect 3694 2864 3700 2876
rect 3752 2864 3758 2916
rect 3878 2864 3884 2916
rect 3936 2904 3942 2916
rect 5166 2904 5172 2916
rect 3936 2876 5172 2904
rect 3936 2864 3942 2876
rect 5166 2864 5172 2876
rect 5224 2864 5230 2916
rect 2038 2796 2044 2848
rect 2096 2796 2102 2848
rect 2682 2836 2688 2848
rect 2643 2808 2688 2836
rect 2682 2796 2688 2808
rect 2740 2796 2746 2848
rect 3970 2836 3976 2848
rect 3931 2808 3976 2836
rect 3970 2796 3976 2808
rect 4028 2796 4034 2848
rect 5626 2836 5632 2848
rect 5587 2808 5632 2836
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 6362 2836 6368 2848
rect 6323 2808 6368 2836
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 6454 2796 6460 2848
rect 6512 2836 6518 2848
rect 6932 2836 6960 2932
rect 7024 2904 7052 3012
rect 7101 3009 7113 3043
rect 7147 3040 7159 3043
rect 8202 3040 8208 3052
rect 7147 3012 8208 3040
rect 7147 3009 7159 3012
rect 7101 3003 7159 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3040 8539 3043
rect 9030 3040 9036 3052
rect 8527 3012 9036 3040
rect 8527 3009 8539 3012
rect 8481 3003 8539 3009
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 9306 3040 9312 3052
rect 9267 3012 9312 3040
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3040 10011 3043
rect 10042 3040 10048 3052
rect 9999 3012 10048 3040
rect 9999 3009 10011 3012
rect 9953 3003 10011 3009
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3009 10287 3043
rect 10229 3003 10287 3009
rect 7466 2932 7472 2984
rect 7524 2972 7530 2984
rect 8110 2972 8116 2984
rect 7524 2944 8116 2972
rect 7524 2932 7530 2944
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 8386 2932 8392 2984
rect 8444 2972 8450 2984
rect 8573 2975 8631 2981
rect 8573 2972 8585 2975
rect 8444 2944 8585 2972
rect 8444 2932 8450 2944
rect 8573 2941 8585 2944
rect 8619 2941 8631 2975
rect 10134 2972 10140 2984
rect 10095 2944 10140 2972
rect 8573 2935 8631 2941
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 7098 2904 7104 2916
rect 7024 2876 7104 2904
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 7558 2864 7564 2916
rect 7616 2904 7622 2916
rect 8202 2904 8208 2916
rect 7616 2876 8208 2904
rect 7616 2864 7622 2876
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 8297 2907 8355 2913
rect 8297 2873 8309 2907
rect 8343 2904 8355 2907
rect 10244 2904 10272 3003
rect 10594 3000 10600 3052
rect 10652 3040 10658 3052
rect 10778 3040 10784 3052
rect 10652 3012 10784 3040
rect 10652 3000 10658 3012
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 10870 3000 10876 3052
rect 10928 3040 10934 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10928 3012 10977 3040
rect 10928 3000 10934 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11422 3000 11428 3052
rect 11480 3040 11486 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11480 3012 11529 3040
rect 11480 3000 11486 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 12342 3000 12348 3052
rect 12400 3040 12406 3052
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 12400 3012 12449 3040
rect 12400 3000 12406 3012
rect 12437 3009 12449 3012
rect 12483 3040 12495 3043
rect 12636 3040 12664 3148
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13262 3136 13268 3188
rect 13320 3176 13326 3188
rect 13357 3179 13415 3185
rect 13357 3176 13369 3179
rect 13320 3148 13369 3176
rect 13320 3136 13326 3148
rect 13357 3145 13369 3148
rect 13403 3145 13415 3179
rect 13357 3139 13415 3145
rect 14093 3179 14151 3185
rect 14093 3145 14105 3179
rect 14139 3176 14151 3179
rect 14642 3176 14648 3188
rect 14139 3148 14648 3176
rect 14139 3145 14151 3148
rect 14093 3139 14151 3145
rect 14642 3136 14648 3148
rect 14700 3136 14706 3188
rect 20346 3176 20352 3188
rect 20307 3148 20352 3176
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 24210 3176 24216 3188
rect 24171 3148 24216 3176
rect 24210 3136 24216 3148
rect 24268 3136 24274 3188
rect 28534 3176 28540 3188
rect 28495 3148 28540 3176
rect 28534 3136 28540 3148
rect 28592 3136 28598 3188
rect 28905 3179 28963 3185
rect 28905 3145 28917 3179
rect 28951 3176 28963 3179
rect 30190 3176 30196 3188
rect 28951 3148 30196 3176
rect 28951 3145 28963 3148
rect 28905 3139 28963 3145
rect 30190 3136 30196 3148
rect 30248 3136 30254 3188
rect 30558 3136 30564 3188
rect 30616 3176 30622 3188
rect 30837 3179 30895 3185
rect 30837 3176 30849 3179
rect 30616 3148 30849 3176
rect 30616 3136 30622 3148
rect 30837 3145 30849 3148
rect 30883 3145 30895 3179
rect 30837 3139 30895 3145
rect 31110 3136 31116 3188
rect 31168 3176 31174 3188
rect 35894 3176 35900 3188
rect 31168 3148 35900 3176
rect 31168 3136 31174 3148
rect 35894 3136 35900 3148
rect 35952 3136 35958 3188
rect 36078 3176 36084 3188
rect 36039 3148 36084 3176
rect 36078 3136 36084 3148
rect 36136 3136 36142 3188
rect 47118 3176 47124 3188
rect 41386 3148 47124 3176
rect 12713 3111 12771 3117
rect 12713 3077 12725 3111
rect 12759 3108 12771 3111
rect 14458 3108 14464 3120
rect 12759 3080 14464 3108
rect 12759 3077 12771 3080
rect 12713 3071 12771 3077
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 18506 3108 18512 3120
rect 18467 3080 18512 3108
rect 18506 3068 18512 3080
rect 18564 3068 18570 3120
rect 20162 3068 20168 3120
rect 20220 3108 20226 3120
rect 20257 3111 20315 3117
rect 20257 3108 20269 3111
rect 20220 3080 20269 3108
rect 20220 3068 20226 3080
rect 20257 3077 20269 3080
rect 20303 3077 20315 3111
rect 22278 3108 22284 3120
rect 22239 3080 22284 3108
rect 20257 3071 20315 3077
rect 22278 3068 22284 3080
rect 22336 3068 22342 3120
rect 22465 3111 22523 3117
rect 22465 3077 22477 3111
rect 22511 3108 22523 3111
rect 22511 3080 27108 3108
rect 22511 3077 22523 3080
rect 22465 3071 22523 3077
rect 12483 3012 12664 3040
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 13262 3000 13268 3052
rect 13320 3040 13326 3052
rect 13909 3043 13967 3049
rect 13909 3040 13921 3043
rect 13320 3012 13921 3040
rect 13320 3000 13326 3012
rect 13909 3009 13921 3012
rect 13955 3009 13967 3043
rect 13909 3003 13967 3009
rect 14921 3043 14979 3049
rect 14921 3009 14933 3043
rect 14967 3040 14979 3043
rect 15838 3040 15844 3052
rect 14967 3012 15844 3040
rect 14967 3009 14979 3012
rect 14921 3003 14979 3009
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 23750 3000 23756 3052
rect 23808 3040 23814 3052
rect 24121 3043 24179 3049
rect 24121 3040 24133 3043
rect 23808 3012 24133 3040
rect 23808 3000 23814 3012
rect 24121 3009 24133 3012
rect 24167 3009 24179 3043
rect 27080 3040 27108 3080
rect 27982 3068 27988 3120
rect 28040 3108 28046 3120
rect 28997 3111 29055 3117
rect 28997 3108 29009 3111
rect 28040 3080 29009 3108
rect 28040 3068 28046 3080
rect 28997 3077 29009 3080
rect 29043 3077 29055 3111
rect 29822 3108 29828 3120
rect 29783 3080 29828 3108
rect 28997 3071 29055 3077
rect 29822 3068 29828 3080
rect 29880 3068 29886 3120
rect 35250 3068 35256 3120
rect 35308 3108 35314 3120
rect 35345 3111 35403 3117
rect 35345 3108 35357 3111
rect 35308 3080 35357 3108
rect 35308 3068 35314 3080
rect 35345 3077 35357 3080
rect 35391 3108 35403 3111
rect 35710 3108 35716 3120
rect 35391 3080 35716 3108
rect 35391 3077 35403 3080
rect 35345 3071 35403 3077
rect 35710 3068 35716 3080
rect 35768 3108 35774 3120
rect 35989 3111 36047 3117
rect 35989 3108 36001 3111
rect 35768 3080 36001 3108
rect 35768 3068 35774 3080
rect 35989 3077 36001 3080
rect 36035 3077 36047 3111
rect 35989 3071 36047 3077
rect 24121 3003 24179 3009
rect 24412 3012 26924 3040
rect 27080 3012 29960 3040
rect 11790 2972 11796 2984
rect 8343 2876 10272 2904
rect 10336 2944 11560 2972
rect 11751 2944 11796 2972
rect 8343 2873 8355 2876
rect 8297 2867 8355 2873
rect 6512 2808 6960 2836
rect 6512 2796 6518 2808
rect 7006 2796 7012 2848
rect 7064 2836 7070 2848
rect 8757 2839 8815 2845
rect 7064 2808 7109 2836
rect 7064 2796 7070 2808
rect 8757 2805 8769 2839
rect 8803 2836 8815 2839
rect 9122 2836 9128 2848
rect 8803 2808 9128 2836
rect 8803 2805 8815 2808
rect 8757 2799 8815 2805
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 9306 2796 9312 2848
rect 9364 2836 9370 2848
rect 9674 2836 9680 2848
rect 9364 2808 9680 2836
rect 9364 2796 9370 2808
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 9769 2839 9827 2845
rect 9769 2805 9781 2839
rect 9815 2836 9827 2839
rect 9950 2836 9956 2848
rect 9815 2808 9956 2836
rect 9815 2805 9827 2808
rect 9769 2799 9827 2805
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 10229 2839 10287 2845
rect 10229 2805 10241 2839
rect 10275 2836 10287 2839
rect 10336 2836 10364 2944
rect 11532 2916 11560 2944
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 16025 2975 16083 2981
rect 16025 2972 16037 2975
rect 14240 2944 16037 2972
rect 14240 2932 14246 2944
rect 16025 2941 16037 2944
rect 16071 2941 16083 2975
rect 16025 2935 16083 2941
rect 18693 2975 18751 2981
rect 18693 2941 18705 2975
rect 18739 2972 18751 2975
rect 24412 2972 24440 3012
rect 18739 2944 24440 2972
rect 18739 2941 18751 2944
rect 18693 2935 18751 2941
rect 24486 2932 24492 2984
rect 24544 2972 24550 2984
rect 25409 2975 25467 2981
rect 25409 2972 25421 2975
rect 24544 2944 25421 2972
rect 24544 2932 24550 2944
rect 25409 2941 25421 2944
rect 25455 2941 25467 2975
rect 25409 2935 25467 2941
rect 11514 2864 11520 2916
rect 11572 2864 11578 2916
rect 14734 2904 14740 2916
rect 14695 2876 14740 2904
rect 14734 2864 14740 2876
rect 14792 2864 14798 2916
rect 14844 2876 15516 2904
rect 10275 2808 10364 2836
rect 10781 2839 10839 2845
rect 10275 2805 10287 2808
rect 10229 2799 10287 2805
rect 10781 2805 10793 2839
rect 10827 2836 10839 2839
rect 10870 2836 10876 2848
rect 10827 2808 10876 2836
rect 10827 2805 10839 2808
rect 10781 2799 10839 2805
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 11238 2796 11244 2848
rect 11296 2836 11302 2848
rect 12434 2836 12440 2848
rect 11296 2808 12440 2836
rect 11296 2796 11302 2808
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 14274 2796 14280 2848
rect 14332 2836 14338 2848
rect 14844 2836 14872 2876
rect 14332 2808 14872 2836
rect 14332 2796 14338 2808
rect 14918 2796 14924 2848
rect 14976 2836 14982 2848
rect 15381 2839 15439 2845
rect 15381 2836 15393 2839
rect 14976 2808 15393 2836
rect 14976 2796 14982 2808
rect 15381 2805 15393 2808
rect 15427 2805 15439 2839
rect 15488 2836 15516 2876
rect 15746 2864 15752 2916
rect 15804 2904 15810 2916
rect 17313 2907 17371 2913
rect 17313 2904 17325 2907
rect 15804 2876 17325 2904
rect 15804 2864 15810 2876
rect 17313 2873 17325 2876
rect 17359 2873 17371 2907
rect 17313 2867 17371 2873
rect 18138 2864 18144 2916
rect 18196 2904 18202 2916
rect 19153 2907 19211 2913
rect 19153 2904 19165 2907
rect 18196 2876 19165 2904
rect 18196 2864 18202 2876
rect 19153 2873 19165 2876
rect 19199 2873 19211 2907
rect 19153 2867 19211 2873
rect 19978 2864 19984 2916
rect 20036 2904 20042 2916
rect 20901 2907 20959 2913
rect 20901 2904 20913 2907
rect 20036 2876 20913 2904
rect 20036 2864 20042 2876
rect 20901 2873 20913 2876
rect 20947 2873 20959 2907
rect 20901 2867 20959 2873
rect 21726 2864 21732 2916
rect 21784 2904 21790 2916
rect 22925 2907 22983 2913
rect 22925 2904 22937 2907
rect 21784 2876 22937 2904
rect 21784 2864 21790 2876
rect 22925 2873 22937 2876
rect 22971 2873 22983 2907
rect 22925 2867 22983 2873
rect 23566 2864 23572 2916
rect 23624 2904 23630 2916
rect 24765 2907 24823 2913
rect 24765 2904 24777 2907
rect 23624 2876 24777 2904
rect 23624 2864 23630 2876
rect 24765 2873 24777 2876
rect 24811 2873 24823 2907
rect 24765 2867 24823 2873
rect 25314 2864 25320 2916
rect 25372 2904 25378 2916
rect 26053 2907 26111 2913
rect 26053 2904 26065 2907
rect 25372 2876 26065 2904
rect 25372 2864 25378 2876
rect 26053 2873 26065 2876
rect 26099 2873 26111 2907
rect 26896 2904 26924 3012
rect 28810 2932 28816 2984
rect 28868 2972 28874 2984
rect 29089 2975 29147 2981
rect 29089 2972 29101 2975
rect 28868 2944 29101 2972
rect 28868 2932 28874 2944
rect 29089 2941 29101 2944
rect 29135 2941 29147 2975
rect 29932 2972 29960 3012
rect 30374 3000 30380 3052
rect 30432 3040 30438 3052
rect 30432 3012 30590 3040
rect 30432 3000 30438 3012
rect 40678 3000 40684 3052
rect 40736 3040 40742 3052
rect 41386 3040 41414 3148
rect 47118 3136 47124 3148
rect 47176 3136 47182 3188
rect 47302 3136 47308 3188
rect 47360 3176 47366 3188
rect 48406 3176 48412 3188
rect 47360 3148 48412 3176
rect 47360 3136 47366 3148
rect 48406 3136 48412 3148
rect 48464 3136 48470 3188
rect 41690 3068 41696 3120
rect 41748 3108 41754 3120
rect 45554 3108 45560 3120
rect 41748 3080 45560 3108
rect 41748 3068 41754 3080
rect 45554 3068 45560 3080
rect 45612 3068 45618 3120
rect 49050 3108 49056 3120
rect 46308 3080 49056 3108
rect 40736 3012 41414 3040
rect 41877 3043 41935 3049
rect 40736 3000 40742 3012
rect 41877 3009 41889 3043
rect 41923 3040 41935 3043
rect 45462 3040 45468 3052
rect 41923 3012 45468 3040
rect 41923 3009 41935 3012
rect 41877 3003 41935 3009
rect 45462 3000 45468 3012
rect 45520 3000 45526 3052
rect 46308 3049 46336 3080
rect 49050 3068 49056 3080
rect 49108 3068 49114 3120
rect 46293 3043 46351 3049
rect 46293 3009 46305 3043
rect 46339 3009 46351 3043
rect 46293 3003 46351 3009
rect 46753 3043 46811 3049
rect 46753 3009 46765 3043
rect 46799 3009 46811 3043
rect 46753 3003 46811 3009
rect 47857 3043 47915 3049
rect 47857 3009 47869 3043
rect 47903 3009 47915 3043
rect 47857 3003 47915 3009
rect 30650 2972 30656 2984
rect 29932 2944 30656 2972
rect 29089 2935 29147 2941
rect 30650 2932 30656 2944
rect 30708 2932 30714 2984
rect 31202 2932 31208 2984
rect 31260 2932 31266 2984
rect 33410 2932 33416 2984
rect 33468 2972 33474 2984
rect 34057 2975 34115 2981
rect 34057 2972 34069 2975
rect 33468 2944 34069 2972
rect 33468 2932 33474 2944
rect 34057 2941 34069 2944
rect 34103 2941 34115 2975
rect 34057 2935 34115 2941
rect 37918 2932 37924 2984
rect 37976 2972 37982 2984
rect 38565 2975 38623 2981
rect 38565 2972 38577 2975
rect 37976 2944 38577 2972
rect 37976 2932 37982 2944
rect 38565 2941 38577 2944
rect 38611 2941 38623 2975
rect 38565 2935 38623 2941
rect 44174 2932 44180 2984
rect 44232 2972 44238 2984
rect 46768 2972 46796 3003
rect 44232 2944 46796 2972
rect 44232 2932 44238 2944
rect 40862 2904 40868 2916
rect 26896 2876 40868 2904
rect 26053 2867 26111 2873
rect 40862 2864 40868 2876
rect 40920 2904 40926 2916
rect 47872 2904 47900 3003
rect 49602 2904 49608 2916
rect 40920 2876 47900 2904
rect 47964 2876 49608 2904
rect 40920 2864 40926 2876
rect 16669 2839 16727 2845
rect 16669 2836 16681 2839
rect 15488 2808 16681 2836
rect 15381 2799 15439 2805
rect 16669 2805 16681 2808
rect 16715 2805 16727 2839
rect 16669 2799 16727 2805
rect 26510 2796 26516 2848
rect 26568 2836 26574 2848
rect 26973 2839 27031 2845
rect 26973 2836 26985 2839
rect 26568 2808 26985 2836
rect 26568 2796 26574 2808
rect 26973 2805 26985 2808
rect 27019 2805 27031 2839
rect 26973 2799 27031 2805
rect 27154 2796 27160 2848
rect 27212 2836 27218 2848
rect 27617 2839 27675 2845
rect 27617 2836 27629 2839
rect 27212 2808 27629 2836
rect 27212 2796 27218 2808
rect 27617 2805 27629 2808
rect 27663 2805 27675 2839
rect 27617 2799 27675 2805
rect 31386 2796 31392 2848
rect 31444 2836 31450 2848
rect 32125 2839 32183 2845
rect 32125 2836 32137 2839
rect 31444 2808 32137 2836
rect 31444 2796 31450 2808
rect 32125 2805 32137 2808
rect 32171 2805 32183 2839
rect 32125 2799 32183 2805
rect 32214 2796 32220 2848
rect 32272 2836 32278 2848
rect 32769 2839 32827 2845
rect 32769 2836 32781 2839
rect 32272 2808 32781 2836
rect 32272 2796 32278 2808
rect 32769 2805 32781 2808
rect 32815 2805 32827 2839
rect 32769 2799 32827 2805
rect 32858 2796 32864 2848
rect 32916 2836 32922 2848
rect 33413 2839 33471 2845
rect 33413 2836 33425 2839
rect 32916 2808 33425 2836
rect 32916 2796 32922 2808
rect 33413 2805 33425 2808
rect 33459 2805 33471 2839
rect 33413 2799 33471 2805
rect 34054 2796 34060 2848
rect 34112 2836 34118 2848
rect 34701 2839 34759 2845
rect 34701 2836 34713 2839
rect 34112 2808 34713 2836
rect 34112 2796 34118 2808
rect 34701 2805 34713 2808
rect 34747 2805 34759 2839
rect 34701 2799 34759 2805
rect 36446 2796 36452 2848
rect 36504 2836 36510 2848
rect 37277 2839 37335 2845
rect 37277 2836 37289 2839
rect 36504 2808 37289 2836
rect 36504 2796 36510 2808
rect 37277 2805 37289 2808
rect 37323 2805 37335 2839
rect 37277 2799 37335 2805
rect 37366 2796 37372 2848
rect 37424 2836 37430 2848
rect 37921 2839 37979 2845
rect 37921 2836 37933 2839
rect 37424 2808 37933 2836
rect 37424 2796 37430 2808
rect 37921 2805 37933 2808
rect 37967 2805 37979 2839
rect 37921 2799 37979 2805
rect 38562 2796 38568 2848
rect 38620 2836 38626 2848
rect 39209 2839 39267 2845
rect 39209 2836 39221 2839
rect 38620 2808 39221 2836
rect 38620 2796 38626 2808
rect 39209 2805 39221 2808
rect 39255 2805 39267 2839
rect 39209 2799 39267 2805
rect 39390 2796 39396 2848
rect 39448 2836 39454 2848
rect 39853 2839 39911 2845
rect 39853 2836 39865 2839
rect 39448 2808 39865 2836
rect 39448 2796 39454 2808
rect 39853 2805 39865 2808
rect 39899 2805 39911 2839
rect 39853 2799 39911 2805
rect 40034 2796 40040 2848
rect 40092 2836 40098 2848
rect 40497 2839 40555 2845
rect 40497 2836 40509 2839
rect 40092 2808 40509 2836
rect 40092 2796 40098 2808
rect 40497 2805 40509 2808
rect 40543 2805 40555 2839
rect 40497 2799 40555 2805
rect 40678 2796 40684 2848
rect 40736 2836 40742 2848
rect 41141 2839 41199 2845
rect 41141 2836 41153 2839
rect 40736 2808 41153 2836
rect 40736 2796 40742 2808
rect 41141 2805 41153 2808
rect 41187 2805 41199 2839
rect 41141 2799 41199 2805
rect 41874 2796 41880 2848
rect 41932 2836 41938 2848
rect 42429 2839 42487 2845
rect 42429 2836 42441 2839
rect 41932 2808 42441 2836
rect 41932 2796 41938 2808
rect 42429 2805 42441 2808
rect 42475 2805 42487 2839
rect 42429 2799 42487 2805
rect 42702 2796 42708 2848
rect 42760 2836 42766 2848
rect 43073 2839 43131 2845
rect 43073 2836 43085 2839
rect 42760 2808 43085 2836
rect 42760 2796 42766 2808
rect 43073 2805 43085 2808
rect 43119 2805 43131 2839
rect 43073 2799 43131 2805
rect 43346 2796 43352 2848
rect 43404 2836 43410 2848
rect 43717 2839 43775 2845
rect 43717 2836 43729 2839
rect 43404 2808 43729 2836
rect 43404 2796 43410 2808
rect 43717 2805 43729 2808
rect 43763 2805 43775 2839
rect 43717 2799 43775 2805
rect 43898 2796 43904 2848
rect 43956 2836 43962 2848
rect 44361 2839 44419 2845
rect 44361 2836 44373 2839
rect 43956 2808 44373 2836
rect 43956 2796 43962 2808
rect 44361 2805 44373 2808
rect 44407 2805 44419 2839
rect 44361 2799 44419 2805
rect 44542 2796 44548 2848
rect 44600 2836 44606 2848
rect 45005 2839 45063 2845
rect 45005 2836 45017 2839
rect 44600 2808 45017 2836
rect 44600 2796 44606 2808
rect 45005 2805 45017 2808
rect 45051 2805 45063 2839
rect 45005 2799 45063 2805
rect 46937 2839 46995 2845
rect 46937 2805 46949 2839
rect 46983 2836 46995 2839
rect 47964 2836 47992 2876
rect 49602 2864 49608 2876
rect 49660 2864 49666 2916
rect 46983 2808 47992 2836
rect 48041 2839 48099 2845
rect 46983 2805 46995 2808
rect 46937 2799 46995 2805
rect 48041 2805 48053 2839
rect 48087 2836 48099 2839
rect 49326 2836 49332 2848
rect 48087 2808 49332 2836
rect 48087 2805 48099 2808
rect 48041 2799 48099 2805
rect 49326 2796 49332 2808
rect 49384 2796 49390 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 937 2635 995 2641
rect 937 2601 949 2635
rect 983 2632 995 2635
rect 1486 2632 1492 2644
rect 983 2604 1492 2632
rect 983 2601 995 2604
rect 937 2595 995 2601
rect 1486 2592 1492 2604
rect 1544 2592 1550 2644
rect 2498 2592 2504 2644
rect 2556 2632 2562 2644
rect 2682 2632 2688 2644
rect 2556 2604 2688 2632
rect 2556 2592 2562 2604
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 2866 2632 2872 2644
rect 2823 2604 2872 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 3142 2632 3148 2644
rect 3103 2604 3148 2632
rect 3142 2592 3148 2604
rect 3200 2592 3206 2644
rect 6730 2592 6736 2644
rect 6788 2632 6794 2644
rect 7558 2632 7564 2644
rect 6788 2604 7564 2632
rect 6788 2592 6794 2604
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 7926 2592 7932 2644
rect 7984 2632 7990 2644
rect 7984 2604 9674 2632
rect 7984 2592 7990 2604
rect 8478 2564 8484 2576
rect 1964 2536 8484 2564
rect 1964 2505 1992 2536
rect 8478 2524 8484 2536
rect 8536 2524 8542 2576
rect 8757 2567 8815 2573
rect 8757 2533 8769 2567
rect 8803 2564 8815 2567
rect 9398 2564 9404 2576
rect 8803 2536 9404 2564
rect 8803 2533 8815 2536
rect 8757 2527 8815 2533
rect 9398 2524 9404 2536
rect 9456 2524 9462 2576
rect 9646 2564 9674 2604
rect 10134 2592 10140 2644
rect 10192 2632 10198 2644
rect 13449 2635 13507 2641
rect 13449 2632 13461 2635
rect 10192 2604 13461 2632
rect 10192 2592 10198 2604
rect 13449 2601 13461 2604
rect 13495 2601 13507 2635
rect 14921 2635 14979 2641
rect 14921 2632 14933 2635
rect 13449 2595 13507 2601
rect 13556 2604 14933 2632
rect 9646 2536 10456 2564
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2465 2007 2499
rect 1949 2459 2007 2465
rect 2038 2456 2044 2508
rect 2096 2496 2102 2508
rect 2498 2496 2504 2508
rect 2096 2468 2504 2496
rect 2096 2456 2102 2468
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 3050 2496 3056 2508
rect 3011 2468 3056 2496
rect 3050 2456 3056 2468
rect 3108 2456 3114 2508
rect 7282 2456 7288 2508
rect 7340 2496 7346 2508
rect 9674 2496 9680 2508
rect 7340 2468 9680 2496
rect 7340 2456 7346 2468
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 9858 2456 9864 2508
rect 9916 2496 9922 2508
rect 10318 2496 10324 2508
rect 9916 2468 10324 2496
rect 9916 2456 9922 2468
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 10428 2496 10456 2536
rect 11054 2524 11060 2576
rect 11112 2564 11118 2576
rect 11974 2564 11980 2576
rect 11112 2536 11980 2564
rect 11112 2524 11118 2536
rect 11974 2524 11980 2536
rect 12032 2524 12038 2576
rect 13556 2564 13584 2604
rect 14921 2601 14933 2604
rect 14967 2601 14979 2635
rect 14921 2595 14979 2601
rect 28997 2635 29055 2641
rect 28997 2601 29009 2635
rect 29043 2632 29055 2635
rect 29178 2632 29184 2644
rect 29043 2604 29184 2632
rect 29043 2601 29055 2604
rect 28997 2595 29055 2601
rect 29178 2592 29184 2604
rect 29236 2592 29242 2644
rect 42518 2592 42524 2644
rect 42576 2632 42582 2644
rect 46842 2632 46848 2644
rect 42576 2604 46848 2632
rect 42576 2592 42582 2604
rect 46842 2592 46848 2604
rect 46900 2592 46906 2644
rect 12176 2536 13584 2564
rect 10428 2468 11008 2496
rect 474 2388 480 2440
rect 532 2428 538 2440
rect 842 2428 848 2440
rect 532 2400 848 2428
rect 532 2388 538 2400
rect 842 2388 848 2400
rect 900 2428 906 2440
rect 2225 2431 2283 2437
rect 2225 2428 2237 2431
rect 900 2400 2237 2428
rect 900 2388 906 2400
rect 2225 2397 2237 2400
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 2314 2388 2320 2440
rect 2372 2428 2378 2440
rect 2961 2431 3019 2437
rect 2961 2428 2973 2431
rect 2372 2400 2973 2428
rect 2372 2388 2378 2400
rect 2961 2397 2973 2400
rect 3007 2397 3019 2431
rect 3234 2428 3240 2440
rect 3195 2400 3240 2428
rect 2961 2391 3019 2397
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 4338 2388 4344 2440
rect 4396 2428 4402 2440
rect 5169 2431 5227 2437
rect 5169 2428 5181 2431
rect 4396 2400 5181 2428
rect 4396 2388 4402 2400
rect 5169 2397 5181 2400
rect 5215 2428 5227 2431
rect 6362 2428 6368 2440
rect 5215 2400 6368 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 6914 2428 6920 2440
rect 6840 2400 6920 2428
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 4249 2363 4307 2369
rect 4249 2360 4261 2363
rect 4212 2332 4261 2360
rect 4212 2320 4218 2332
rect 4249 2329 4261 2332
rect 4295 2360 4307 2363
rect 4706 2360 4712 2372
rect 4295 2332 4712 2360
rect 4295 2329 4307 2332
rect 4249 2323 4307 2329
rect 4706 2320 4712 2332
rect 4764 2320 4770 2372
rect 5626 2320 5632 2372
rect 5684 2360 5690 2372
rect 6840 2369 6868 2400
rect 6914 2388 6920 2400
rect 6972 2388 6978 2440
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 8757 2431 8815 2437
rect 8757 2428 8769 2431
rect 8168 2400 8769 2428
rect 8168 2388 8174 2400
rect 8757 2397 8769 2400
rect 8803 2397 8815 2431
rect 8757 2391 8815 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9088 2400 10732 2428
rect 9088 2388 9094 2400
rect 6825 2363 6883 2369
rect 6825 2360 6837 2363
rect 5684 2332 6837 2360
rect 5684 2320 5690 2332
rect 6825 2329 6837 2332
rect 6871 2329 6883 2363
rect 6825 2323 6883 2329
rect 7006 2320 7012 2372
rect 7064 2360 7070 2372
rect 7745 2363 7803 2369
rect 7745 2360 7757 2363
rect 7064 2332 7757 2360
rect 7064 2320 7070 2332
rect 7745 2329 7757 2332
rect 7791 2329 7803 2363
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 7745 2323 7803 2329
rect 7944 2332 9413 2360
rect 2958 2252 2964 2304
rect 3016 2292 3022 2304
rect 3694 2292 3700 2304
rect 3016 2264 3700 2292
rect 3016 2252 3022 2264
rect 3694 2252 3700 2264
rect 3752 2252 3758 2304
rect 4522 2292 4528 2304
rect 4483 2264 4528 2292
rect 4522 2252 4528 2264
rect 4580 2252 4586 2304
rect 5445 2295 5503 2301
rect 5445 2261 5457 2295
rect 5491 2292 5503 2295
rect 6914 2292 6920 2304
rect 5491 2264 6920 2292
rect 5491 2261 5503 2264
rect 5445 2255 5503 2261
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 7098 2292 7104 2304
rect 7059 2264 7104 2292
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 7374 2252 7380 2304
rect 7432 2292 7438 2304
rect 7944 2292 7972 2332
rect 9401 2329 9413 2332
rect 9447 2360 9459 2363
rect 10042 2360 10048 2372
rect 9447 2332 10048 2360
rect 9447 2329 9459 2332
rect 9401 2323 9459 2329
rect 10042 2320 10048 2332
rect 10100 2320 10106 2372
rect 10318 2360 10324 2372
rect 10279 2332 10324 2360
rect 10318 2320 10324 2332
rect 10376 2320 10382 2372
rect 10704 2360 10732 2400
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 10873 2431 10931 2437
rect 10873 2428 10885 2431
rect 10836 2400 10885 2428
rect 10836 2388 10842 2400
rect 10873 2397 10885 2400
rect 10919 2397 10931 2431
rect 10980 2428 11008 2468
rect 11146 2456 11152 2508
rect 11204 2496 11210 2508
rect 11701 2499 11759 2505
rect 11701 2496 11713 2499
rect 11204 2468 11713 2496
rect 11204 2456 11210 2468
rect 11701 2465 11713 2468
rect 11747 2465 11759 2499
rect 11701 2459 11759 2465
rect 11330 2428 11336 2440
rect 10980 2400 11336 2428
rect 10873 2391 10931 2397
rect 11330 2388 11336 2400
rect 11388 2388 11394 2440
rect 11974 2428 11980 2440
rect 11935 2400 11980 2428
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 12176 2360 12204 2536
rect 13998 2524 14004 2576
rect 14056 2564 14062 2576
rect 15565 2567 15623 2573
rect 15565 2564 15577 2567
rect 14056 2536 15577 2564
rect 14056 2524 14062 2536
rect 15565 2533 15577 2536
rect 15611 2533 15623 2567
rect 15565 2527 15623 2533
rect 16666 2524 16672 2576
rect 16724 2564 16730 2576
rect 17313 2567 17371 2573
rect 17313 2564 17325 2567
rect 16724 2536 17325 2564
rect 16724 2524 16730 2536
rect 17313 2533 17325 2536
rect 17359 2533 17371 2567
rect 17313 2527 17371 2533
rect 23842 2524 23848 2576
rect 23900 2564 23906 2576
rect 25041 2567 25099 2573
rect 25041 2564 25053 2567
rect 23900 2536 25053 2564
rect 23900 2524 23906 2536
rect 25041 2533 25053 2536
rect 25087 2533 25099 2567
rect 25041 2527 25099 2533
rect 43254 2524 43260 2576
rect 43312 2564 43318 2576
rect 46750 2564 46756 2576
rect 43312 2536 46756 2564
rect 43312 2524 43318 2536
rect 46750 2524 46756 2536
rect 46808 2524 46814 2576
rect 46937 2567 46995 2573
rect 46937 2533 46949 2567
rect 46983 2564 46995 2567
rect 49418 2564 49424 2576
rect 46983 2536 49424 2564
rect 46983 2533 46995 2536
rect 46937 2527 46995 2533
rect 49418 2524 49424 2536
rect 49476 2524 49482 2576
rect 15378 2496 15384 2508
rect 14384 2468 15384 2496
rect 12342 2388 12348 2440
rect 12400 2428 12406 2440
rect 12437 2431 12495 2437
rect 12437 2428 12449 2431
rect 12400 2400 12449 2428
rect 12400 2388 12406 2400
rect 12437 2397 12449 2400
rect 12483 2428 12495 2431
rect 12526 2428 12532 2440
rect 12483 2400 12532 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 12526 2388 12532 2400
rect 12584 2388 12590 2440
rect 13357 2438 13415 2439
rect 13096 2433 13415 2438
rect 14384 2437 14412 2468
rect 15378 2456 15384 2468
rect 15436 2456 15442 2508
rect 22922 2456 22928 2508
rect 22980 2496 22986 2508
rect 24397 2499 24455 2505
rect 24397 2496 24409 2499
rect 22980 2468 24409 2496
rect 22980 2456 22986 2468
rect 24397 2465 24409 2468
rect 24443 2465 24455 2499
rect 24397 2459 24455 2465
rect 24762 2456 24768 2508
rect 24820 2496 24826 2508
rect 25685 2499 25743 2505
rect 25685 2496 25697 2499
rect 24820 2468 25697 2496
rect 24820 2456 24826 2468
rect 25685 2465 25697 2468
rect 25731 2465 25743 2499
rect 25685 2459 25743 2465
rect 26878 2456 26884 2508
rect 26936 2496 26942 2508
rect 27617 2499 27675 2505
rect 27617 2496 27629 2499
rect 26936 2468 27629 2496
rect 26936 2456 26942 2468
rect 27617 2465 27629 2468
rect 27663 2465 27675 2499
rect 30926 2496 30932 2508
rect 27617 2459 27675 2465
rect 28552 2468 30932 2496
rect 13096 2428 13369 2433
rect 12636 2410 13369 2428
rect 12636 2400 13124 2410
rect 10704 2332 12204 2360
rect 12250 2320 12256 2372
rect 12308 2360 12314 2372
rect 12636 2360 12664 2400
rect 13357 2399 13369 2410
rect 13403 2399 13415 2433
rect 13357 2393 13415 2399
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2397 13599 2431
rect 13541 2391 13599 2397
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2428 15163 2431
rect 15470 2428 15476 2440
rect 15151 2400 15476 2428
rect 15151 2397 15163 2400
rect 15105 2391 15163 2397
rect 12308 2332 12664 2360
rect 12308 2320 12314 2332
rect 12710 2320 12716 2372
rect 12768 2360 12774 2372
rect 12768 2332 12813 2360
rect 12768 2320 12774 2332
rect 7432 2264 7972 2292
rect 8021 2295 8079 2301
rect 7432 2252 7438 2264
rect 8021 2261 8033 2295
rect 8067 2292 8079 2295
rect 9214 2292 9220 2304
rect 8067 2264 9220 2292
rect 8067 2261 8079 2264
rect 8021 2255 8079 2261
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 9674 2292 9680 2304
rect 9635 2264 9680 2292
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 13556 2292 13584 2391
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 15654 2388 15660 2440
rect 15712 2428 15718 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 15712 2400 16681 2428
rect 15712 2388 15718 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 17586 2388 17592 2440
rect 17644 2428 17650 2440
rect 17957 2431 18015 2437
rect 17957 2428 17969 2431
rect 17644 2400 17969 2428
rect 17644 2388 17650 2400
rect 17957 2397 17969 2400
rect 18003 2397 18015 2431
rect 18598 2428 18604 2440
rect 18559 2400 18604 2428
rect 17957 2391 18015 2397
rect 18598 2388 18604 2400
rect 18656 2388 18662 2440
rect 18782 2388 18788 2440
rect 18840 2428 18846 2440
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 18840 2400 19257 2428
rect 18840 2388 18846 2400
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19889 2431 19947 2437
rect 19889 2428 19901 2431
rect 19392 2400 19901 2428
rect 19392 2388 19398 2400
rect 19889 2397 19901 2400
rect 19935 2397 19947 2431
rect 19889 2391 19947 2397
rect 20254 2388 20260 2440
rect 20312 2428 20318 2440
rect 20533 2431 20591 2437
rect 20533 2428 20545 2431
rect 20312 2400 20545 2428
rect 20312 2388 20318 2400
rect 20533 2397 20545 2400
rect 20579 2397 20591 2431
rect 20533 2391 20591 2397
rect 21174 2388 21180 2440
rect 21232 2428 21238 2440
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 21232 2400 21833 2428
rect 21232 2388 21238 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 22094 2388 22100 2440
rect 22152 2428 22158 2440
rect 22465 2431 22523 2437
rect 22465 2428 22477 2431
rect 22152 2400 22477 2428
rect 22152 2388 22158 2400
rect 22465 2397 22477 2400
rect 22511 2397 22523 2431
rect 22465 2391 22523 2397
rect 22646 2388 22652 2440
rect 22704 2428 22710 2440
rect 23201 2431 23259 2437
rect 23201 2428 23213 2431
rect 22704 2400 23213 2428
rect 22704 2388 22710 2400
rect 23201 2397 23213 2400
rect 23247 2397 23259 2431
rect 23201 2391 23259 2397
rect 25774 2388 25780 2440
rect 25832 2428 25838 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 25832 2400 26985 2428
rect 25832 2388 25838 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 27706 2388 27712 2440
rect 27764 2428 27770 2440
rect 28261 2431 28319 2437
rect 28261 2428 28273 2431
rect 27764 2400 28273 2428
rect 27764 2388 27770 2400
rect 28261 2397 28273 2400
rect 28307 2397 28319 2431
rect 28261 2391 28319 2397
rect 17402 2320 17408 2372
rect 17460 2360 17466 2372
rect 28552 2360 28580 2468
rect 30926 2456 30932 2468
rect 30984 2456 30990 2508
rect 41322 2456 41328 2508
rect 41380 2496 41386 2508
rect 41380 2468 46796 2496
rect 41380 2456 41386 2468
rect 29822 2388 29828 2440
rect 29880 2428 29886 2440
rect 30653 2431 30711 2437
rect 30653 2428 30665 2431
rect 29880 2400 30665 2428
rect 29880 2388 29886 2400
rect 30653 2397 30665 2400
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31297 2431 31355 2437
rect 31297 2428 31309 2431
rect 30800 2400 31309 2428
rect 30800 2388 30806 2400
rect 31297 2397 31309 2400
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 31662 2388 31668 2440
rect 31720 2428 31726 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31720 2400 32137 2428
rect 31720 2388 31726 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 32582 2388 32588 2440
rect 32640 2428 32646 2440
rect 32769 2431 32827 2437
rect 32769 2428 32781 2431
rect 32640 2400 32781 2428
rect 32640 2388 32646 2400
rect 32769 2397 32781 2400
rect 32815 2397 32827 2431
rect 33778 2428 33784 2440
rect 33739 2400 33784 2428
rect 32769 2391 32827 2397
rect 33778 2388 33784 2400
rect 33836 2388 33842 2440
rect 34330 2388 34336 2440
rect 34388 2428 34394 2440
rect 34701 2431 34759 2437
rect 34701 2428 34713 2431
rect 34388 2400 34713 2428
rect 34388 2388 34394 2400
rect 34701 2397 34713 2400
rect 34747 2397 34759 2431
rect 34701 2391 34759 2397
rect 34974 2388 34980 2440
rect 35032 2428 35038 2440
rect 35345 2431 35403 2437
rect 35345 2428 35357 2431
rect 35032 2400 35357 2428
rect 35032 2388 35038 2400
rect 35345 2397 35357 2400
rect 35391 2397 35403 2431
rect 35345 2391 35403 2397
rect 35526 2388 35532 2440
rect 35584 2428 35590 2440
rect 35989 2431 36047 2437
rect 35989 2428 36001 2431
rect 35584 2400 36001 2428
rect 35584 2388 35590 2400
rect 35989 2397 36001 2400
rect 36035 2397 36047 2431
rect 35989 2391 36047 2397
rect 36722 2388 36728 2440
rect 36780 2428 36786 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36780 2400 37289 2428
rect 36780 2388 36786 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 37642 2388 37648 2440
rect 37700 2428 37706 2440
rect 37921 2431 37979 2437
rect 37921 2428 37933 2431
rect 37700 2400 37933 2428
rect 37700 2388 37706 2400
rect 37921 2397 37933 2400
rect 37967 2397 37979 2431
rect 38838 2428 38844 2440
rect 38799 2400 38844 2428
rect 37921 2391 37979 2397
rect 38838 2388 38844 2400
rect 38896 2388 38902 2440
rect 39758 2388 39764 2440
rect 39816 2428 39822 2440
rect 39853 2431 39911 2437
rect 39853 2428 39865 2431
rect 39816 2400 39865 2428
rect 39816 2388 39822 2400
rect 39853 2397 39865 2400
rect 39899 2397 39911 2431
rect 40954 2428 40960 2440
rect 40915 2400 40960 2428
rect 39853 2391 39911 2397
rect 40954 2388 40960 2400
rect 41012 2388 41018 2440
rect 41417 2431 41475 2437
rect 41417 2397 41429 2431
rect 41463 2428 41475 2431
rect 41506 2428 41512 2440
rect 41463 2400 41512 2428
rect 41463 2397 41475 2400
rect 41417 2391 41475 2397
rect 41506 2388 41512 2400
rect 41564 2388 41570 2440
rect 42426 2428 42432 2440
rect 42387 2400 42432 2428
rect 42426 2388 42432 2400
rect 42484 2388 42490 2440
rect 43441 2431 43499 2437
rect 43441 2397 43453 2431
rect 43487 2428 43499 2431
rect 43622 2428 43628 2440
rect 43487 2400 43628 2428
rect 43487 2397 43499 2400
rect 43441 2391 43499 2397
rect 43622 2388 43628 2400
rect 43680 2388 43686 2440
rect 44085 2431 44143 2437
rect 44085 2397 44097 2431
rect 44131 2428 44143 2431
rect 44266 2428 44272 2440
rect 44131 2400 44272 2428
rect 44131 2397 44143 2400
rect 44085 2391 44143 2397
rect 44266 2388 44272 2400
rect 44324 2388 44330 2440
rect 44818 2388 44824 2440
rect 44876 2428 44882 2440
rect 46768 2437 46796 2468
rect 45005 2431 45063 2437
rect 45005 2428 45017 2431
rect 44876 2400 45017 2428
rect 44876 2388 44882 2400
rect 45005 2397 45017 2400
rect 45051 2397 45063 2431
rect 46017 2431 46075 2437
rect 46017 2428 46029 2431
rect 45005 2391 45063 2397
rect 45526 2400 46029 2428
rect 17460 2332 28580 2360
rect 17460 2320 17466 2332
rect 29178 2320 29184 2372
rect 29236 2360 29242 2372
rect 30009 2363 30067 2369
rect 30009 2360 30021 2363
rect 29236 2332 30021 2360
rect 29236 2320 29242 2332
rect 30009 2329 30021 2332
rect 30055 2329 30067 2363
rect 30009 2323 30067 2329
rect 14182 2292 14188 2304
rect 12124 2264 13584 2292
rect 14143 2264 14188 2292
rect 12124 2252 12130 2264
rect 14182 2252 14188 2264
rect 14240 2252 14246 2304
rect 17770 2252 17776 2304
rect 17828 2292 17834 2304
rect 29196 2292 29224 2320
rect 17828 2264 29224 2292
rect 30101 2295 30159 2301
rect 17828 2252 17834 2264
rect 30101 2261 30113 2295
rect 30147 2292 30159 2295
rect 45526 2292 45554 2400
rect 46017 2397 46029 2400
rect 46063 2397 46075 2431
rect 46017 2391 46075 2397
rect 46753 2431 46811 2437
rect 46753 2397 46765 2431
rect 46799 2397 46811 2431
rect 46753 2391 46811 2397
rect 47118 2388 47124 2440
rect 47176 2428 47182 2440
rect 47857 2431 47915 2437
rect 47857 2428 47869 2431
rect 47176 2400 47869 2428
rect 47176 2388 47182 2400
rect 47857 2397 47869 2400
rect 47903 2397 47915 2431
rect 47857 2391 47915 2397
rect 49694 2360 49700 2372
rect 46216 2332 49700 2360
rect 46216 2301 46244 2332
rect 49694 2320 49700 2332
rect 49752 2320 49758 2372
rect 30147 2264 45554 2292
rect 46201 2295 46259 2301
rect 30147 2261 30159 2264
rect 30101 2255 30159 2261
rect 46201 2261 46213 2295
rect 46247 2261 46259 2295
rect 46201 2255 46259 2261
rect 48041 2295 48099 2301
rect 48041 2261 48053 2295
rect 48087 2292 48099 2295
rect 49234 2292 49240 2304
rect 48087 2264 49240 2292
rect 48087 2261 48099 2264
rect 48041 2255 48099 2261
rect 49234 2252 49240 2264
rect 49292 2252 49298 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 14 2048 20 2100
rect 72 2088 78 2100
rect 27890 2088 27896 2100
rect 72 2060 27896 2088
rect 72 2048 78 2060
rect 27890 2048 27896 2060
rect 27948 2048 27954 2100
rect 5902 1980 5908 2032
rect 5960 2020 5966 2032
rect 9398 2020 9404 2032
rect 5960 1992 9404 2020
rect 5960 1980 5966 1992
rect 9398 1980 9404 1992
rect 9456 1980 9462 2032
rect 10042 1980 10048 2032
rect 10100 2020 10106 2032
rect 13906 2020 13912 2032
rect 10100 1992 13912 2020
rect 10100 1980 10106 1992
rect 13906 1980 13912 1992
rect 13964 1980 13970 2032
rect 7558 1912 7564 1964
rect 7616 1952 7622 1964
rect 8294 1952 8300 1964
rect 7616 1924 8300 1952
rect 7616 1912 7622 1924
rect 8294 1912 8300 1924
rect 8352 1912 8358 1964
rect 8386 1912 8392 1964
rect 8444 1952 8450 1964
rect 14182 1952 14188 1964
rect 8444 1924 14188 1952
rect 8444 1912 8450 1924
rect 14182 1912 14188 1924
rect 14240 1912 14246 1964
rect 8849 1887 8907 1893
rect 8849 1853 8861 1887
rect 8895 1884 8907 1887
rect 12342 1884 12348 1896
rect 8895 1856 12348 1884
rect 8895 1853 8907 1856
rect 8849 1847 8907 1853
rect 12342 1844 12348 1856
rect 12400 1844 12406 1896
rect 12710 1844 12716 1896
rect 12768 1884 12774 1896
rect 17402 1884 17408 1896
rect 12768 1856 17408 1884
rect 12768 1844 12774 1856
rect 17402 1844 17408 1856
rect 17460 1844 17466 1896
rect 3142 1776 3148 1828
rect 3200 1816 3206 1828
rect 3602 1816 3608 1828
rect 3200 1788 3608 1816
rect 3200 1776 3206 1788
rect 3602 1776 3608 1788
rect 3660 1776 3666 1828
rect 6914 1776 6920 1828
rect 6972 1816 6978 1828
rect 13538 1816 13544 1828
rect 6972 1788 13544 1816
rect 6972 1776 6978 1788
rect 13538 1776 13544 1788
rect 13596 1776 13602 1828
rect 4706 1708 4712 1760
rect 4764 1748 4770 1760
rect 5626 1748 5632 1760
rect 4764 1720 5632 1748
rect 4764 1708 4770 1720
rect 5626 1708 5632 1720
rect 5684 1708 5690 1760
rect 7098 1708 7104 1760
rect 7156 1748 7162 1760
rect 15102 1748 15108 1760
rect 7156 1720 15108 1748
rect 7156 1708 7162 1720
rect 15102 1708 15108 1720
rect 15160 1708 15166 1760
rect 3602 1640 3608 1692
rect 3660 1680 3666 1692
rect 3878 1680 3884 1692
rect 3660 1652 3884 1680
rect 3660 1640 3666 1652
rect 3878 1640 3884 1652
rect 3936 1640 3942 1692
rect 7377 1683 7435 1689
rect 7377 1649 7389 1683
rect 7423 1680 7435 1683
rect 7423 1652 9628 1680
rect 7423 1649 7435 1652
rect 7377 1643 7435 1649
rect 7282 1572 7288 1624
rect 7340 1612 7346 1624
rect 8018 1612 8024 1624
rect 7340 1584 8024 1612
rect 7340 1572 7346 1584
rect 8018 1572 8024 1584
rect 8076 1572 8082 1624
rect 8294 1572 8300 1624
rect 8352 1612 8358 1624
rect 9490 1612 9496 1624
rect 8352 1584 9496 1612
rect 8352 1572 8358 1584
rect 9490 1572 9496 1584
rect 9548 1572 9554 1624
rect 9600 1612 9628 1652
rect 9674 1640 9680 1692
rect 9732 1680 9738 1692
rect 20162 1680 20168 1692
rect 9732 1652 20168 1680
rect 9732 1640 9738 1652
rect 20162 1640 20168 1652
rect 20220 1640 20226 1692
rect 11974 1612 11980 1624
rect 9600 1584 11980 1612
rect 11974 1572 11980 1584
rect 12032 1572 12038 1624
rect 13354 1572 13360 1624
rect 13412 1612 13418 1624
rect 15010 1612 15016 1624
rect 13412 1584 15016 1612
rect 13412 1572 13418 1584
rect 15010 1572 15016 1584
rect 15068 1572 15074 1624
rect 4522 1504 4528 1556
rect 4580 1544 4586 1556
rect 13262 1544 13268 1556
rect 4580 1516 13268 1544
rect 4580 1504 4586 1516
rect 13262 1504 13268 1516
rect 13320 1504 13326 1556
rect 7374 1476 7380 1488
rect 6886 1448 7380 1476
rect 4522 1300 4528 1352
rect 4580 1340 4586 1352
rect 5166 1340 5172 1352
rect 4580 1312 5172 1340
rect 4580 1300 4586 1312
rect 5166 1300 5172 1312
rect 5224 1300 5230 1352
rect 6886 1340 6914 1448
rect 7374 1436 7380 1448
rect 7432 1436 7438 1488
rect 9214 1436 9220 1488
rect 9272 1476 9278 1488
rect 18598 1476 18604 1488
rect 9272 1448 18604 1476
rect 9272 1436 9278 1448
rect 18598 1436 18604 1448
rect 18656 1436 18662 1488
rect 7006 1368 7012 1420
rect 7064 1408 7070 1420
rect 7742 1408 7748 1420
rect 7064 1380 7748 1408
rect 7064 1368 7070 1380
rect 7742 1368 7748 1380
rect 7800 1368 7806 1420
rect 8386 1408 8392 1420
rect 8312 1380 8392 1408
rect 7374 1340 7380 1352
rect 5920 1312 6914 1340
rect 7335 1312 7380 1340
rect 5920 1216 5948 1312
rect 7374 1300 7380 1312
rect 7432 1300 7438 1352
rect 7742 1232 7748 1284
rect 7800 1272 7806 1284
rect 8312 1272 8340 1380
rect 8386 1368 8392 1380
rect 8444 1368 8450 1420
rect 9030 1368 9036 1420
rect 9088 1408 9094 1420
rect 9088 1380 9260 1408
rect 9088 1368 9094 1380
rect 9232 1352 9260 1380
rect 9306 1368 9312 1420
rect 9364 1408 9370 1420
rect 9490 1408 9496 1420
rect 9364 1380 9496 1408
rect 9364 1368 9370 1380
rect 9490 1368 9496 1380
rect 9548 1368 9554 1420
rect 10042 1368 10048 1420
rect 10100 1408 10106 1420
rect 10594 1408 10600 1420
rect 10100 1380 10600 1408
rect 10100 1368 10106 1380
rect 10594 1368 10600 1380
rect 10652 1368 10658 1420
rect 11330 1368 11336 1420
rect 11388 1408 11394 1420
rect 17310 1408 17316 1420
rect 11388 1380 17316 1408
rect 11388 1368 11394 1380
rect 17310 1368 17316 1380
rect 17368 1368 17374 1420
rect 9214 1300 9220 1352
rect 9272 1300 9278 1352
rect 9766 1300 9772 1352
rect 9824 1340 9830 1352
rect 12342 1340 12348 1352
rect 9824 1312 12348 1340
rect 9824 1300 9830 1312
rect 12342 1300 12348 1312
rect 12400 1300 12406 1352
rect 12434 1300 12440 1352
rect 12492 1340 12498 1352
rect 14642 1340 14648 1352
rect 12492 1312 14648 1340
rect 12492 1300 12498 1312
rect 14642 1300 14648 1312
rect 14700 1300 14706 1352
rect 44450 1300 44456 1352
rect 44508 1340 44514 1352
rect 46474 1340 46480 1352
rect 44508 1312 46480 1340
rect 44508 1300 44514 1312
rect 46474 1300 46480 1312
rect 46532 1300 46538 1352
rect 7800 1244 8340 1272
rect 7800 1232 7806 1244
rect 10134 1232 10140 1284
rect 10192 1272 10198 1284
rect 14734 1272 14740 1284
rect 10192 1244 14740 1272
rect 10192 1232 10198 1244
rect 14734 1232 14740 1244
rect 14792 1232 14798 1284
rect 4154 1164 4160 1216
rect 4212 1204 4218 1216
rect 4798 1204 4804 1216
rect 4212 1176 4804 1204
rect 4212 1164 4218 1176
rect 4798 1164 4804 1176
rect 4856 1164 4862 1216
rect 5902 1164 5908 1216
rect 5960 1164 5966 1216
rect 10318 1164 10324 1216
rect 10376 1204 10382 1216
rect 10778 1204 10784 1216
rect 10376 1176 10784 1204
rect 10376 1164 10382 1176
rect 10778 1164 10784 1176
rect 10836 1164 10842 1216
rect 8386 1096 8392 1148
rect 8444 1136 8450 1148
rect 11054 1136 11060 1148
rect 8444 1108 11060 1136
rect 8444 1096 8450 1108
rect 11054 1096 11060 1108
rect 11112 1096 11118 1148
rect 9674 1028 9680 1080
rect 9732 1068 9738 1080
rect 11698 1068 11704 1080
rect 9732 1040 11704 1068
rect 9732 1028 9738 1040
rect 11698 1028 11704 1040
rect 11756 1028 11762 1080
rect 12802 1028 12808 1080
rect 12860 1068 12866 1080
rect 14918 1068 14924 1080
rect 12860 1040 14924 1068
rect 12860 1028 12866 1040
rect 14918 1028 14924 1040
rect 14976 1028 14982 1080
rect 10686 960 10692 1012
rect 10744 1000 10750 1012
rect 12618 1000 12624 1012
rect 10744 972 12624 1000
rect 10744 960 10750 972
rect 12618 960 12624 972
rect 12676 960 12682 1012
rect 5258 892 5264 944
rect 5316 932 5322 944
rect 6914 932 6920 944
rect 5316 904 6920 932
rect 5316 892 5322 904
rect 6914 892 6920 904
rect 6972 892 6978 944
rect 8846 932 8852 944
rect 8807 904 8852 932
rect 8846 892 8852 904
rect 8904 892 8910 944
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 1492 47243 1544 47252
rect 1492 47209 1501 47243
rect 1501 47209 1535 47243
rect 1535 47209 1544 47243
rect 1492 47200 1544 47209
rect 1860 47200 1912 47252
rect 3056 47200 3108 47252
rect 4620 47243 4672 47252
rect 4620 47209 4629 47243
rect 4629 47209 4663 47243
rect 4663 47209 4672 47243
rect 4620 47200 4672 47209
rect 4712 47200 4764 47252
rect 5540 47200 5592 47252
rect 6920 47200 6972 47252
rect 8300 47243 8352 47252
rect 8300 47209 8309 47243
rect 8309 47209 8343 47243
rect 8343 47209 8352 47243
rect 8300 47200 8352 47209
rect 9312 47200 9364 47252
rect 10600 47200 10652 47252
rect 11796 47200 11848 47252
rect 13084 47200 13136 47252
rect 14280 47200 14332 47252
rect 15568 47200 15620 47252
rect 16856 47200 16908 47252
rect 18052 47200 18104 47252
rect 19340 47200 19392 47252
rect 20720 47200 20772 47252
rect 22100 47243 22152 47252
rect 22100 47209 22109 47243
rect 22109 47209 22143 47243
rect 22143 47209 22152 47243
rect 22100 47200 22152 47209
rect 23020 47200 23072 47252
rect 24308 47200 24360 47252
rect 25596 47200 25648 47252
rect 26792 47200 26844 47252
rect 28080 47200 28132 47252
rect 29276 47200 29328 47252
rect 30564 47200 30616 47252
rect 31760 47200 31812 47252
rect 33140 47200 33192 47252
rect 33508 47200 33560 47252
rect 34520 47200 34572 47252
rect 35532 47200 35584 47252
rect 38016 47200 38068 47252
rect 38660 47200 38712 47252
rect 39304 47200 39356 47252
rect 40500 47200 40552 47252
rect 41788 47200 41840 47252
rect 43076 47200 43128 47252
rect 44272 47200 44324 47252
rect 45652 47200 45704 47252
rect 41052 47132 41104 47184
rect 40224 47064 40276 47116
rect 46848 47132 46900 47184
rect 48412 47200 48464 47252
rect 49240 47132 49292 47184
rect 1676 47039 1728 47048
rect 1676 47005 1685 47039
rect 1685 47005 1719 47039
rect 1719 47005 1728 47039
rect 1676 46996 1728 47005
rect 1952 46996 2004 47048
rect 2872 47039 2924 47048
rect 2872 47005 2881 47039
rect 2881 47005 2915 47039
rect 2915 47005 2924 47039
rect 2872 46996 2924 47005
rect 3792 47039 3844 47048
rect 3792 47005 3801 47039
rect 3801 47005 3835 47039
rect 3835 47005 3844 47039
rect 3792 46996 3844 47005
rect 4804 47039 4856 47048
rect 4804 47005 4813 47039
rect 4813 47005 4847 47039
rect 4847 47005 4856 47039
rect 4804 46996 4856 47005
rect 5816 46996 5868 47048
rect 6368 47039 6420 47048
rect 6368 47005 6377 47039
rect 6377 47005 6411 47039
rect 6411 47005 6420 47039
rect 6368 46996 6420 47005
rect 7380 47039 7432 47048
rect 7380 47005 7389 47039
rect 7389 47005 7423 47039
rect 7423 47005 7432 47039
rect 7380 46996 7432 47005
rect 8024 46996 8076 47048
rect 9772 46996 9824 47048
rect 10600 46996 10652 47048
rect 12900 46996 12952 47048
rect 13084 46996 13136 47048
rect 14372 47039 14424 47048
rect 14372 47005 14381 47039
rect 14381 47005 14415 47039
rect 14415 47005 14424 47039
rect 14372 46996 14424 47005
rect 15660 47039 15712 47048
rect 15660 47005 15669 47039
rect 15669 47005 15703 47039
rect 15703 47005 15712 47039
rect 15660 46996 15712 47005
rect 17776 46996 17828 47048
rect 18420 47039 18472 47048
rect 18420 47005 18429 47039
rect 18429 47005 18463 47039
rect 18463 47005 18472 47039
rect 18420 46996 18472 47005
rect 20444 46996 20496 47048
rect 20628 47039 20680 47048
rect 20628 47005 20637 47039
rect 20637 47005 20671 47039
rect 20671 47005 20680 47039
rect 20628 46996 20680 47005
rect 21916 47039 21968 47048
rect 21916 47005 21925 47039
rect 21925 47005 21959 47039
rect 21959 47005 21968 47039
rect 21916 46996 21968 47005
rect 23112 47039 23164 47048
rect 23112 47005 23121 47039
rect 23121 47005 23155 47039
rect 23155 47005 23164 47039
rect 23112 46996 23164 47005
rect 24400 47039 24452 47048
rect 24400 47005 24409 47039
rect 24409 47005 24443 47039
rect 24443 47005 24452 47039
rect 24400 46996 24452 47005
rect 25688 47039 25740 47048
rect 25688 47005 25697 47039
rect 25697 47005 25731 47039
rect 25731 47005 25740 47039
rect 25688 46996 25740 47005
rect 26976 47039 27028 47048
rect 26976 47005 26985 47039
rect 26985 47005 27019 47039
rect 27019 47005 27028 47039
rect 26976 46996 27028 47005
rect 28172 47039 28224 47048
rect 28172 47005 28181 47039
rect 28181 47005 28215 47039
rect 28215 47005 28224 47039
rect 28172 46996 28224 47005
rect 29552 47039 29604 47048
rect 29552 47005 29561 47039
rect 29561 47005 29595 47039
rect 29595 47005 29604 47039
rect 29552 46996 29604 47005
rect 30656 47039 30708 47048
rect 30656 47005 30665 47039
rect 30665 47005 30699 47039
rect 30699 47005 30708 47039
rect 30656 46996 30708 47005
rect 32404 47039 32456 47048
rect 32404 47005 32413 47039
rect 32413 47005 32447 47039
rect 32447 47005 32456 47039
rect 32404 46996 32456 47005
rect 33416 47039 33468 47048
rect 33416 47005 33425 47039
rect 33425 47005 33459 47039
rect 33459 47005 33468 47039
rect 33416 46996 33468 47005
rect 34704 47039 34756 47048
rect 8944 46928 8996 46980
rect 15200 46971 15252 46980
rect 15200 46937 15209 46971
rect 15209 46937 15243 46971
rect 15243 46937 15252 46971
rect 15200 46928 15252 46937
rect 33140 46928 33192 46980
rect 34704 47005 34713 47039
rect 34713 47005 34747 47039
rect 34747 47005 34756 47039
rect 34704 46996 34756 47005
rect 35624 47039 35676 47048
rect 35624 47005 35633 47039
rect 35633 47005 35667 47039
rect 35667 47005 35676 47039
rect 35624 46996 35676 47005
rect 37556 47039 37608 47048
rect 34612 46928 34664 46980
rect 37556 47005 37565 47039
rect 37565 47005 37599 47039
rect 37599 47005 37608 47039
rect 37556 46996 37608 47005
rect 38660 46996 38712 47048
rect 38752 46996 38804 47048
rect 39856 47039 39908 47048
rect 39856 47005 39865 47039
rect 39865 47005 39899 47039
rect 39899 47005 39908 47039
rect 39856 46996 39908 47005
rect 41144 46996 41196 47048
rect 41328 47039 41380 47048
rect 41328 47005 41337 47039
rect 41337 47005 41371 47039
rect 41371 47005 41380 47039
rect 41328 46996 41380 47005
rect 41880 46996 41932 47048
rect 43168 47039 43220 47048
rect 43168 47005 43177 47039
rect 43177 47005 43211 47039
rect 43211 47005 43220 47039
rect 43168 46996 43220 47005
rect 44180 47039 44232 47048
rect 44180 47005 44189 47039
rect 44189 47005 44223 47039
rect 44223 47005 44232 47039
rect 44180 46996 44232 47005
rect 42708 46928 42760 46980
rect 45744 46928 45796 46980
rect 47952 46996 48004 47048
rect 1032 46860 1084 46912
rect 28816 46860 28868 46912
rect 31300 46860 31352 46912
rect 34796 46860 34848 46912
rect 36820 46860 36872 46912
rect 40960 46860 41012 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 572 46656 624 46708
rect 2228 46656 2280 46708
rect 3516 46656 3568 46708
rect 4804 46656 4856 46708
rect 6368 46656 6420 46708
rect 7196 46656 7248 46708
rect 8484 46656 8536 46708
rect 9864 46656 9916 46708
rect 10968 46656 11020 46708
rect 12348 46656 12400 46708
rect 13452 46656 13504 46708
rect 14740 46656 14792 46708
rect 15936 46699 15988 46708
rect 15936 46665 15945 46699
rect 15945 46665 15979 46699
rect 15979 46665 15988 46699
rect 15936 46656 15988 46665
rect 17224 46656 17276 46708
rect 18512 46656 18564 46708
rect 19984 46699 20036 46708
rect 19984 46665 19993 46699
rect 19993 46665 20027 46699
rect 20027 46665 20036 46699
rect 19984 46656 20036 46665
rect 20444 46656 20496 46708
rect 20996 46656 21048 46708
rect 22192 46656 22244 46708
rect 23480 46656 23532 46708
rect 24676 46656 24728 46708
rect 25964 46656 26016 46708
rect 27252 46656 27304 46708
rect 29736 46656 29788 46708
rect 32404 46656 32456 46708
rect 33416 46656 33468 46708
rect 34704 46656 34756 46708
rect 35992 46656 36044 46708
rect 37188 46656 37240 46708
rect 37556 46656 37608 46708
rect 38660 46699 38712 46708
rect 38660 46665 38669 46699
rect 38669 46665 38703 46699
rect 38703 46665 38712 46699
rect 38660 46656 38712 46665
rect 39672 46656 39724 46708
rect 42248 46656 42300 46708
rect 43444 46656 43496 46708
rect 44732 46699 44784 46708
rect 44732 46665 44741 46699
rect 44741 46665 44775 46699
rect 44775 46665 44784 46699
rect 44732 46656 44784 46665
rect 46204 46699 46256 46708
rect 32036 46588 32088 46640
rect 41052 46588 41104 46640
rect 41144 46588 41196 46640
rect 46204 46665 46213 46699
rect 46213 46665 46247 46699
rect 46247 46665 46256 46699
rect 46204 46656 46256 46665
rect 48872 46656 48924 46708
rect 48044 46588 48096 46640
rect 2504 46520 2556 46572
rect 2596 46563 2648 46572
rect 2596 46529 2605 46563
rect 2605 46529 2639 46563
rect 2639 46529 2648 46563
rect 2596 46520 2648 46529
rect 3056 46520 3108 46572
rect 4160 46563 4212 46572
rect 4160 46529 4169 46563
rect 4169 46529 4203 46563
rect 4203 46529 4212 46563
rect 4160 46520 4212 46529
rect 6368 46563 6420 46572
rect 6368 46529 6377 46563
rect 6377 46529 6411 46563
rect 6411 46529 6420 46563
rect 6368 46520 6420 46529
rect 7748 46520 7800 46572
rect 8116 46520 8168 46572
rect 9864 46520 9916 46572
rect 11704 46520 11756 46572
rect 12808 46563 12860 46572
rect 12808 46529 12817 46563
rect 12817 46529 12851 46563
rect 12851 46529 12860 46563
rect 12808 46520 12860 46529
rect 13820 46563 13872 46572
rect 13820 46529 13829 46563
rect 13829 46529 13863 46563
rect 13863 46529 13872 46563
rect 13820 46520 13872 46529
rect 15108 46563 15160 46572
rect 15108 46529 15117 46563
rect 15117 46529 15151 46563
rect 15151 46529 15160 46563
rect 15108 46520 15160 46529
rect 15936 46520 15988 46572
rect 16672 46520 16724 46572
rect 17960 46563 18012 46572
rect 17960 46529 17969 46563
rect 17969 46529 18003 46563
rect 18003 46529 18012 46563
rect 17960 46520 18012 46529
rect 18696 46563 18748 46572
rect 18696 46529 18705 46563
rect 18705 46529 18739 46563
rect 18739 46529 18748 46563
rect 18696 46520 18748 46529
rect 19984 46520 20036 46572
rect 20720 46563 20772 46572
rect 20720 46529 20729 46563
rect 20729 46529 20763 46563
rect 20763 46529 20772 46563
rect 20720 46520 20772 46529
rect 21088 46520 21140 46572
rect 22560 46563 22612 46572
rect 22560 46529 22569 46563
rect 22569 46529 22603 46563
rect 22603 46529 22612 46563
rect 22560 46520 22612 46529
rect 23020 46520 23072 46572
rect 23756 46520 23808 46572
rect 24952 46520 25004 46572
rect 26240 46520 26292 46572
rect 27436 46563 27488 46572
rect 27436 46529 27445 46563
rect 27445 46529 27479 46563
rect 27479 46529 27488 46563
rect 27436 46520 27488 46529
rect 27528 46520 27580 46572
rect 28816 46520 28868 46572
rect 29828 46563 29880 46572
rect 29828 46529 29837 46563
rect 29837 46529 29871 46563
rect 29871 46529 29880 46563
rect 29828 46520 29880 46529
rect 31300 46520 31352 46572
rect 31760 46520 31812 46572
rect 34336 46563 34388 46572
rect 34336 46529 34345 46563
rect 34345 46529 34379 46563
rect 34379 46529 34388 46563
rect 34336 46520 34388 46529
rect 34796 46520 34848 46572
rect 36268 46520 36320 46572
rect 37372 46520 37424 46572
rect 39120 46520 39172 46572
rect 39764 46563 39816 46572
rect 39764 46529 39773 46563
rect 39773 46529 39807 46563
rect 39807 46529 39816 46563
rect 39764 46520 39816 46529
rect 40500 46563 40552 46572
rect 40500 46529 40509 46563
rect 40509 46529 40543 46563
rect 40543 46529 40552 46563
rect 40500 46520 40552 46529
rect 6000 46384 6052 46436
rect 3608 46359 3660 46368
rect 3608 46325 3617 46359
rect 3617 46325 3651 46359
rect 3651 46325 3660 46359
rect 3608 46316 3660 46325
rect 9404 46359 9456 46368
rect 9404 46325 9413 46359
rect 9413 46325 9447 46359
rect 9447 46325 9456 46359
rect 9404 46316 9456 46325
rect 11244 46316 11296 46368
rect 40132 46452 40184 46504
rect 32220 46384 32272 46436
rect 41052 46384 41104 46436
rect 41236 46520 41288 46572
rect 41788 46563 41840 46572
rect 41788 46529 41797 46563
rect 41797 46529 41831 46563
rect 41831 46529 41840 46563
rect 41788 46520 41840 46529
rect 42432 46563 42484 46572
rect 42432 46529 42441 46563
rect 42441 46529 42475 46563
rect 42475 46529 42484 46563
rect 42432 46520 42484 46529
rect 43536 46563 43588 46572
rect 43536 46529 43545 46563
rect 43545 46529 43579 46563
rect 43579 46529 43588 46563
rect 43536 46520 43588 46529
rect 44548 46563 44600 46572
rect 44548 46529 44557 46563
rect 44557 46529 44591 46563
rect 44591 46529 44600 46563
rect 44548 46520 44600 46529
rect 45284 46563 45336 46572
rect 45284 46529 45293 46563
rect 45293 46529 45327 46563
rect 45327 46529 45336 46563
rect 45284 46520 45336 46529
rect 46020 46563 46072 46572
rect 46020 46529 46029 46563
rect 46029 46529 46063 46563
rect 46063 46529 46072 46563
rect 46020 46520 46072 46529
rect 47860 46563 47912 46572
rect 14188 46316 14240 46368
rect 16672 46359 16724 46368
rect 16672 46325 16681 46359
rect 16681 46325 16715 46359
rect 16715 46325 16724 46359
rect 16672 46316 16724 46325
rect 24768 46316 24820 46368
rect 29000 46359 29052 46368
rect 29000 46325 29009 46359
rect 29009 46325 29043 46359
rect 29043 46325 29052 46359
rect 29000 46316 29052 46325
rect 40040 46316 40092 46368
rect 42708 46316 42760 46368
rect 45100 46316 45152 46368
rect 46204 46316 46256 46368
rect 47860 46529 47869 46563
rect 47869 46529 47903 46563
rect 47903 46529 47912 46563
rect 47860 46520 47912 46529
rect 48044 46427 48096 46436
rect 48044 46393 48053 46427
rect 48053 46393 48087 46427
rect 48087 46393 48096 46427
rect 48044 46384 48096 46393
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 1676 46112 1728 46164
rect 2504 46112 2556 46164
rect 3792 46155 3844 46164
rect 3792 46121 3801 46155
rect 3801 46121 3835 46155
rect 3835 46121 3844 46155
rect 3792 46112 3844 46121
rect 7380 46112 7432 46164
rect 12808 46112 12860 46164
rect 12900 46155 12952 46164
rect 12900 46121 12909 46155
rect 12909 46121 12943 46155
rect 12943 46121 12952 46155
rect 17776 46155 17828 46164
rect 12900 46112 12952 46121
rect 17776 46121 17785 46155
rect 17785 46121 17819 46155
rect 17819 46121 17828 46155
rect 17776 46112 17828 46121
rect 18420 46155 18472 46164
rect 18420 46121 18429 46155
rect 18429 46121 18463 46155
rect 18463 46121 18472 46155
rect 18420 46112 18472 46121
rect 20628 46112 20680 46164
rect 21916 46112 21968 46164
rect 26976 46112 27028 46164
rect 28172 46112 28224 46164
rect 28448 46112 28500 46164
rect 29552 46155 29604 46164
rect 29552 46121 29561 46155
rect 29561 46121 29595 46155
rect 29595 46121 29604 46155
rect 29552 46112 29604 46121
rect 30656 46112 30708 46164
rect 30932 46112 30984 46164
rect 32036 46112 32088 46164
rect 35440 46112 35492 46164
rect 35624 46112 35676 46164
rect 3056 45976 3108 46028
rect 8944 46019 8996 46028
rect 2044 45908 2096 45960
rect 2780 45951 2832 45960
rect 2780 45917 2789 45951
rect 2789 45917 2823 45951
rect 2823 45917 2832 45951
rect 2780 45908 2832 45917
rect 6920 45908 6972 45960
rect 8944 45985 8953 46019
rect 8953 45985 8987 46019
rect 8987 45985 8996 46019
rect 8944 45976 8996 45985
rect 29000 46044 29052 46096
rect 31852 46044 31904 46096
rect 8392 45951 8444 45960
rect 8392 45917 8401 45951
rect 8401 45917 8435 45951
rect 8435 45917 8444 45951
rect 8392 45908 8444 45917
rect 11152 45908 11204 45960
rect 5264 45840 5316 45892
rect 6460 45840 6512 45892
rect 9312 45840 9364 45892
rect 9404 45840 9456 45892
rect 11520 45840 11572 45892
rect 12900 45840 12952 45892
rect 15200 45908 15252 45960
rect 15844 45908 15896 45960
rect 17408 45908 17460 45960
rect 20720 45908 20772 45960
rect 21548 45951 21600 45960
rect 21548 45917 21557 45951
rect 21557 45917 21591 45951
rect 21591 45917 21600 45951
rect 21548 45908 21600 45917
rect 24860 45951 24912 45960
rect 24860 45917 24869 45951
rect 24869 45917 24903 45951
rect 24903 45917 24912 45951
rect 24860 45908 24912 45917
rect 26976 45908 27028 45960
rect 29736 45951 29788 45960
rect 14188 45840 14240 45892
rect 4988 45772 5040 45824
rect 5816 45815 5868 45824
rect 5816 45781 5825 45815
rect 5825 45781 5859 45815
rect 5859 45781 5868 45815
rect 5816 45772 5868 45781
rect 7748 45815 7800 45824
rect 7748 45781 7757 45815
rect 7757 45781 7791 45815
rect 7791 45781 7800 45815
rect 7748 45772 7800 45781
rect 9864 45772 9916 45824
rect 14280 45772 14332 45824
rect 16580 45840 16632 45892
rect 19432 45840 19484 45892
rect 22744 45840 22796 45892
rect 25136 45883 25188 45892
rect 25136 45849 25170 45883
rect 25170 45849 25188 45883
rect 25136 45840 25188 45849
rect 26424 45840 26476 45892
rect 29736 45917 29745 45951
rect 29745 45917 29779 45951
rect 29779 45917 29788 45951
rect 29736 45908 29788 45917
rect 30472 45908 30524 45960
rect 31392 45840 31444 45892
rect 14740 45772 14792 45824
rect 15108 45772 15160 45824
rect 15936 45815 15988 45824
rect 15936 45781 15945 45815
rect 15945 45781 15979 45815
rect 15979 45781 15988 45815
rect 15936 45772 15988 45781
rect 23756 45815 23808 45824
rect 23756 45781 23765 45815
rect 23765 45781 23799 45815
rect 23799 45781 23808 45815
rect 23756 45772 23808 45781
rect 26240 45815 26292 45824
rect 26240 45781 26249 45815
rect 26249 45781 26283 45815
rect 26283 45781 26292 45815
rect 26240 45772 26292 45781
rect 29736 45772 29788 45824
rect 33232 45908 33284 45960
rect 33324 45908 33376 45960
rect 34336 45908 34388 45960
rect 39120 46112 39172 46164
rect 39856 46112 39908 46164
rect 41328 46112 41380 46164
rect 41880 46155 41932 46164
rect 41880 46121 41889 46155
rect 41889 46121 41923 46155
rect 41923 46121 41932 46155
rect 41880 46112 41932 46121
rect 43168 46112 43220 46164
rect 44180 46112 44232 46164
rect 45560 46112 45612 46164
rect 46480 46112 46532 46164
rect 47308 46155 47360 46164
rect 47308 46121 47317 46155
rect 47317 46121 47351 46155
rect 47351 46121 47360 46155
rect 47308 46112 47360 46121
rect 35992 45951 36044 45960
rect 35992 45917 36001 45951
rect 36001 45917 36035 45951
rect 36035 45917 36044 45951
rect 35992 45908 36044 45917
rect 39948 46044 40000 46096
rect 40132 46044 40184 46096
rect 45100 46044 45152 46096
rect 46756 46044 46808 46096
rect 31944 45840 31996 45892
rect 39120 45951 39172 45960
rect 39120 45917 39129 45951
rect 39129 45917 39163 45951
rect 39163 45917 39172 45951
rect 39120 45908 39172 45917
rect 39672 45908 39724 45960
rect 41512 45908 41564 45960
rect 41696 45951 41748 45960
rect 41696 45917 41705 45951
rect 41705 45917 41739 45951
rect 41739 45917 41748 45951
rect 41696 45908 41748 45917
rect 43904 45908 43956 45960
rect 46480 45908 46532 45960
rect 47860 45951 47912 45960
rect 47860 45917 47869 45951
rect 47869 45917 47903 45951
rect 47903 45917 47912 45951
rect 47860 45908 47912 45917
rect 36452 45840 36504 45892
rect 33140 45772 33192 45824
rect 34796 45815 34848 45824
rect 34796 45781 34805 45815
rect 34805 45781 34839 45815
rect 34839 45781 34848 45815
rect 34796 45772 34848 45781
rect 35440 45772 35492 45824
rect 44732 45840 44784 45892
rect 45284 45840 45336 45892
rect 37372 45815 37424 45824
rect 37372 45781 37381 45815
rect 37381 45781 37415 45815
rect 37415 45781 37424 45815
rect 37372 45772 37424 45781
rect 48044 45815 48096 45824
rect 48044 45781 48053 45815
rect 48053 45781 48087 45815
rect 48087 45781 48096 45815
rect 48044 45772 48096 45781
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 5264 45611 5316 45620
rect 5264 45577 5273 45611
rect 5273 45577 5307 45611
rect 5307 45577 5316 45611
rect 5264 45568 5316 45577
rect 6460 45611 6512 45620
rect 6460 45577 6469 45611
rect 6469 45577 6503 45611
rect 6503 45577 6512 45611
rect 6460 45568 6512 45577
rect 9312 45611 9364 45620
rect 2780 45500 2832 45552
rect 2504 45432 2556 45484
rect 4528 45475 4580 45484
rect 4528 45441 4537 45475
rect 4537 45441 4571 45475
rect 4571 45441 4580 45475
rect 4528 45432 4580 45441
rect 4712 45475 4764 45484
rect 4712 45441 4721 45475
rect 4721 45441 4755 45475
rect 4755 45441 4764 45475
rect 4712 45432 4764 45441
rect 5816 45432 5868 45484
rect 7748 45500 7800 45552
rect 9312 45577 9321 45611
rect 9321 45577 9355 45611
rect 9355 45577 9364 45611
rect 9312 45568 9364 45577
rect 11520 45611 11572 45620
rect 11520 45577 11529 45611
rect 11529 45577 11563 45611
rect 11563 45577 11572 45611
rect 11520 45568 11572 45577
rect 14280 45611 14332 45620
rect 14280 45577 14289 45611
rect 14289 45577 14323 45611
rect 14323 45577 14332 45611
rect 14280 45568 14332 45577
rect 22744 45611 22796 45620
rect 22744 45577 22753 45611
rect 22753 45577 22787 45611
rect 22787 45577 22796 45611
rect 22744 45568 22796 45577
rect 25136 45568 25188 45620
rect 28448 45568 28500 45620
rect 30472 45568 30524 45620
rect 31392 45568 31444 45620
rect 4620 45364 4672 45416
rect 4804 45407 4856 45416
rect 4804 45373 4813 45407
rect 4813 45373 4847 45407
rect 4847 45373 4856 45407
rect 4804 45364 4856 45373
rect 1952 45339 2004 45348
rect 1952 45305 1961 45339
rect 1961 45305 1995 45339
rect 1995 45305 2004 45339
rect 1952 45296 2004 45305
rect 4160 45296 4212 45348
rect 4988 45364 5040 45416
rect 6460 45364 6512 45416
rect 7196 45475 7248 45484
rect 7196 45441 7205 45475
rect 7205 45441 7239 45475
rect 7239 45441 7248 45475
rect 8392 45500 8444 45552
rect 10048 45500 10100 45552
rect 7196 45432 7248 45441
rect 6736 45296 6788 45348
rect 8300 45364 8352 45416
rect 8852 45475 8904 45484
rect 8852 45441 8861 45475
rect 8861 45441 8895 45475
rect 8895 45441 8904 45475
rect 8852 45432 8904 45441
rect 9864 45432 9916 45484
rect 10416 45475 10468 45484
rect 2688 45228 2740 45280
rect 7012 45296 7064 45348
rect 8024 45339 8076 45348
rect 8024 45305 8033 45339
rect 8033 45305 8067 45339
rect 8067 45305 8076 45339
rect 8024 45296 8076 45305
rect 9404 45364 9456 45416
rect 10416 45441 10425 45475
rect 10425 45441 10459 45475
rect 10459 45441 10468 45475
rect 10416 45432 10468 45441
rect 12808 45500 12860 45552
rect 11244 45364 11296 45416
rect 12900 45475 12952 45484
rect 9772 45339 9824 45348
rect 9772 45305 9781 45339
rect 9781 45305 9815 45339
rect 9815 45305 9824 45339
rect 9772 45296 9824 45305
rect 10600 45339 10652 45348
rect 10600 45305 10609 45339
rect 10609 45305 10643 45339
rect 10643 45305 10652 45339
rect 10600 45296 10652 45305
rect 11980 45407 12032 45416
rect 11980 45373 11989 45407
rect 11989 45373 12023 45407
rect 12023 45373 12032 45407
rect 11980 45364 12032 45373
rect 12164 45364 12216 45416
rect 12900 45441 12909 45475
rect 12909 45441 12943 45475
rect 12943 45441 12952 45475
rect 12900 45432 12952 45441
rect 13728 45475 13780 45484
rect 13728 45441 13737 45475
rect 13737 45441 13771 45475
rect 13771 45441 13780 45475
rect 13728 45432 13780 45441
rect 14740 45432 14792 45484
rect 16580 45500 16632 45552
rect 15016 45475 15068 45484
rect 15016 45441 15025 45475
rect 15025 45441 15059 45475
rect 15059 45441 15068 45475
rect 15016 45432 15068 45441
rect 15108 45407 15160 45416
rect 12440 45296 12492 45348
rect 13084 45339 13136 45348
rect 13084 45305 13093 45339
rect 13093 45305 13127 45339
rect 13127 45305 13136 45339
rect 13084 45296 13136 45305
rect 11980 45228 12032 45280
rect 12900 45228 12952 45280
rect 15108 45373 15117 45407
rect 15117 45373 15151 45407
rect 15151 45373 15160 45407
rect 15108 45364 15160 45373
rect 14464 45296 14516 45348
rect 15936 45432 15988 45484
rect 18604 45475 18656 45484
rect 18604 45441 18638 45475
rect 18638 45441 18656 45475
rect 18604 45432 18656 45441
rect 17408 45364 17460 45416
rect 18328 45407 18380 45416
rect 18328 45373 18337 45407
rect 18337 45373 18371 45407
rect 18371 45373 18380 45407
rect 18328 45364 18380 45373
rect 16212 45228 16264 45280
rect 17868 45228 17920 45280
rect 19432 45296 19484 45348
rect 20720 45296 20772 45348
rect 21548 45296 21600 45348
rect 19708 45271 19760 45280
rect 19708 45237 19717 45271
rect 19717 45237 19751 45271
rect 19751 45237 19760 45271
rect 19708 45228 19760 45237
rect 19984 45228 20036 45280
rect 23756 45500 23808 45552
rect 23940 45500 23992 45552
rect 23020 45432 23072 45484
rect 23848 45432 23900 45484
rect 26240 45500 26292 45552
rect 28540 45500 28592 45552
rect 23664 45364 23716 45416
rect 26332 45432 26384 45484
rect 28264 45432 28316 45484
rect 29000 45432 29052 45484
rect 31208 45500 31260 45552
rect 31944 45500 31996 45552
rect 32128 45568 32180 45620
rect 40224 45568 40276 45620
rect 33324 45500 33376 45552
rect 30932 45432 30984 45484
rect 33140 45432 33192 45484
rect 33232 45475 33284 45484
rect 33232 45441 33241 45475
rect 33241 45441 33275 45475
rect 33275 45441 33284 45475
rect 35992 45500 36044 45552
rect 36176 45500 36228 45552
rect 33232 45432 33284 45441
rect 33508 45475 33560 45484
rect 33508 45441 33542 45475
rect 33542 45441 33560 45475
rect 33508 45432 33560 45441
rect 35716 45432 35768 45484
rect 39120 45500 39172 45552
rect 41236 45568 41288 45620
rect 41696 45568 41748 45620
rect 42432 45611 42484 45620
rect 42432 45577 42441 45611
rect 42441 45577 42475 45611
rect 42475 45577 42484 45611
rect 42432 45568 42484 45577
rect 43536 45568 43588 45620
rect 43904 45611 43956 45620
rect 43904 45577 43913 45611
rect 43913 45577 43947 45611
rect 43947 45577 43956 45611
rect 43904 45568 43956 45577
rect 44548 45568 44600 45620
rect 49700 45568 49752 45620
rect 23756 45296 23808 45348
rect 27436 45364 27488 45416
rect 27988 45364 28040 45416
rect 31116 45407 31168 45416
rect 31116 45373 31125 45407
rect 31125 45373 31159 45407
rect 31159 45373 31168 45407
rect 31116 45364 31168 45373
rect 25688 45339 25740 45348
rect 25688 45305 25697 45339
rect 25697 45305 25731 45339
rect 25731 45305 25740 45339
rect 25688 45296 25740 45305
rect 30196 45339 30248 45348
rect 26332 45228 26384 45280
rect 26976 45228 27028 45280
rect 30196 45305 30205 45339
rect 30205 45305 30239 45339
rect 30239 45305 30248 45339
rect 35348 45364 35400 45416
rect 38660 45432 38712 45484
rect 36176 45407 36228 45416
rect 36176 45373 36185 45407
rect 36185 45373 36219 45407
rect 36219 45373 36228 45407
rect 36176 45364 36228 45373
rect 30196 45296 30248 45305
rect 33140 45296 33192 45348
rect 34612 45271 34664 45280
rect 34612 45237 34621 45271
rect 34621 45237 34655 45271
rect 34655 45237 34664 45271
rect 35348 45271 35400 45280
rect 34612 45228 34664 45237
rect 35348 45237 35357 45271
rect 35357 45237 35391 45271
rect 35391 45237 35400 45271
rect 35348 45228 35400 45237
rect 35992 45296 36044 45348
rect 40040 45364 40092 45416
rect 41512 45432 41564 45484
rect 44456 45475 44508 45484
rect 44456 45441 44465 45475
rect 44465 45441 44499 45475
rect 44499 45441 44508 45475
rect 44456 45432 44508 45441
rect 45100 45475 45152 45484
rect 45100 45441 45109 45475
rect 45109 45441 45143 45475
rect 45143 45441 45152 45475
rect 45100 45432 45152 45441
rect 46020 45475 46072 45484
rect 46020 45441 46029 45475
rect 46029 45441 46063 45475
rect 46063 45441 46072 45475
rect 46020 45432 46072 45441
rect 45652 45364 45704 45416
rect 45836 45296 45888 45348
rect 45928 45296 45980 45348
rect 38660 45271 38712 45280
rect 38660 45237 38669 45271
rect 38669 45237 38703 45271
rect 38703 45237 38712 45271
rect 38660 45228 38712 45237
rect 39672 45271 39724 45280
rect 39672 45237 39681 45271
rect 39681 45237 39715 45271
rect 39715 45237 39724 45271
rect 39672 45228 39724 45237
rect 46480 45228 46532 45280
rect 46848 45228 46900 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 2504 45067 2556 45076
rect 2504 45033 2513 45067
rect 2513 45033 2547 45067
rect 2547 45033 2556 45067
rect 2504 45024 2556 45033
rect 4620 45024 4672 45076
rect 5448 45024 5500 45076
rect 6920 45067 6972 45076
rect 6920 45033 6929 45067
rect 6929 45033 6963 45067
rect 6963 45033 6972 45067
rect 6920 45024 6972 45033
rect 8392 45024 8444 45076
rect 14372 45067 14424 45076
rect 14372 45033 14381 45067
rect 14381 45033 14415 45067
rect 14415 45033 14424 45067
rect 14372 45024 14424 45033
rect 15660 45067 15712 45076
rect 15660 45033 15669 45067
rect 15669 45033 15703 45067
rect 15703 45033 15712 45067
rect 15660 45024 15712 45033
rect 18328 45024 18380 45076
rect 4988 44999 5040 45008
rect 4988 44965 4997 44999
rect 4997 44965 5031 44999
rect 5031 44965 5040 44999
rect 4988 44956 5040 44965
rect 10416 44956 10468 45008
rect 4804 44888 4856 44940
rect 7012 44888 7064 44940
rect 2688 44863 2740 44872
rect 2688 44829 2697 44863
rect 2697 44829 2731 44863
rect 2731 44829 2740 44863
rect 2688 44820 2740 44829
rect 2044 44727 2096 44736
rect 2044 44693 2053 44727
rect 2053 44693 2087 44727
rect 2087 44693 2096 44727
rect 2044 44684 2096 44693
rect 2688 44684 2740 44736
rect 3056 44863 3108 44872
rect 3056 44829 3065 44863
rect 3065 44829 3099 44863
rect 3099 44829 3108 44863
rect 3056 44820 3108 44829
rect 3608 44820 3660 44872
rect 12532 44888 12584 44940
rect 13728 44956 13780 45008
rect 16672 44956 16724 45008
rect 17132 44956 17184 45008
rect 17316 44888 17368 44940
rect 17868 44888 17920 44940
rect 18604 44956 18656 45008
rect 18788 44956 18840 45008
rect 20720 45024 20772 45076
rect 22100 45024 22152 45076
rect 22560 45024 22612 45076
rect 23112 45024 23164 45076
rect 24584 45024 24636 45076
rect 26976 45067 27028 45076
rect 26976 45033 26985 45067
rect 26985 45033 27019 45067
rect 27019 45033 27028 45067
rect 26976 45024 27028 45033
rect 28264 45067 28316 45076
rect 28264 45033 28273 45067
rect 28273 45033 28307 45067
rect 28307 45033 28316 45067
rect 28264 45024 28316 45033
rect 28356 45024 28408 45076
rect 28816 45024 28868 45076
rect 4344 44752 4396 44804
rect 4712 44752 4764 44804
rect 5264 44752 5316 44804
rect 14188 44863 14240 44872
rect 14188 44829 14197 44863
rect 14197 44829 14231 44863
rect 14231 44829 14240 44863
rect 14188 44820 14240 44829
rect 14924 44820 14976 44872
rect 16212 44820 16264 44872
rect 18052 44820 18104 44872
rect 18328 44863 18380 44872
rect 18328 44829 18337 44863
rect 18337 44829 18371 44863
rect 18371 44829 18380 44863
rect 18328 44820 18380 44829
rect 19708 44820 19760 44872
rect 20352 44863 20404 44872
rect 20352 44829 20361 44863
rect 20361 44829 20395 44863
rect 20395 44829 20404 44863
rect 20352 44820 20404 44829
rect 21548 44888 21600 44940
rect 24768 44956 24820 45008
rect 28356 44888 28408 44940
rect 28540 44888 28592 44940
rect 33232 45024 33284 45076
rect 33508 45067 33560 45076
rect 33508 45033 33517 45067
rect 33517 45033 33551 45067
rect 33551 45033 33560 45067
rect 33508 45024 33560 45033
rect 34336 45024 34388 45076
rect 35348 45024 35400 45076
rect 36452 45067 36504 45076
rect 31760 44999 31812 45008
rect 31760 44965 31769 44999
rect 31769 44965 31803 44999
rect 31803 44965 31812 44999
rect 31760 44956 31812 44965
rect 3884 44727 3936 44736
rect 3884 44693 3893 44727
rect 3893 44693 3927 44727
rect 3927 44693 3936 44727
rect 3884 44684 3936 44693
rect 6460 44684 6512 44736
rect 8300 44727 8352 44736
rect 8300 44693 8309 44727
rect 8309 44693 8343 44727
rect 8343 44693 8352 44727
rect 8300 44684 8352 44693
rect 9680 44684 9732 44736
rect 10784 44727 10836 44736
rect 10784 44693 10793 44727
rect 10793 44693 10827 44727
rect 10827 44693 10836 44727
rect 10784 44684 10836 44693
rect 11244 44727 11296 44736
rect 11244 44693 11253 44727
rect 11253 44693 11287 44727
rect 11287 44693 11296 44727
rect 11244 44684 11296 44693
rect 13728 44684 13780 44736
rect 15016 44684 15068 44736
rect 16212 44727 16264 44736
rect 16212 44693 16221 44727
rect 16221 44693 16255 44727
rect 16255 44693 16264 44727
rect 16212 44684 16264 44693
rect 17316 44684 17368 44736
rect 19432 44752 19484 44804
rect 24584 44863 24636 44872
rect 24584 44829 24593 44863
rect 24593 44829 24627 44863
rect 24627 44829 24636 44863
rect 24584 44820 24636 44829
rect 28448 44863 28500 44872
rect 28448 44829 28457 44863
rect 28457 44829 28491 44863
rect 28491 44829 28500 44863
rect 28448 44820 28500 44829
rect 20904 44752 20956 44804
rect 23572 44752 23624 44804
rect 27344 44752 27396 44804
rect 20996 44684 21048 44736
rect 23940 44684 23992 44736
rect 24400 44727 24452 44736
rect 24400 44693 24409 44727
rect 24409 44693 24443 44727
rect 24443 44693 24452 44727
rect 24400 44684 24452 44693
rect 28540 44684 28592 44736
rect 28816 44863 28868 44872
rect 28816 44829 28825 44863
rect 28825 44829 28859 44863
rect 28859 44829 28868 44863
rect 29000 44863 29052 44872
rect 28816 44820 28868 44829
rect 29000 44829 29009 44863
rect 29009 44829 29043 44863
rect 29043 44829 29052 44863
rect 29000 44820 29052 44829
rect 28908 44752 28960 44804
rect 32220 44888 32272 44940
rect 34796 44956 34848 45008
rect 35900 44956 35952 45008
rect 36452 45033 36461 45067
rect 36461 45033 36495 45067
rect 36495 45033 36504 45067
rect 36452 45024 36504 45033
rect 39120 45024 39172 45076
rect 43904 45067 43956 45076
rect 43904 45033 43913 45067
rect 43913 45033 43947 45067
rect 43947 45033 43956 45067
rect 43904 45024 43956 45033
rect 45100 45067 45152 45076
rect 45100 45033 45109 45067
rect 45109 45033 45143 45067
rect 45143 45033 45152 45067
rect 45100 45024 45152 45033
rect 46020 45067 46072 45076
rect 46020 45033 46029 45067
rect 46029 45033 46063 45067
rect 46063 45033 46072 45067
rect 46020 45024 46072 45033
rect 47584 45024 47636 45076
rect 39672 44956 39724 45008
rect 33140 44931 33192 44940
rect 29736 44752 29788 44804
rect 30472 44752 30524 44804
rect 31208 44820 31260 44872
rect 33140 44897 33149 44931
rect 33149 44897 33183 44931
rect 33183 44897 33192 44931
rect 33140 44888 33192 44897
rect 36176 44888 36228 44940
rect 44456 44888 44508 44940
rect 33232 44820 33284 44872
rect 34612 44820 34664 44872
rect 35716 44863 35768 44872
rect 35716 44829 35725 44863
rect 35725 44829 35759 44863
rect 35759 44829 35768 44863
rect 35716 44820 35768 44829
rect 35808 44820 35860 44872
rect 36084 44863 36136 44872
rect 36084 44829 36093 44863
rect 36093 44829 36127 44863
rect 36127 44829 36136 44863
rect 36084 44820 36136 44829
rect 37372 44820 37424 44872
rect 45744 44820 45796 44872
rect 47308 44888 47360 44940
rect 47676 44863 47728 44872
rect 47676 44829 47685 44863
rect 47685 44829 47719 44863
rect 47719 44829 47728 44863
rect 47676 44820 47728 44829
rect 31024 44684 31076 44736
rect 32220 44727 32272 44736
rect 32220 44693 32229 44727
rect 32229 44693 32263 44727
rect 32263 44693 32272 44727
rect 32220 44684 32272 44693
rect 34704 44684 34756 44736
rect 35808 44684 35860 44736
rect 40500 44684 40552 44736
rect 44364 44727 44416 44736
rect 44364 44693 44373 44727
rect 44373 44693 44407 44727
rect 44407 44693 44416 44727
rect 44364 44684 44416 44693
rect 46848 44684 46900 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 8852 44480 8904 44532
rect 6736 44412 6788 44464
rect 9680 44412 9732 44464
rect 10784 44412 10836 44464
rect 2780 44276 2832 44328
rect 4344 44319 4396 44328
rect 4344 44285 4353 44319
rect 4353 44285 4387 44319
rect 4387 44285 4396 44319
rect 4344 44276 4396 44285
rect 4804 44276 4856 44328
rect 3056 44208 3108 44260
rect 2780 44140 2832 44192
rect 4988 44140 5040 44192
rect 6460 44140 6512 44192
rect 10232 44387 10284 44396
rect 10232 44353 10241 44387
rect 10241 44353 10275 44387
rect 10275 44353 10284 44387
rect 10232 44344 10284 44353
rect 11704 44387 11756 44396
rect 11704 44353 11713 44387
rect 11713 44353 11747 44387
rect 11747 44353 11756 44387
rect 11704 44344 11756 44353
rect 11980 44387 12032 44396
rect 11980 44353 11989 44387
rect 11989 44353 12023 44387
rect 12023 44353 12032 44387
rect 11980 44344 12032 44353
rect 12164 44344 12216 44396
rect 13176 44480 13228 44532
rect 14464 44523 14516 44532
rect 14464 44489 14473 44523
rect 14473 44489 14507 44523
rect 14507 44489 14516 44523
rect 14464 44480 14516 44489
rect 14924 44480 14976 44532
rect 15844 44523 15896 44532
rect 15844 44489 15853 44523
rect 15853 44489 15887 44523
rect 15887 44489 15896 44523
rect 15844 44480 15896 44489
rect 16212 44480 16264 44532
rect 18328 44480 18380 44532
rect 20536 44480 20588 44532
rect 20904 44523 20956 44532
rect 20904 44489 20913 44523
rect 20913 44489 20947 44523
rect 20947 44489 20956 44523
rect 20904 44480 20956 44489
rect 20996 44480 21048 44532
rect 45652 44480 45704 44532
rect 45836 44480 45888 44532
rect 47860 44480 47912 44532
rect 12624 44412 12676 44464
rect 19524 44387 19576 44396
rect 19524 44353 19533 44387
rect 19533 44353 19567 44387
rect 19567 44353 19576 44387
rect 19524 44344 19576 44353
rect 20168 44387 20220 44396
rect 20168 44353 20177 44387
rect 20177 44353 20211 44387
rect 20211 44353 20220 44387
rect 20168 44344 20220 44353
rect 20260 44344 20312 44396
rect 12440 44276 12492 44328
rect 13176 44276 13228 44328
rect 15936 44276 15988 44328
rect 19432 44276 19484 44328
rect 20536 44319 20588 44328
rect 20536 44285 20545 44319
rect 20545 44285 20579 44319
rect 20579 44285 20588 44319
rect 20536 44276 20588 44285
rect 22100 44344 22152 44396
rect 22284 44387 22336 44396
rect 22284 44353 22293 44387
rect 22293 44353 22327 44387
rect 22327 44353 22336 44387
rect 22284 44344 22336 44353
rect 23572 44387 23624 44396
rect 21272 44276 21324 44328
rect 22192 44276 22244 44328
rect 23572 44353 23581 44387
rect 23581 44353 23615 44387
rect 23615 44353 23624 44387
rect 23572 44344 23624 44353
rect 23756 44387 23808 44396
rect 23756 44353 23765 44387
rect 23765 44353 23799 44387
rect 23799 44353 23808 44387
rect 23756 44344 23808 44353
rect 24768 44344 24820 44396
rect 24860 44344 24912 44396
rect 25136 44344 25188 44396
rect 27344 44344 27396 44396
rect 28724 44412 28776 44464
rect 30472 44455 30524 44464
rect 30472 44421 30481 44455
rect 30481 44421 30515 44455
rect 30515 44421 30524 44455
rect 30472 44412 30524 44421
rect 29092 44344 29144 44396
rect 31760 44412 31812 44464
rect 34336 44412 34388 44464
rect 44732 44455 44784 44464
rect 44732 44421 44741 44455
rect 44741 44421 44775 44455
rect 44775 44421 44784 44455
rect 44732 44412 44784 44421
rect 30932 44387 30984 44396
rect 30932 44353 30941 44387
rect 30941 44353 30975 44387
rect 30975 44353 30984 44387
rect 30932 44344 30984 44353
rect 31208 44387 31260 44396
rect 31208 44353 31217 44387
rect 31217 44353 31251 44387
rect 31251 44353 31260 44387
rect 31208 44344 31260 44353
rect 31392 44344 31444 44396
rect 47676 44412 47728 44464
rect 45744 44344 45796 44396
rect 46940 44344 46992 44396
rect 23480 44276 23532 44328
rect 24676 44276 24728 44328
rect 28080 44276 28132 44328
rect 29000 44276 29052 44328
rect 30196 44276 30248 44328
rect 31116 44276 31168 44328
rect 31300 44276 31352 44328
rect 10784 44140 10836 44192
rect 11612 44140 11664 44192
rect 13268 44140 13320 44192
rect 17224 44140 17276 44192
rect 18788 44140 18840 44192
rect 19524 44140 19576 44192
rect 22008 44140 22060 44192
rect 23480 44140 23532 44192
rect 23664 44140 23716 44192
rect 23940 44140 23992 44192
rect 24584 44140 24636 44192
rect 30748 44208 30800 44260
rect 31208 44208 31260 44260
rect 44364 44208 44416 44260
rect 26424 44183 26476 44192
rect 26424 44149 26433 44183
rect 26433 44149 26467 44183
rect 26467 44149 26476 44183
rect 26424 44140 26476 44149
rect 28080 44140 28132 44192
rect 30104 44140 30156 44192
rect 35624 44140 35676 44192
rect 46940 44183 46992 44192
rect 46940 44149 46949 44183
rect 46949 44149 46983 44183
rect 46983 44149 46992 44183
rect 46940 44140 46992 44149
rect 48044 44183 48096 44192
rect 48044 44149 48053 44183
rect 48053 44149 48087 44183
rect 48087 44149 48096 44183
rect 48044 44140 48096 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 2872 43936 2924 43988
rect 5448 43936 5500 43988
rect 11152 43936 11204 43988
rect 3884 43911 3936 43920
rect 3884 43877 3893 43911
rect 3893 43877 3927 43911
rect 3927 43877 3936 43911
rect 3884 43868 3936 43877
rect 4620 43868 4672 43920
rect 7012 43868 7064 43920
rect 4988 43800 5040 43852
rect 2044 43732 2096 43784
rect 8208 43800 8260 43852
rect 2964 43707 3016 43716
rect 2964 43673 2982 43707
rect 2982 43673 3016 43707
rect 2964 43664 3016 43673
rect 3516 43664 3568 43716
rect 4804 43596 4856 43648
rect 46940 43936 46992 43988
rect 47216 43936 47268 43988
rect 47952 43936 48004 43988
rect 11980 43800 12032 43852
rect 35072 43868 35124 43920
rect 38660 43868 38712 43920
rect 39764 43868 39816 43920
rect 45652 43911 45704 43920
rect 45652 43877 45661 43911
rect 45661 43877 45695 43911
rect 45695 43877 45704 43911
rect 45652 43868 45704 43877
rect 46204 43911 46256 43920
rect 46204 43877 46213 43911
rect 46213 43877 46247 43911
rect 46247 43877 46256 43911
rect 46204 43868 46256 43877
rect 46664 43868 46716 43920
rect 11612 43775 11664 43784
rect 11612 43741 11630 43775
rect 11630 43741 11664 43775
rect 11612 43732 11664 43741
rect 12900 43800 12952 43852
rect 13176 43843 13228 43852
rect 13176 43809 13185 43843
rect 13185 43809 13219 43843
rect 13219 43809 13228 43843
rect 13176 43800 13228 43809
rect 15108 43800 15160 43852
rect 12164 43732 12216 43784
rect 13820 43732 13872 43784
rect 16672 43800 16724 43852
rect 16764 43732 16816 43784
rect 18328 43800 18380 43852
rect 18604 43800 18656 43852
rect 21180 43800 21232 43852
rect 21272 43800 21324 43852
rect 17132 43775 17184 43784
rect 17132 43741 17141 43775
rect 17141 43741 17175 43775
rect 17175 43741 17184 43775
rect 17132 43732 17184 43741
rect 17224 43775 17276 43784
rect 17224 43741 17233 43775
rect 17233 43741 17267 43775
rect 17267 43741 17276 43775
rect 17224 43732 17276 43741
rect 17408 43775 17460 43784
rect 17408 43741 17417 43775
rect 17417 43741 17451 43775
rect 17451 43741 17460 43775
rect 17408 43732 17460 43741
rect 18052 43732 18104 43784
rect 20168 43732 20220 43784
rect 20260 43732 20312 43784
rect 22192 43732 22244 43784
rect 22928 43732 22980 43784
rect 24768 43843 24820 43852
rect 24768 43809 24777 43843
rect 24777 43809 24811 43843
rect 24811 43809 24820 43843
rect 24768 43800 24820 43809
rect 25136 43843 25188 43852
rect 25136 43809 25145 43843
rect 25145 43809 25179 43843
rect 25179 43809 25188 43843
rect 25136 43800 25188 43809
rect 27344 43843 27396 43852
rect 27344 43809 27353 43843
rect 27353 43809 27387 43843
rect 27387 43809 27396 43843
rect 27344 43800 27396 43809
rect 23572 43775 23624 43784
rect 23572 43741 23581 43775
rect 23581 43741 23615 43775
rect 23615 43741 23624 43775
rect 23572 43732 23624 43741
rect 13268 43664 13320 43716
rect 15752 43707 15804 43716
rect 15752 43673 15761 43707
rect 15761 43673 15795 43707
rect 15795 43673 15804 43707
rect 15752 43664 15804 43673
rect 17500 43664 17552 43716
rect 22284 43664 22336 43716
rect 23756 43732 23808 43784
rect 23848 43775 23900 43784
rect 23848 43741 23857 43775
rect 23857 43741 23891 43775
rect 23891 43741 23900 43775
rect 23848 43732 23900 43741
rect 24584 43775 24636 43784
rect 24584 43741 24593 43775
rect 24593 43741 24627 43775
rect 24627 43741 24636 43775
rect 24584 43732 24636 43741
rect 24676 43775 24728 43784
rect 24676 43741 24685 43775
rect 24685 43741 24719 43775
rect 24719 43741 24728 43775
rect 24676 43732 24728 43741
rect 26424 43732 26476 43784
rect 29828 43800 29880 43852
rect 32404 43800 32456 43852
rect 33324 43800 33376 43852
rect 35900 43800 35952 43852
rect 35992 43800 36044 43852
rect 28632 43775 28684 43784
rect 28632 43741 28641 43775
rect 28641 43741 28675 43775
rect 28675 43741 28684 43775
rect 28632 43732 28684 43741
rect 29000 43775 29052 43784
rect 28540 43664 28592 43716
rect 29000 43741 29009 43775
rect 29009 43741 29043 43775
rect 29043 43741 29052 43775
rect 29000 43732 29052 43741
rect 31576 43732 31628 43784
rect 32864 43775 32916 43784
rect 32864 43741 32873 43775
rect 32873 43741 32907 43775
rect 32907 43741 32916 43775
rect 32864 43732 32916 43741
rect 33140 43732 33192 43784
rect 10232 43596 10284 43648
rect 11704 43596 11756 43648
rect 11796 43596 11848 43648
rect 13360 43596 13412 43648
rect 13636 43596 13688 43648
rect 15200 43596 15252 43648
rect 16948 43596 17000 43648
rect 21272 43639 21324 43648
rect 21272 43605 21281 43639
rect 21281 43605 21315 43639
rect 21315 43605 21324 43639
rect 21272 43596 21324 43605
rect 23204 43596 23256 43648
rect 23296 43596 23348 43648
rect 28080 43596 28132 43648
rect 28264 43639 28316 43648
rect 28264 43605 28273 43639
rect 28273 43605 28307 43639
rect 28307 43605 28316 43639
rect 28264 43596 28316 43605
rect 29276 43596 29328 43648
rect 30380 43639 30432 43648
rect 30380 43605 30389 43639
rect 30389 43605 30423 43639
rect 30423 43605 30432 43639
rect 30380 43596 30432 43605
rect 31116 43596 31168 43648
rect 31852 43596 31904 43648
rect 34060 43664 34112 43716
rect 35256 43732 35308 43784
rect 35624 43732 35676 43784
rect 35716 43775 35768 43784
rect 35716 43741 35725 43775
rect 35725 43741 35759 43775
rect 35759 43741 35768 43775
rect 47308 43775 47360 43784
rect 35716 43732 35768 43741
rect 47308 43741 47317 43775
rect 47317 43741 47351 43775
rect 47351 43741 47360 43775
rect 47308 43732 47360 43741
rect 36268 43664 36320 43716
rect 36360 43664 36412 43716
rect 32496 43639 32548 43648
rect 32496 43605 32505 43639
rect 32505 43605 32539 43639
rect 32539 43605 32548 43639
rect 32496 43596 32548 43605
rect 34796 43596 34848 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 2320 43299 2372 43308
rect 2320 43265 2329 43299
rect 2329 43265 2363 43299
rect 2363 43265 2372 43299
rect 2320 43256 2372 43265
rect 2964 43392 3016 43444
rect 5816 43435 5868 43444
rect 2688 43299 2740 43308
rect 2688 43265 2697 43299
rect 2697 43265 2731 43299
rect 2731 43265 2740 43299
rect 2688 43256 2740 43265
rect 2872 43299 2924 43308
rect 2872 43265 2881 43299
rect 2881 43265 2915 43299
rect 2915 43265 2924 43299
rect 2872 43256 2924 43265
rect 3516 43299 3568 43308
rect 3516 43265 3525 43299
rect 3525 43265 3559 43299
rect 3559 43265 3568 43299
rect 3516 43256 3568 43265
rect 5448 43324 5500 43376
rect 5816 43401 5825 43435
rect 5825 43401 5859 43435
rect 5859 43401 5868 43435
rect 5816 43392 5868 43401
rect 6368 43392 6420 43444
rect 8116 43435 8168 43444
rect 8116 43401 8125 43435
rect 8125 43401 8159 43435
rect 8159 43401 8168 43435
rect 8116 43392 8168 43401
rect 9680 43392 9732 43444
rect 10048 43392 10100 43444
rect 11796 43324 11848 43376
rect 4712 43299 4764 43308
rect 4712 43265 4746 43299
rect 4746 43265 4764 43299
rect 4712 43256 4764 43265
rect 4988 43256 5040 43308
rect 6828 43256 6880 43308
rect 7012 43299 7064 43308
rect 7012 43265 7046 43299
rect 7046 43265 7064 43299
rect 8944 43299 8996 43308
rect 7012 43256 7064 43265
rect 8944 43265 8953 43299
rect 8953 43265 8987 43299
rect 8987 43265 8996 43299
rect 8944 43256 8996 43265
rect 10508 43256 10560 43308
rect 12164 43367 12216 43376
rect 12164 43333 12173 43367
rect 12173 43333 12207 43367
rect 12207 43333 12216 43367
rect 12164 43324 12216 43333
rect 12072 43256 12124 43308
rect 13636 43324 13688 43376
rect 13360 43299 13412 43308
rect 13360 43265 13394 43299
rect 13394 43265 13412 43299
rect 13360 43256 13412 43265
rect 13820 43392 13872 43444
rect 15200 43392 15252 43444
rect 15844 43392 15896 43444
rect 16672 43392 16724 43444
rect 17960 43392 18012 43444
rect 18696 43392 18748 43444
rect 16948 43367 17000 43376
rect 16948 43333 16982 43367
rect 16982 43333 17000 43367
rect 16948 43324 17000 43333
rect 848 43052 900 43104
rect 18604 43256 18656 43308
rect 2780 43120 2832 43172
rect 4804 43052 4856 43104
rect 9220 43095 9272 43104
rect 9220 43061 9229 43095
rect 9229 43061 9263 43095
rect 9263 43061 9272 43095
rect 9220 43052 9272 43061
rect 23112 43392 23164 43444
rect 23388 43392 23440 43444
rect 24952 43392 25004 43444
rect 26332 43435 26384 43444
rect 26332 43401 26341 43435
rect 26341 43401 26375 43435
rect 26375 43401 26384 43435
rect 26332 43392 26384 43401
rect 27528 43392 27580 43444
rect 29828 43392 29880 43444
rect 33140 43392 33192 43444
rect 33232 43392 33284 43444
rect 35072 43435 35124 43444
rect 35072 43401 35081 43435
rect 35081 43401 35115 43435
rect 35115 43401 35124 43435
rect 35072 43392 35124 43401
rect 36360 43435 36412 43444
rect 36360 43401 36369 43435
rect 36369 43401 36403 43435
rect 36403 43401 36412 43435
rect 36360 43392 36412 43401
rect 20628 43324 20680 43376
rect 19340 43256 19392 43308
rect 20168 43256 20220 43308
rect 20536 43299 20588 43308
rect 20536 43265 20545 43299
rect 20545 43265 20579 43299
rect 20579 43265 20588 43299
rect 20536 43256 20588 43265
rect 21088 43256 21140 43308
rect 21180 43256 21232 43308
rect 21916 43256 21968 43308
rect 23296 43324 23348 43376
rect 24860 43324 24912 43376
rect 28264 43324 28316 43376
rect 30104 43367 30156 43376
rect 30104 43333 30113 43367
rect 30113 43333 30147 43367
rect 30147 43333 30156 43367
rect 30104 43324 30156 43333
rect 32864 43324 32916 43376
rect 20628 43231 20680 43240
rect 20628 43197 20637 43231
rect 20637 43197 20671 43231
rect 20671 43197 20680 43231
rect 20628 43188 20680 43197
rect 19616 43052 19668 43104
rect 20352 43120 20404 43172
rect 23204 43299 23256 43308
rect 23204 43265 23238 43299
rect 23238 43265 23256 43299
rect 23204 43256 23256 43265
rect 25228 43299 25280 43308
rect 25228 43265 25262 43299
rect 25262 43265 25280 43299
rect 25228 43256 25280 43265
rect 27988 43188 28040 43240
rect 28908 43256 28960 43308
rect 31576 43299 31628 43308
rect 31576 43265 31585 43299
rect 31585 43265 31619 43299
rect 31619 43265 31628 43299
rect 31576 43256 31628 43265
rect 32404 43299 32456 43308
rect 32404 43265 32413 43299
rect 32413 43265 32447 43299
rect 32447 43265 32456 43299
rect 32404 43256 32456 43265
rect 33140 43256 33192 43308
rect 35716 43256 35768 43308
rect 35900 43299 35952 43308
rect 35900 43265 35909 43299
rect 35909 43265 35943 43299
rect 35943 43265 35952 43299
rect 35900 43256 35952 43265
rect 38660 43256 38712 43308
rect 46940 43256 46992 43308
rect 31944 43188 31996 43240
rect 35256 43188 35308 43240
rect 36084 43188 36136 43240
rect 21088 43095 21140 43104
rect 21088 43061 21097 43095
rect 21097 43061 21131 43095
rect 21131 43061 21140 43095
rect 21088 43052 21140 43061
rect 21364 43052 21416 43104
rect 35348 43120 35400 43172
rect 48044 43163 48096 43172
rect 48044 43129 48053 43163
rect 48053 43129 48087 43163
rect 48087 43129 48096 43163
rect 48044 43120 48096 43129
rect 31300 43052 31352 43104
rect 46940 43095 46992 43104
rect 46940 43061 46949 43095
rect 46949 43061 46983 43095
rect 46983 43061 46992 43095
rect 46940 43052 46992 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 4712 42848 4764 42900
rect 7012 42848 7064 42900
rect 8944 42848 8996 42900
rect 10508 42891 10560 42900
rect 10508 42857 10517 42891
rect 10517 42857 10551 42891
rect 10551 42857 10560 42891
rect 10508 42848 10560 42857
rect 11980 42891 12032 42900
rect 11980 42857 11989 42891
rect 11989 42857 12023 42891
rect 12023 42857 12032 42891
rect 11980 42848 12032 42857
rect 2320 42780 2372 42832
rect 2688 42755 2740 42764
rect 2688 42721 2697 42755
rect 2697 42721 2731 42755
rect 2731 42721 2740 42755
rect 2688 42712 2740 42721
rect 2596 42644 2648 42696
rect 4252 42780 4304 42832
rect 4620 42780 4672 42832
rect 9220 42780 9272 42832
rect 4528 42712 4580 42764
rect 2780 42653 2814 42674
rect 2814 42653 2832 42674
rect 2780 42622 2832 42653
rect 4712 42644 4764 42696
rect 4896 42644 4948 42696
rect 6736 42755 6788 42764
rect 6736 42721 6745 42755
rect 6745 42721 6779 42755
rect 6779 42721 6788 42755
rect 6736 42712 6788 42721
rect 2320 42551 2372 42560
rect 2320 42517 2329 42551
rect 2329 42517 2363 42551
rect 2363 42517 2372 42551
rect 2320 42508 2372 42517
rect 3240 42508 3292 42560
rect 5816 42644 5868 42696
rect 6368 42687 6420 42696
rect 6368 42653 6377 42687
rect 6377 42653 6411 42687
rect 6411 42653 6420 42687
rect 6368 42644 6420 42653
rect 6552 42687 6604 42696
rect 6552 42653 6561 42687
rect 6561 42653 6595 42687
rect 6595 42653 6604 42687
rect 6552 42644 6604 42653
rect 8116 42712 8168 42764
rect 17132 42712 17184 42764
rect 20628 42848 20680 42900
rect 20996 42891 21048 42900
rect 20996 42857 21005 42891
rect 21005 42857 21039 42891
rect 21039 42857 21048 42891
rect 20996 42848 21048 42857
rect 23296 42891 23348 42900
rect 23296 42857 23305 42891
rect 23305 42857 23339 42891
rect 23339 42857 23348 42891
rect 23296 42848 23348 42857
rect 25228 42848 25280 42900
rect 30104 42848 30156 42900
rect 34060 42891 34112 42900
rect 34060 42857 34069 42891
rect 34069 42857 34103 42891
rect 34103 42857 34112 42891
rect 34060 42848 34112 42857
rect 41512 42848 41564 42900
rect 36268 42823 36320 42832
rect 36268 42789 36277 42823
rect 36277 42789 36311 42823
rect 36311 42789 36320 42823
rect 36268 42780 36320 42789
rect 19340 42712 19392 42764
rect 19616 42755 19668 42764
rect 19616 42721 19625 42755
rect 19625 42721 19659 42755
rect 19659 42721 19668 42755
rect 19616 42712 19668 42721
rect 21916 42755 21968 42764
rect 21916 42721 21925 42755
rect 21925 42721 21959 42755
rect 21959 42721 21968 42755
rect 21916 42712 21968 42721
rect 24768 42755 24820 42764
rect 24768 42721 24777 42755
rect 24777 42721 24811 42755
rect 24811 42721 24820 42755
rect 24768 42712 24820 42721
rect 8208 42687 8260 42696
rect 7104 42576 7156 42628
rect 8208 42653 8217 42687
rect 8217 42653 8251 42687
rect 8251 42653 8260 42687
rect 8208 42644 8260 42653
rect 9128 42644 9180 42696
rect 10508 42687 10560 42696
rect 10508 42653 10517 42687
rect 10517 42653 10551 42687
rect 10551 42653 10560 42687
rect 10508 42644 10560 42653
rect 17408 42644 17460 42696
rect 6368 42508 6420 42560
rect 7748 42551 7800 42560
rect 7748 42517 7757 42551
rect 7757 42517 7791 42551
rect 7791 42517 7800 42551
rect 7748 42508 7800 42517
rect 9680 42551 9732 42560
rect 9680 42517 9689 42551
rect 9689 42517 9723 42551
rect 9723 42517 9732 42551
rect 9680 42508 9732 42517
rect 18696 42644 18748 42696
rect 21088 42644 21140 42696
rect 23848 42644 23900 42696
rect 18328 42576 18380 42628
rect 23388 42619 23440 42628
rect 23388 42585 23397 42619
rect 23397 42585 23431 42619
rect 23431 42585 23440 42619
rect 23388 42576 23440 42585
rect 24216 42576 24268 42628
rect 18512 42508 18564 42560
rect 23572 42508 23624 42560
rect 26332 42644 26384 42696
rect 26792 42644 26844 42696
rect 31116 42644 31168 42696
rect 32680 42687 32732 42696
rect 32680 42653 32689 42687
rect 32689 42653 32723 42687
rect 32723 42653 32732 42687
rect 32680 42644 32732 42653
rect 32496 42576 32548 42628
rect 34796 42576 34848 42628
rect 30472 42508 30524 42560
rect 31944 42551 31996 42560
rect 31944 42517 31953 42551
rect 31953 42517 31987 42551
rect 31987 42517 31996 42551
rect 31944 42508 31996 42517
rect 47308 42551 47360 42560
rect 47308 42517 47317 42551
rect 47317 42517 47351 42551
rect 47351 42517 47360 42551
rect 47308 42508 47360 42517
rect 48044 42551 48096 42560
rect 48044 42517 48053 42551
rect 48053 42517 48087 42551
rect 48087 42517 48096 42551
rect 48044 42508 48096 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 4252 42347 4304 42356
rect 4252 42313 4261 42347
rect 4261 42313 4295 42347
rect 4295 42313 4304 42347
rect 4252 42304 4304 42313
rect 2320 42236 2372 42288
rect 1952 42168 2004 42220
rect 4988 42304 5040 42356
rect 6920 42304 6972 42356
rect 9956 42304 10008 42356
rect 10140 42304 10192 42356
rect 10508 42304 10560 42356
rect 26792 42304 26844 42356
rect 9128 42279 9180 42288
rect 9128 42245 9137 42279
rect 9137 42245 9171 42279
rect 9171 42245 9180 42279
rect 9128 42236 9180 42245
rect 20076 42236 20128 42288
rect 20536 42236 20588 42288
rect 14464 42168 14516 42220
rect 12440 42100 12492 42152
rect 27988 42168 28040 42220
rect 32680 42236 32732 42288
rect 30472 42211 30524 42220
rect 30472 42177 30506 42211
rect 30506 42177 30524 42211
rect 30472 42168 30524 42177
rect 2596 42032 2648 42084
rect 1492 42007 1544 42016
rect 1492 41973 1501 42007
rect 1501 41973 1535 42007
rect 1535 41973 1544 42007
rect 1492 41964 1544 41973
rect 6552 41964 6604 42016
rect 24216 42007 24268 42016
rect 24216 41973 24225 42007
rect 24225 41973 24259 42007
rect 24259 41973 24268 42007
rect 24216 41964 24268 41973
rect 31576 42007 31628 42016
rect 31576 41973 31585 42007
rect 31585 41973 31619 42007
rect 31619 41973 31628 42007
rect 31576 41964 31628 41973
rect 34704 41964 34756 42016
rect 48044 42007 48096 42016
rect 48044 41973 48053 42007
rect 48053 41973 48087 42007
rect 48087 41973 48096 42007
rect 48044 41964 48096 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1952 41803 2004 41812
rect 1952 41769 1961 41803
rect 1961 41769 1995 41803
rect 1995 41769 2004 41803
rect 1952 41760 2004 41769
rect 4712 41760 4764 41812
rect 12256 41760 12308 41812
rect 47308 41760 47360 41812
rect 2780 41692 2832 41744
rect 9680 41692 9732 41744
rect 31116 41735 31168 41744
rect 31116 41701 31125 41735
rect 31125 41701 31159 41735
rect 31159 41701 31168 41735
rect 31116 41692 31168 41701
rect 31852 41624 31904 41676
rect 2596 41556 2648 41608
rect 9220 41556 9272 41608
rect 30748 41556 30800 41608
rect 31300 41599 31352 41608
rect 31300 41565 31309 41599
rect 31309 41565 31343 41599
rect 31343 41565 31352 41599
rect 31300 41556 31352 41565
rect 31668 41599 31720 41608
rect 31668 41565 31677 41599
rect 31677 41565 31711 41599
rect 31711 41565 31720 41599
rect 31668 41556 31720 41565
rect 48044 41599 48096 41608
rect 48044 41565 48053 41599
rect 48053 41565 48087 41599
rect 48087 41565 48096 41599
rect 48044 41556 48096 41565
rect 31944 41488 31996 41540
rect 46296 41488 46348 41540
rect 24584 41420 24636 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 30748 41259 30800 41268
rect 30748 41225 30757 41259
rect 30757 41225 30791 41259
rect 30791 41225 30800 41259
rect 30748 41216 30800 41225
rect 48044 41123 48096 41132
rect 48044 41089 48053 41123
rect 48053 41089 48087 41123
rect 48087 41089 48096 41123
rect 48044 41080 48096 41089
rect 47032 40944 47084 40996
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 18604 40672 18656 40724
rect 46940 40672 46992 40724
rect 48044 40672 48096 40724
rect 48044 40375 48096 40384
rect 48044 40341 48053 40375
rect 48053 40341 48087 40375
rect 48087 40341 48096 40375
rect 48044 40332 48096 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 15200 40060 15252 40112
rect 48044 40103 48096 40112
rect 48044 40069 48053 40103
rect 48053 40069 48087 40103
rect 48087 40069 48096 40103
rect 48044 40060 48096 40069
rect 11980 39992 12032 40044
rect 48136 39788 48188 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 48044 39355 48096 39364
rect 48044 39321 48053 39355
rect 48053 39321 48087 39355
rect 48087 39321 48096 39355
rect 48044 39312 48096 39321
rect 45560 39244 45612 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 48044 38947 48096 38956
rect 48044 38913 48053 38947
rect 48053 38913 48087 38947
rect 48087 38913 48096 38947
rect 48044 38904 48096 38913
rect 47768 38768 47820 38820
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 27988 38471 28040 38480
rect 27988 38437 27997 38471
rect 27997 38437 28031 38471
rect 28031 38437 28040 38471
rect 27988 38428 28040 38437
rect 23388 38224 23440 38276
rect 48044 38267 48096 38276
rect 48044 38233 48053 38267
rect 48053 38233 48087 38267
rect 48087 38233 48096 38267
rect 48044 38224 48096 38233
rect 46572 38156 46624 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 48044 37859 48096 37868
rect 48044 37825 48053 37859
rect 48053 37825 48087 37859
rect 48087 37825 48096 37859
rect 48044 37816 48096 37825
rect 47860 37723 47912 37732
rect 47860 37689 47869 37723
rect 47869 37689 47903 37723
rect 47903 37689 47912 37723
rect 47860 37680 47912 37689
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 48044 37408 48096 37460
rect 48044 37111 48096 37120
rect 48044 37077 48053 37111
rect 48053 37077 48087 37111
rect 48087 37077 48096 37111
rect 48044 37068 48096 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 48044 36771 48096 36780
rect 48044 36737 48053 36771
rect 48053 36737 48087 36771
rect 48087 36737 48096 36771
rect 48044 36728 48096 36737
rect 45836 36592 45888 36644
rect 11152 36524 11204 36576
rect 24216 36524 24268 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 9956 36363 10008 36372
rect 9956 36329 9965 36363
rect 9965 36329 9999 36363
rect 9999 36329 10008 36363
rect 9956 36320 10008 36329
rect 11152 36116 11204 36168
rect 15200 36048 15252 36100
rect 48044 36091 48096 36100
rect 48044 36057 48053 36091
rect 48053 36057 48087 36091
rect 48087 36057 48096 36091
rect 48044 36048 48096 36057
rect 1492 36023 1544 36032
rect 1492 35989 1501 36023
rect 1501 35989 1535 36023
rect 1535 35989 1544 36023
rect 1492 35980 1544 35989
rect 47952 36023 48004 36032
rect 47952 35989 47961 36023
rect 47961 35989 47995 36023
rect 47995 35989 48004 36023
rect 47952 35980 48004 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 48044 35683 48096 35692
rect 48044 35649 48053 35683
rect 48053 35649 48087 35683
rect 48087 35649 48096 35683
rect 48044 35640 48096 35649
rect 45928 35504 45980 35556
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 48044 35003 48096 35012
rect 48044 34969 48053 35003
rect 48053 34969 48087 35003
rect 48087 34969 48096 35003
rect 48044 34960 48096 34969
rect 47124 34892 47176 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 48044 34595 48096 34604
rect 48044 34561 48053 34595
rect 48053 34561 48087 34595
rect 48087 34561 48096 34595
rect 48044 34552 48096 34561
rect 47584 34484 47636 34536
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 48044 34144 48096 34196
rect 48044 33847 48096 33856
rect 48044 33813 48053 33847
rect 48053 33813 48087 33847
rect 48087 33813 48096 33847
rect 48044 33804 48096 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 48044 33507 48096 33516
rect 48044 33473 48053 33507
rect 48053 33473 48087 33507
rect 48087 33473 48096 33507
rect 48044 33464 48096 33473
rect 47400 33328 47452 33380
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 48044 32827 48096 32836
rect 48044 32793 48053 32827
rect 48053 32793 48087 32827
rect 48087 32793 48096 32827
rect 48044 32784 48096 32793
rect 47216 32716 47268 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 23388 32487 23440 32496
rect 23388 32453 23397 32487
rect 23397 32453 23431 32487
rect 23431 32453 23440 32487
rect 23388 32444 23440 32453
rect 19892 32376 19944 32428
rect 48044 32419 48096 32428
rect 48044 32385 48053 32419
rect 48053 32385 48087 32419
rect 48087 32385 48096 32419
rect 48044 32376 48096 32385
rect 46020 32240 46072 32292
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 15200 31900 15252 31952
rect 19892 31764 19944 31816
rect 48044 31807 48096 31816
rect 48044 31773 48053 31807
rect 48053 31773 48087 31807
rect 48087 31773 48096 31807
rect 48044 31764 48096 31773
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 48044 31331 48096 31340
rect 48044 31297 48053 31331
rect 48053 31297 48087 31331
rect 48087 31297 48096 31331
rect 48044 31288 48096 31297
rect 45652 31152 45704 31204
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 48044 30880 48096 30932
rect 1492 30583 1544 30592
rect 1492 30549 1501 30583
rect 1501 30549 1535 30583
rect 1535 30549 1544 30583
rect 1492 30540 1544 30549
rect 2872 30583 2924 30592
rect 2872 30549 2881 30583
rect 2881 30549 2915 30583
rect 2915 30549 2924 30583
rect 2872 30540 2924 30549
rect 17224 30540 17276 30592
rect 48044 30583 48096 30592
rect 48044 30549 48053 30583
rect 48053 30549 48087 30583
rect 48087 30549 48096 30583
rect 48044 30540 48096 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 48044 30243 48096 30252
rect 48044 30209 48053 30243
rect 48053 30209 48087 30243
rect 48087 30209 48096 30243
rect 48044 30200 48096 30209
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 48044 29563 48096 29572
rect 48044 29529 48053 29563
rect 48053 29529 48087 29563
rect 48087 29529 48096 29563
rect 48044 29520 48096 29529
rect 45744 29452 45796 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 48044 29155 48096 29164
rect 48044 29121 48053 29155
rect 48053 29121 48087 29155
rect 48087 29121 48096 29155
rect 48044 29112 48096 29121
rect 46664 28976 46716 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 48044 28475 48096 28484
rect 48044 28441 48053 28475
rect 48053 28441 48087 28475
rect 48087 28441 48096 28475
rect 48044 28432 48096 28441
rect 44640 28364 44692 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 48228 28024 48280 28076
rect 48320 27820 48372 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 48228 27548 48280 27600
rect 48044 27276 48096 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 48044 26979 48096 26988
rect 48044 26945 48053 26979
rect 48053 26945 48087 26979
rect 48087 26945 48096 26979
rect 48044 26936 48096 26945
rect 47308 26868 47360 26920
rect 47768 26868 47820 26920
rect 47952 26868 48004 26920
rect 48228 26868 48280 26920
rect 47032 26800 47084 26852
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 47952 26571 48004 26580
rect 47952 26537 47961 26571
rect 47961 26537 47995 26571
rect 47995 26537 48004 26571
rect 47952 26528 48004 26537
rect 48044 26299 48096 26308
rect 48044 26265 48053 26299
rect 48053 26265 48087 26299
rect 48087 26265 48096 26299
rect 48044 26256 48096 26265
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 48044 25891 48096 25900
rect 48044 25857 48053 25891
rect 48053 25857 48087 25891
rect 48087 25857 48096 25891
rect 48044 25848 48096 25857
rect 47676 25712 47728 25764
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19984 25347 20036 25356
rect 19984 25313 19993 25347
rect 19993 25313 20027 25347
rect 20027 25313 20036 25347
rect 19984 25304 20036 25313
rect 1676 25279 1728 25288
rect 1676 25245 1685 25279
rect 1685 25245 1719 25279
rect 1719 25245 1728 25279
rect 1676 25236 1728 25245
rect 48044 25211 48096 25220
rect 1492 25143 1544 25152
rect 1492 25109 1501 25143
rect 1501 25109 1535 25143
rect 1535 25109 1544 25143
rect 1492 25100 1544 25109
rect 48044 25177 48053 25211
rect 48053 25177 48087 25211
rect 48087 25177 48096 25211
rect 48044 25168 48096 25177
rect 28540 25100 28592 25152
rect 47492 25100 47544 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1676 24896 1728 24948
rect 2688 24760 2740 24812
rect 8300 24760 8352 24812
rect 48044 24803 48096 24812
rect 48044 24769 48053 24803
rect 48053 24769 48087 24803
rect 48087 24769 48096 24803
rect 48044 24760 48096 24769
rect 47860 24667 47912 24676
rect 47860 24633 47869 24667
rect 47869 24633 47903 24667
rect 47903 24633 47912 24667
rect 47860 24624 47912 24633
rect 2688 24599 2740 24608
rect 2688 24565 2697 24599
rect 2697 24565 2731 24599
rect 2731 24565 2740 24599
rect 2688 24556 2740 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 48044 24123 48096 24132
rect 48044 24089 48053 24123
rect 48053 24089 48087 24123
rect 48087 24089 48096 24123
rect 48044 24080 48096 24089
rect 45376 24012 45428 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 48044 23035 48096 23044
rect 48044 23001 48053 23035
rect 48053 23001 48087 23035
rect 48087 23001 48096 23035
rect 48044 22992 48096 23001
rect 44272 22924 44324 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 48044 22627 48096 22636
rect 48044 22593 48053 22627
rect 48053 22593 48087 22627
rect 48087 22593 48096 22627
rect 48044 22584 48096 22593
rect 47768 22448 47820 22500
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 48228 22108 48280 22160
rect 48412 22108 48464 22160
rect 48044 22040 48096 22092
rect 47952 21972 48004 22024
rect 48228 21972 48280 22024
rect 48044 21947 48096 21956
rect 48044 21913 48053 21947
rect 48053 21913 48087 21947
rect 48087 21913 48096 21947
rect 48044 21904 48096 21913
rect 45468 21836 45520 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 48228 21632 48280 21684
rect 48044 21539 48096 21548
rect 48044 21505 48053 21539
rect 48053 21505 48087 21539
rect 48087 21505 48096 21539
rect 48044 21496 48096 21505
rect 47952 21428 48004 21480
rect 48136 21360 48188 21412
rect 45836 21292 45888 21344
rect 46112 21292 46164 21344
rect 46756 21292 46808 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 45928 21020 45980 21072
rect 47492 20927 47544 20936
rect 47492 20893 47501 20927
rect 47501 20893 47535 20927
rect 47535 20893 47544 20927
rect 47492 20884 47544 20893
rect 48136 20927 48188 20936
rect 48136 20893 48145 20927
rect 48145 20893 48179 20927
rect 48179 20893 48188 20927
rect 48136 20884 48188 20893
rect 46480 20816 46532 20868
rect 46848 20791 46900 20800
rect 46848 20757 46857 20791
rect 46857 20757 46891 20791
rect 46891 20757 46900 20791
rect 46848 20748 46900 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1216 20544 1268 20596
rect 2596 20544 2648 20596
rect 46296 20544 46348 20596
rect 47952 20544 48004 20596
rect 48228 20544 48280 20596
rect 46848 20408 46900 20460
rect 48228 20408 48280 20460
rect 47584 20204 47636 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 40684 19932 40736 19984
rect 47768 19864 47820 19916
rect 1952 19796 2004 19848
rect 45928 19839 45980 19848
rect 44824 19728 44876 19780
rect 45928 19805 45937 19839
rect 45937 19805 45971 19839
rect 45971 19805 45980 19839
rect 45928 19796 45980 19805
rect 46296 19839 46348 19848
rect 46296 19805 46305 19839
rect 46305 19805 46339 19839
rect 46339 19805 46348 19839
rect 46296 19796 46348 19805
rect 46388 19839 46440 19848
rect 46388 19805 46397 19839
rect 46397 19805 46431 19839
rect 46431 19805 46440 19839
rect 46388 19796 46440 19805
rect 46848 19796 46900 19848
rect 47584 19839 47636 19848
rect 47584 19805 47593 19839
rect 47593 19805 47627 19839
rect 47627 19805 47636 19839
rect 47584 19796 47636 19805
rect 47952 19839 48004 19848
rect 47952 19805 47961 19839
rect 47961 19805 47995 19839
rect 47995 19805 48004 19839
rect 47952 19796 48004 19805
rect 46204 19728 46256 19780
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 6552 19456 6604 19508
rect 14556 19388 14608 19440
rect 40684 19388 40736 19440
rect 46388 19388 46440 19440
rect 1124 19252 1176 19304
rect 39304 19320 39356 19372
rect 46204 19320 46256 19372
rect 46480 19363 46532 19372
rect 46480 19329 46489 19363
rect 46489 19329 46523 19363
rect 46523 19329 46532 19363
rect 46480 19320 46532 19329
rect 46940 19320 46992 19372
rect 48044 19320 48096 19372
rect 47400 19184 47452 19236
rect 48136 19184 48188 19236
rect 47584 19116 47636 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 47124 18912 47176 18964
rect 47400 18912 47452 18964
rect 47216 18844 47268 18896
rect 45928 18776 45980 18828
rect 46848 18776 46900 18828
rect 47768 18776 47820 18828
rect 46296 18751 46348 18760
rect 46296 18717 46305 18751
rect 46305 18717 46339 18751
rect 46339 18717 46348 18751
rect 46296 18708 46348 18717
rect 47584 18751 47636 18760
rect 47584 18717 47593 18751
rect 47593 18717 47627 18751
rect 47627 18717 47636 18751
rect 47584 18708 47636 18717
rect 46480 18615 46532 18624
rect 46480 18581 46489 18615
rect 46489 18581 46523 18615
rect 46523 18581 46532 18615
rect 46480 18572 46532 18581
rect 47032 18615 47084 18624
rect 47032 18581 47041 18615
rect 47041 18581 47075 18615
rect 47075 18581 47084 18615
rect 47032 18572 47084 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 16120 18368 16172 18420
rect 47032 18368 47084 18420
rect 45560 18232 45612 18284
rect 46112 18232 46164 18284
rect 46296 18232 46348 18284
rect 46480 18275 46532 18284
rect 46480 18241 46489 18275
rect 46489 18241 46523 18275
rect 46523 18241 46532 18275
rect 46480 18232 46532 18241
rect 45928 18164 45980 18216
rect 46112 18071 46164 18080
rect 46112 18037 46121 18071
rect 46121 18037 46155 18071
rect 46155 18037 46164 18071
rect 46112 18028 46164 18037
rect 47768 18232 47820 18284
rect 48136 18275 48188 18284
rect 48136 18241 48145 18275
rect 48145 18241 48179 18275
rect 48179 18241 48188 18275
rect 48136 18232 48188 18241
rect 47584 18028 47636 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 47952 17756 48004 17808
rect 46848 17688 46900 17740
rect 47768 17688 47820 17740
rect 47952 17663 48004 17672
rect 45560 17552 45612 17604
rect 45836 17552 45888 17604
rect 46480 17552 46532 17604
rect 47952 17629 47961 17663
rect 47961 17629 47995 17663
rect 47995 17629 48004 17663
rect 47952 17620 48004 17629
rect 45928 17527 45980 17536
rect 45928 17493 45937 17527
rect 45937 17493 45971 17527
rect 45971 17493 45980 17527
rect 45928 17484 45980 17493
rect 46572 17484 46624 17536
rect 46756 17484 46808 17536
rect 47032 17527 47084 17536
rect 47032 17493 47041 17527
rect 47041 17493 47075 17527
rect 47075 17493 47084 17527
rect 47032 17484 47084 17493
rect 47952 17484 48004 17536
rect 48228 17484 48280 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 45928 17280 45980 17332
rect 14004 17212 14056 17264
rect 47032 17212 47084 17264
rect 47124 17212 47176 17264
rect 47492 17212 47544 17264
rect 45652 17076 45704 17128
rect 45928 17076 45980 17128
rect 46756 17144 46808 17196
rect 47768 17144 47820 17196
rect 48228 17144 48280 17196
rect 47584 17076 47636 17128
rect 46756 17008 46808 17060
rect 46572 16940 46624 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 46296 16736 46348 16788
rect 46480 16779 46532 16788
rect 46480 16745 46489 16779
rect 46489 16745 46523 16779
rect 46523 16745 46532 16779
rect 46480 16736 46532 16745
rect 46296 16575 46348 16584
rect 46296 16541 46305 16575
rect 46305 16541 46339 16575
rect 46339 16541 46348 16575
rect 46296 16532 46348 16541
rect 47400 16575 47452 16584
rect 47400 16541 47409 16575
rect 47409 16541 47443 16575
rect 47443 16541 47452 16575
rect 47400 16532 47452 16541
rect 47584 16575 47636 16584
rect 47584 16541 47593 16575
rect 47593 16541 47627 16575
rect 47627 16541 47636 16575
rect 47584 16532 47636 16541
rect 48044 16575 48096 16584
rect 48044 16541 48053 16575
rect 48053 16541 48087 16575
rect 48087 16541 48096 16575
rect 48044 16532 48096 16541
rect 45928 16464 45980 16516
rect 46848 16464 46900 16516
rect 47032 16439 47084 16448
rect 47032 16405 47041 16439
rect 47041 16405 47075 16439
rect 47075 16405 47084 16439
rect 47032 16396 47084 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 13268 16192 13320 16244
rect 47032 16192 47084 16244
rect 47768 16235 47820 16244
rect 47768 16201 47777 16235
rect 47777 16201 47811 16235
rect 47811 16201 47820 16235
rect 47768 16192 47820 16201
rect 45928 16099 45980 16108
rect 45928 16065 45937 16099
rect 45937 16065 45971 16099
rect 45971 16065 45980 16099
rect 45928 16056 45980 16065
rect 46480 16056 46532 16108
rect 46756 16056 46808 16108
rect 47584 15920 47636 15972
rect 46296 15852 46348 15904
rect 46848 15852 46900 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 48136 15648 48188 15700
rect 46020 15580 46072 15632
rect 46480 15580 46532 15632
rect 33140 15512 33192 15564
rect 47400 15555 47452 15564
rect 47400 15521 47409 15555
rect 47409 15521 47443 15555
rect 47443 15521 47452 15555
rect 47400 15512 47452 15521
rect 47492 15512 47544 15564
rect 46296 15487 46348 15496
rect 46296 15453 46305 15487
rect 46305 15453 46339 15487
rect 46339 15453 46348 15487
rect 46296 15444 46348 15453
rect 48044 15487 48096 15496
rect 48044 15453 48053 15487
rect 48053 15453 48087 15487
rect 48087 15453 48096 15487
rect 48044 15444 48096 15453
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 45560 15104 45612 15156
rect 46848 15104 46900 15156
rect 45560 14968 45612 15020
rect 46572 14968 46624 15020
rect 48412 15036 48464 15088
rect 47032 15011 47084 15020
rect 47032 14977 47041 15011
rect 47041 14977 47075 15011
rect 47075 14977 47084 15011
rect 47032 14968 47084 14977
rect 48044 14968 48096 15020
rect 48136 15011 48188 15020
rect 48136 14977 48145 15011
rect 48145 14977 48179 15011
rect 48179 14977 48188 15011
rect 48136 14968 48188 14977
rect 37924 14900 37976 14952
rect 47400 14900 47452 14952
rect 46480 14764 46532 14816
rect 47584 14764 47636 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 47032 14560 47084 14612
rect 47400 14467 47452 14476
rect 47400 14433 47409 14467
rect 47409 14433 47443 14467
rect 47443 14433 47452 14467
rect 47400 14424 47452 14433
rect 46020 14356 46072 14408
rect 46756 14356 46808 14408
rect 47584 14399 47636 14408
rect 47584 14365 47593 14399
rect 47593 14365 47627 14399
rect 47627 14365 47636 14399
rect 47584 14356 47636 14365
rect 47768 14356 47820 14408
rect 48044 14399 48096 14408
rect 48044 14365 48053 14399
rect 48053 14365 48087 14399
rect 48087 14365 48096 14399
rect 48044 14356 48096 14365
rect 27344 14288 27396 14340
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 47768 14016 47820 14068
rect 46480 13923 46532 13932
rect 664 13812 716 13864
rect 46480 13889 46489 13923
rect 46489 13889 46523 13923
rect 46523 13889 46532 13923
rect 46480 13880 46532 13889
rect 46848 13923 46900 13932
rect 46848 13889 46857 13923
rect 46857 13889 46891 13923
rect 46891 13889 46900 13923
rect 46848 13880 46900 13889
rect 47032 13923 47084 13932
rect 47032 13889 47041 13923
rect 47041 13889 47075 13923
rect 47075 13889 47084 13923
rect 47032 13880 47084 13889
rect 48044 13880 48096 13932
rect 4620 13812 4672 13864
rect 36636 13812 36688 13864
rect 47400 13812 47452 13864
rect 1492 13787 1544 13796
rect 1492 13753 1501 13787
rect 1501 13753 1535 13787
rect 1535 13753 1544 13787
rect 1492 13744 1544 13753
rect 47584 13676 47636 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 48044 13472 48096 13524
rect 48228 13472 48280 13524
rect 46940 13336 46992 13388
rect 46296 13311 46348 13320
rect 46296 13277 46305 13311
rect 46305 13277 46339 13311
rect 46339 13277 46348 13311
rect 46296 13268 46348 13277
rect 46572 13268 46624 13320
rect 47584 13311 47636 13320
rect 47584 13277 47593 13311
rect 47593 13277 47627 13311
rect 47627 13277 47636 13311
rect 47584 13268 47636 13277
rect 48044 13311 48096 13320
rect 48044 13277 48053 13311
rect 48053 13277 48087 13311
rect 48087 13277 48096 13311
rect 48044 13268 48096 13277
rect 46480 13175 46532 13184
rect 46480 13141 46489 13175
rect 46489 13141 46523 13175
rect 46523 13141 46532 13175
rect 46480 13132 46532 13141
rect 47032 13175 47084 13184
rect 47032 13141 47041 13175
rect 47041 13141 47075 13175
rect 47075 13141 47084 13175
rect 47032 13132 47084 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 8300 12928 8352 12980
rect 47032 12928 47084 12980
rect 45192 12860 45244 12912
rect 45836 12860 45888 12912
rect 46480 12835 46532 12844
rect 46480 12801 46489 12835
rect 46489 12801 46523 12835
rect 46523 12801 46532 12835
rect 46480 12792 46532 12801
rect 47952 12860 48004 12912
rect 46940 12792 46992 12844
rect 48044 12792 48096 12844
rect 45652 12724 45704 12776
rect 46572 12767 46624 12776
rect 46572 12733 46581 12767
rect 46581 12733 46615 12767
rect 46615 12733 46624 12767
rect 46572 12724 46624 12733
rect 46020 12588 46072 12640
rect 46388 12588 46440 12640
rect 46848 12656 46900 12708
rect 46756 12588 46808 12640
rect 47584 12588 47636 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 45284 12384 45336 12436
rect 46020 12248 46072 12300
rect 46572 12248 46624 12300
rect 46296 12223 46348 12232
rect 46296 12189 46305 12223
rect 46305 12189 46339 12223
rect 46339 12189 46348 12223
rect 46296 12180 46348 12189
rect 46480 12180 46532 12232
rect 46848 12180 46900 12232
rect 47584 12223 47636 12232
rect 47584 12189 47593 12223
rect 47593 12189 47627 12223
rect 47627 12189 47636 12223
rect 47584 12180 47636 12189
rect 48044 12248 48096 12300
rect 45560 12044 45612 12096
rect 46020 12044 46072 12096
rect 46112 12044 46164 12096
rect 47032 12087 47084 12096
rect 47032 12053 47041 12087
rect 47041 12053 47075 12087
rect 47075 12053 47084 12087
rect 47032 12044 47084 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 25228 11840 25280 11892
rect 47032 11840 47084 11892
rect 45928 11772 45980 11824
rect 45284 11704 45336 11756
rect 46940 11747 46992 11756
rect 46940 11713 46949 11747
rect 46949 11713 46983 11747
rect 46983 11713 46992 11747
rect 48136 11747 48188 11756
rect 46940 11704 46992 11713
rect 48136 11713 48145 11747
rect 48145 11713 48179 11747
rect 48179 11713 48188 11747
rect 48136 11704 48188 11713
rect 45560 11636 45612 11688
rect 46848 11568 46900 11620
rect 1860 11500 1912 11552
rect 48136 11568 48188 11620
rect 47584 11500 47636 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 46940 11296 46992 11348
rect 45928 11228 45980 11280
rect 46112 11228 46164 11280
rect 45744 11203 45796 11212
rect 45744 11169 45753 11203
rect 45753 11169 45787 11203
rect 45787 11169 45796 11203
rect 45744 11160 45796 11169
rect 45836 11092 45888 11144
rect 46112 11092 46164 11144
rect 46848 11160 46900 11212
rect 47584 11135 47636 11144
rect 1584 11024 1636 11076
rect 2596 11067 2648 11076
rect 2596 11033 2605 11067
rect 2605 11033 2639 11067
rect 2639 11033 2648 11067
rect 2596 11024 2648 11033
rect 3424 11024 3476 11076
rect 3976 11024 4028 11076
rect 4620 11024 4672 11076
rect 5448 11024 5500 11076
rect 15292 11024 15344 11076
rect 47584 11101 47593 11135
rect 47593 11101 47627 11135
rect 47627 11101 47636 11135
rect 47584 11092 47636 11101
rect 48044 11135 48096 11144
rect 48044 11101 48053 11135
rect 48053 11101 48087 11135
rect 48087 11101 48096 11135
rect 48044 11092 48096 11101
rect 45192 10956 45244 11008
rect 45744 10956 45796 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 46848 10752 46900 10804
rect 45928 10616 45980 10668
rect 46388 10616 46440 10668
rect 48228 10616 48280 10668
rect 3884 10480 3936 10532
rect 1676 10412 1728 10464
rect 2136 10412 2188 10464
rect 2228 10412 2280 10464
rect 3516 10412 3568 10464
rect 4068 10412 4120 10464
rect 4712 10412 4764 10464
rect 5356 10455 5408 10464
rect 5356 10421 5365 10455
rect 5365 10421 5399 10455
rect 5399 10421 5408 10455
rect 5356 10412 5408 10421
rect 46940 10412 46992 10464
rect 47584 10412 47636 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 45744 10251 45796 10260
rect 45744 10217 45753 10251
rect 45753 10217 45787 10251
rect 45787 10217 45796 10251
rect 45744 10208 45796 10217
rect 2504 10004 2556 10056
rect 3884 10004 3936 10056
rect 4160 10004 4212 10056
rect 46296 10047 46348 10056
rect 46296 10013 46305 10047
rect 46305 10013 46339 10047
rect 46339 10013 46348 10047
rect 46296 10004 46348 10013
rect 47400 10047 47452 10056
rect 47400 10013 47409 10047
rect 47409 10013 47443 10047
rect 47443 10013 47452 10047
rect 47400 10004 47452 10013
rect 47584 10047 47636 10056
rect 47584 10013 47593 10047
rect 47593 10013 47627 10047
rect 47627 10013 47636 10047
rect 47584 10004 47636 10013
rect 48044 10047 48096 10056
rect 48044 10013 48053 10047
rect 48053 10013 48087 10047
rect 48087 10013 48096 10047
rect 48044 10004 48096 10013
rect 940 9936 992 9988
rect 2044 9936 2096 9988
rect 756 9868 808 9920
rect 1216 9868 1268 9920
rect 1400 9911 1452 9920
rect 1400 9877 1409 9911
rect 1409 9877 1443 9911
rect 1443 9877 1452 9911
rect 1400 9868 1452 9877
rect 2412 9868 2464 9920
rect 2780 9868 2832 9920
rect 5172 9911 5224 9920
rect 5172 9877 5181 9911
rect 5181 9877 5215 9911
rect 5215 9877 5224 9911
rect 5172 9868 5224 9877
rect 5540 9868 5592 9920
rect 6460 9911 6512 9920
rect 6460 9877 6469 9911
rect 6469 9877 6503 9911
rect 6503 9877 6512 9911
rect 6460 9868 6512 9877
rect 46480 9911 46532 9920
rect 46480 9877 46489 9911
rect 46489 9877 46523 9911
rect 46523 9877 46532 9911
rect 46480 9868 46532 9877
rect 47032 9911 47084 9920
rect 47032 9877 47041 9911
rect 47041 9877 47075 9911
rect 47075 9877 47084 9911
rect 47032 9868 47084 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 1216 9664 1268 9716
rect 2688 9664 2740 9716
rect 6460 9664 6512 9716
rect 47032 9664 47084 9716
rect 1308 9596 1360 9648
rect 6276 9596 6328 9648
rect 7380 9596 7432 9648
rect 8300 9596 8352 9648
rect 46664 9596 46716 9648
rect 46940 9596 46992 9648
rect 46480 9571 46532 9580
rect 46480 9537 46489 9571
rect 46489 9537 46523 9571
rect 46523 9537 46532 9571
rect 46480 9528 46532 9537
rect 1952 9460 2004 9512
rect 8392 9460 8444 9512
rect 27344 9460 27396 9512
rect 45836 9503 45888 9512
rect 45836 9469 45845 9503
rect 45845 9469 45879 9503
rect 45879 9469 45888 9503
rect 45836 9460 45888 9469
rect 46756 9460 46808 9512
rect 48044 9528 48096 9580
rect 48136 9571 48188 9580
rect 48136 9537 48145 9571
rect 48145 9537 48179 9571
rect 48179 9537 48188 9571
rect 48136 9528 48188 9537
rect 4528 9392 4580 9444
rect 5080 9392 5132 9444
rect 7012 9392 7064 9444
rect 45560 9392 45612 9444
rect 1492 9367 1544 9376
rect 1492 9333 1501 9367
rect 1501 9333 1535 9367
rect 1535 9333 1544 9367
rect 1492 9324 1544 9333
rect 1768 9324 1820 9376
rect 2872 9324 2924 9376
rect 3700 9367 3752 9376
rect 3700 9333 3709 9367
rect 3709 9333 3743 9367
rect 3743 9333 3752 9367
rect 3700 9324 3752 9333
rect 4620 9324 4672 9376
rect 4804 9324 4856 9376
rect 5264 9324 5316 9376
rect 6368 9367 6420 9376
rect 6368 9333 6377 9367
rect 6377 9333 6411 9367
rect 6411 9333 6420 9367
rect 6368 9324 6420 9333
rect 6736 9324 6788 9376
rect 47952 9367 48004 9376
rect 47952 9333 47961 9367
rect 47961 9333 47995 9367
rect 47995 9333 48004 9367
rect 47952 9324 48004 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 5724 9120 5776 9172
rect 6736 9120 6788 9172
rect 45836 9120 45888 9172
rect 46388 9163 46440 9172
rect 46388 9129 46397 9163
rect 46397 9129 46431 9163
rect 46431 9129 46440 9163
rect 46388 9120 46440 9129
rect 46756 9120 46808 9172
rect 47400 9120 47452 9172
rect 388 8916 440 8968
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 5632 8916 5684 8968
rect 9680 8916 9732 8968
rect 33140 8916 33192 8968
rect 2320 8780 2372 8832
rect 4988 8848 5040 8900
rect 7288 8848 7340 8900
rect 8116 8848 8168 8900
rect 8944 8891 8996 8900
rect 8944 8857 8953 8891
rect 8953 8857 8987 8891
rect 8987 8857 8996 8891
rect 8944 8848 8996 8857
rect 45652 9052 45704 9104
rect 47216 9052 47268 9104
rect 47400 9027 47452 9036
rect 47400 8993 47409 9027
rect 47409 8993 47443 9027
rect 47443 8993 47452 9027
rect 47400 8984 47452 8993
rect 45192 8916 45244 8968
rect 46204 8959 46256 8968
rect 46204 8925 46213 8959
rect 46213 8925 46247 8959
rect 46247 8925 46256 8959
rect 46204 8916 46256 8925
rect 46296 8916 46348 8968
rect 48320 8984 48372 9036
rect 2964 8823 3016 8832
rect 2964 8789 2973 8823
rect 2973 8789 3007 8823
rect 3007 8789 3016 8823
rect 2964 8780 3016 8789
rect 3608 8780 3660 8832
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 4896 8823 4948 8832
rect 4896 8789 4905 8823
rect 4905 8789 4939 8823
rect 4939 8789 4948 8823
rect 4896 8780 4948 8789
rect 5908 8780 5960 8832
rect 6184 8780 6236 8832
rect 7196 8780 7248 8832
rect 7748 8780 7800 8832
rect 9220 8780 9272 8832
rect 37648 8848 37700 8900
rect 9680 8780 9732 8832
rect 48044 8959 48096 8968
rect 48044 8925 48053 8959
rect 48053 8925 48087 8959
rect 48087 8925 48096 8959
rect 48044 8916 48096 8925
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 5080 8576 5132 8628
rect 8944 8576 8996 8628
rect 44640 8619 44692 8628
rect 4896 8508 4948 8560
rect 4988 8508 5040 8560
rect 5172 8508 5224 8560
rect 37648 8508 37700 8560
rect 44640 8585 44649 8619
rect 44649 8585 44683 8619
rect 44683 8585 44692 8619
rect 44640 8576 44692 8585
rect 46756 8508 46808 8560
rect 48044 8576 48096 8628
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 3332 8440 3384 8492
rect 4712 8440 4764 8492
rect 5080 8440 5132 8492
rect 7840 8372 7892 8424
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 4712 8347 4764 8356
rect 4712 8313 4721 8347
rect 4721 8313 4755 8347
rect 4755 8313 4764 8347
rect 4712 8304 4764 8313
rect 5172 8347 5224 8356
rect 5172 8313 5181 8347
rect 5181 8313 5215 8347
rect 5215 8313 5224 8347
rect 5172 8304 5224 8313
rect 5816 8347 5868 8356
rect 5816 8313 5825 8347
rect 5825 8313 5859 8347
rect 5859 8313 5868 8347
rect 5816 8304 5868 8313
rect 7656 8347 7708 8356
rect 7656 8313 7665 8347
rect 7665 8313 7699 8347
rect 7699 8313 7708 8347
rect 7656 8304 7708 8313
rect 3240 8236 3292 8288
rect 3884 8236 3936 8288
rect 6092 8236 6144 8288
rect 8208 8279 8260 8288
rect 8208 8245 8217 8279
rect 8217 8245 8251 8279
rect 8251 8245 8260 8279
rect 8208 8236 8260 8245
rect 8668 8236 8720 8288
rect 9312 8279 9364 8288
rect 9312 8245 9321 8279
rect 9321 8245 9355 8279
rect 9355 8245 9364 8279
rect 9312 8236 9364 8245
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 10416 8279 10468 8288
rect 10416 8245 10425 8279
rect 10425 8245 10459 8279
rect 10459 8245 10468 8279
rect 10416 8236 10468 8245
rect 46664 8440 46716 8492
rect 46388 8415 46440 8424
rect 46388 8381 46397 8415
rect 46397 8381 46431 8415
rect 46431 8381 46440 8415
rect 46388 8372 46440 8381
rect 45560 8304 45612 8356
rect 45744 8304 45796 8356
rect 47492 8304 47544 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1492 8032 1544 8084
rect 2044 8032 2096 8084
rect 45744 8032 45796 8084
rect 47124 8032 47176 8084
rect 47676 7964 47728 8016
rect 756 7896 808 7948
rect 7564 7896 7616 7948
rect 14832 7896 14884 7948
rect 30380 7896 30432 7948
rect 47216 7896 47268 7948
rect 296 7828 348 7880
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 2504 7828 2556 7880
rect 2780 7828 2832 7880
rect 4068 7828 4120 7880
rect 4528 7828 4580 7880
rect 15384 7828 15436 7880
rect 36636 7828 36688 7880
rect 45652 7871 45704 7880
rect 45652 7837 45661 7871
rect 45661 7837 45695 7871
rect 45695 7837 45704 7871
rect 45652 7828 45704 7837
rect 46112 7828 46164 7880
rect 47400 7871 47452 7880
rect 47400 7837 47409 7871
rect 47409 7837 47443 7871
rect 47443 7837 47452 7871
rect 47400 7828 47452 7837
rect 47584 7871 47636 7880
rect 47584 7837 47593 7871
rect 47593 7837 47627 7871
rect 47627 7837 47636 7871
rect 47584 7828 47636 7837
rect 48044 7871 48096 7880
rect 48044 7837 48053 7871
rect 48053 7837 48087 7871
rect 48087 7837 48096 7871
rect 48044 7828 48096 7837
rect 6552 7760 6604 7812
rect 15844 7760 15896 7812
rect 39304 7760 39356 7812
rect 44548 7760 44600 7812
rect 44640 7760 44692 7812
rect 45468 7760 45520 7812
rect 2044 7692 2096 7744
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 3056 7735 3108 7744
rect 3056 7701 3065 7735
rect 3065 7701 3099 7735
rect 3099 7701 3108 7735
rect 3056 7692 3108 7701
rect 3792 7735 3844 7744
rect 3792 7701 3801 7735
rect 3801 7701 3835 7735
rect 3835 7701 3844 7735
rect 3792 7692 3844 7701
rect 4436 7735 4488 7744
rect 4436 7701 4445 7735
rect 4445 7701 4479 7735
rect 4479 7701 4488 7735
rect 4436 7692 4488 7701
rect 6644 7735 6696 7744
rect 6644 7701 6653 7735
rect 6653 7701 6687 7735
rect 6687 7701 6696 7735
rect 6644 7692 6696 7701
rect 7472 7735 7524 7744
rect 7472 7701 7481 7735
rect 7481 7701 7515 7735
rect 7515 7701 7524 7735
rect 7472 7692 7524 7701
rect 8024 7735 8076 7744
rect 8024 7701 8033 7735
rect 8033 7701 8067 7735
rect 8067 7701 8076 7735
rect 8024 7692 8076 7701
rect 9588 7692 9640 7744
rect 9772 7735 9824 7744
rect 9772 7701 9781 7735
rect 9781 7701 9815 7735
rect 9815 7701 9824 7735
rect 9772 7692 9824 7701
rect 10140 7692 10192 7744
rect 10784 7735 10836 7744
rect 10784 7701 10793 7735
rect 10793 7701 10827 7735
rect 10827 7701 10836 7735
rect 10784 7692 10836 7701
rect 11336 7735 11388 7744
rect 11336 7701 11345 7735
rect 11345 7701 11379 7735
rect 11379 7701 11388 7735
rect 11336 7692 11388 7701
rect 43076 7692 43128 7744
rect 44272 7735 44324 7744
rect 44272 7701 44281 7735
rect 44281 7701 44315 7735
rect 44315 7701 44324 7735
rect 44272 7692 44324 7701
rect 47032 7735 47084 7744
rect 47032 7701 47041 7735
rect 47041 7701 47075 7735
rect 47075 7701 47084 7735
rect 47032 7692 47084 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 2688 7531 2740 7540
rect 2688 7497 2697 7531
rect 2697 7497 2731 7531
rect 2731 7497 2740 7531
rect 2688 7488 2740 7497
rect 6828 7488 6880 7540
rect 11060 7488 11112 7540
rect 47032 7488 47084 7540
rect 2320 7420 2372 7472
rect 44272 7420 44324 7472
rect 2228 7352 2280 7404
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 4712 7352 4764 7404
rect 5264 7352 5316 7404
rect 5632 7352 5684 7404
rect 6000 7352 6052 7404
rect 6368 7352 6420 7404
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 7748 7352 7800 7404
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 9496 7352 9548 7404
rect 10416 7352 10468 7404
rect 12164 7352 12216 7404
rect 43076 7352 43128 7404
rect 43168 7352 43220 7404
rect 44088 7352 44140 7404
rect 45652 7420 45704 7472
rect 45100 7395 45152 7404
rect 45100 7361 45109 7395
rect 45109 7361 45143 7395
rect 45143 7361 45152 7395
rect 45100 7352 45152 7361
rect 45928 7352 45980 7404
rect 47952 7420 48004 7472
rect 1400 7216 1452 7268
rect 8576 7284 8628 7336
rect 16764 7284 16816 7336
rect 46388 7327 46440 7336
rect 46388 7293 46397 7327
rect 46397 7293 46431 7327
rect 46431 7293 46440 7327
rect 46388 7284 46440 7293
rect 46756 7327 46808 7336
rect 46756 7293 46765 7327
rect 46765 7293 46799 7327
rect 46799 7293 46808 7327
rect 46756 7284 46808 7293
rect 2320 7216 2372 7268
rect 10232 7216 10284 7268
rect 11980 7216 12032 7268
rect 12808 7216 12860 7268
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 2780 7148 2832 7200
rect 3976 7148 4028 7200
rect 4988 7191 5040 7200
rect 4988 7157 4997 7191
rect 4997 7157 5031 7191
rect 5031 7157 5040 7191
rect 4988 7148 5040 7157
rect 5632 7191 5684 7200
rect 5632 7157 5641 7191
rect 5641 7157 5675 7191
rect 5675 7157 5684 7191
rect 5632 7148 5684 7157
rect 6368 7191 6420 7200
rect 6368 7157 6377 7191
rect 6377 7157 6411 7191
rect 6411 7157 6420 7191
rect 6368 7148 6420 7157
rect 6920 7148 6972 7200
rect 7932 7148 7984 7200
rect 8300 7148 8352 7200
rect 10692 7148 10744 7200
rect 11704 7148 11756 7200
rect 42800 7191 42852 7200
rect 42800 7157 42809 7191
rect 42809 7157 42843 7191
rect 42843 7157 42852 7191
rect 42800 7148 42852 7157
rect 43168 7148 43220 7200
rect 44088 7216 44140 7268
rect 45100 7216 45152 7268
rect 45192 7216 45244 7268
rect 45468 7216 45520 7268
rect 46020 7148 46072 7200
rect 47860 7148 47912 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3424 6944 3476 6996
rect 572 6876 624 6928
rect 3516 6876 3568 6928
rect 4160 6876 4212 6928
rect 4436 6876 4488 6928
rect 4896 6876 4948 6928
rect 480 6740 532 6792
rect 2136 6808 2188 6860
rect 2596 6808 2648 6860
rect 14372 6944 14424 6996
rect 44456 6919 44508 6928
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 2320 6740 2372 6792
rect 3240 6740 3292 6792
rect 3792 6740 3844 6792
rect 4436 6740 4488 6792
rect 4528 6740 4580 6792
rect 5356 6740 5408 6792
rect 3424 6672 3476 6724
rect 5908 6740 5960 6792
rect 1400 6604 1452 6656
rect 2136 6647 2188 6656
rect 2136 6613 2145 6647
rect 2145 6613 2179 6647
rect 2179 6613 2188 6647
rect 2136 6604 2188 6613
rect 2780 6604 2832 6656
rect 3516 6604 3568 6656
rect 4896 6604 4948 6656
rect 6184 6672 6236 6724
rect 7196 6740 7248 6792
rect 7656 6740 7708 6792
rect 7288 6672 7340 6724
rect 8760 6808 8812 6860
rect 44456 6885 44465 6919
rect 44465 6885 44499 6919
rect 44499 6885 44508 6919
rect 44456 6876 44508 6885
rect 10968 6808 11020 6860
rect 44180 6808 44232 6860
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 8852 6740 8904 6792
rect 9864 6740 9916 6792
rect 10232 6740 10284 6792
rect 10600 6740 10652 6792
rect 11336 6740 11388 6792
rect 11612 6740 11664 6792
rect 13268 6783 13320 6792
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 42800 6740 42852 6792
rect 45376 6808 45428 6860
rect 47216 6808 47268 6860
rect 47400 6851 47452 6860
rect 47400 6817 47409 6851
rect 47409 6817 47443 6851
rect 47443 6817 47452 6851
rect 47400 6808 47452 6817
rect 44824 6740 44876 6792
rect 45652 6783 45704 6792
rect 45652 6749 45661 6783
rect 45661 6749 45695 6783
rect 45695 6749 45704 6783
rect 45652 6740 45704 6749
rect 43260 6715 43312 6724
rect 5540 6604 5592 6656
rect 6460 6604 6512 6656
rect 7104 6604 7156 6656
rect 7932 6604 7984 6656
rect 9036 6647 9088 6656
rect 9036 6613 9045 6647
rect 9045 6613 9079 6647
rect 9079 6613 9088 6647
rect 9036 6604 9088 6613
rect 9128 6604 9180 6656
rect 10416 6604 10468 6656
rect 11520 6647 11572 6656
rect 11520 6613 11529 6647
rect 11529 6613 11563 6647
rect 11563 6613 11572 6647
rect 11520 6604 11572 6613
rect 11796 6604 11848 6656
rect 43260 6681 43269 6715
rect 43269 6681 43303 6715
rect 43303 6681 43312 6715
rect 43260 6672 43312 6681
rect 17040 6604 17092 6656
rect 45744 6604 45796 6656
rect 46296 6604 46348 6656
rect 46756 6740 46808 6792
rect 47676 6740 47728 6792
rect 48044 6783 48096 6792
rect 48044 6749 48053 6783
rect 48053 6749 48087 6783
rect 48087 6749 48096 6783
rect 48044 6740 48096 6749
rect 46940 6715 46992 6724
rect 46940 6681 46949 6715
rect 46949 6681 46983 6715
rect 46983 6681 46992 6715
rect 46940 6672 46992 6681
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2044 6400 2096 6452
rect 2412 6400 2464 6452
rect 2504 6400 2556 6452
rect 1860 6264 1912 6316
rect 1584 6196 1636 6248
rect 1860 6128 1912 6180
rect 3240 6264 3292 6316
rect 4344 6332 4396 6384
rect 4528 6332 4580 6384
rect 8116 6400 8168 6452
rect 11428 6400 11480 6452
rect 23020 6400 23072 6452
rect 44088 6400 44140 6452
rect 44272 6400 44324 6452
rect 45468 6400 45520 6452
rect 45928 6443 45980 6452
rect 45928 6409 45937 6443
rect 45937 6409 45971 6443
rect 45971 6409 45980 6443
rect 45928 6400 45980 6409
rect 4252 6307 4304 6316
rect 4252 6273 4261 6307
rect 4261 6273 4295 6307
rect 4295 6273 4304 6307
rect 4252 6264 4304 6273
rect 4804 6264 4856 6316
rect 4160 6196 4212 6248
rect 8484 6332 8536 6384
rect 5724 6264 5776 6316
rect 7012 6264 7064 6316
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 8392 6264 8444 6316
rect 5448 6196 5500 6248
rect 11060 6332 11112 6384
rect 14004 6375 14056 6384
rect 14004 6341 14013 6375
rect 14013 6341 14047 6375
rect 14047 6341 14056 6375
rect 14004 6332 14056 6341
rect 14556 6375 14608 6384
rect 14556 6341 14565 6375
rect 14565 6341 14599 6375
rect 14599 6341 14608 6375
rect 14556 6332 14608 6341
rect 44456 6332 44508 6384
rect 48044 6400 48096 6452
rect 9680 6264 9732 6316
rect 10140 6264 10192 6316
rect 9404 6196 9456 6248
rect 10784 6264 10836 6316
rect 11244 6264 11296 6316
rect 17224 6264 17276 6316
rect 23664 6264 23716 6316
rect 12256 6239 12308 6248
rect 12256 6205 12265 6239
rect 12265 6205 12299 6239
rect 12299 6205 12308 6239
rect 12256 6196 12308 6205
rect 14372 6196 14424 6248
rect 39304 6196 39356 6248
rect 10968 6128 11020 6180
rect 11336 6128 11388 6180
rect 43168 6196 43220 6248
rect 44548 6264 44600 6316
rect 44916 6264 44968 6316
rect 45192 6307 45244 6316
rect 45192 6273 45201 6307
rect 45201 6273 45235 6307
rect 45235 6273 45244 6307
rect 45192 6264 45244 6273
rect 46848 6307 46900 6316
rect 46848 6273 46857 6307
rect 46857 6273 46891 6307
rect 46891 6273 46900 6307
rect 46848 6264 46900 6273
rect 47492 6264 47544 6316
rect 45560 6196 45612 6248
rect 43260 6128 43312 6180
rect 1124 6060 1176 6112
rect 1584 6060 1636 6112
rect 2412 6060 2464 6112
rect 3792 6060 3844 6112
rect 5080 6060 5132 6112
rect 5724 6060 5776 6112
rect 6184 6060 6236 6112
rect 6276 6060 6328 6112
rect 7012 6060 7064 6112
rect 7564 6060 7616 6112
rect 8208 6060 8260 6112
rect 8392 6060 8444 6112
rect 9036 6103 9088 6112
rect 9036 6069 9045 6103
rect 9045 6069 9079 6103
rect 9079 6069 9088 6103
rect 9036 6060 9088 6069
rect 10324 6103 10376 6112
rect 10324 6069 10333 6103
rect 10333 6069 10367 6103
rect 10367 6069 10376 6103
rect 10324 6060 10376 6069
rect 12532 6060 12584 6112
rect 13084 6060 13136 6112
rect 15200 6103 15252 6112
rect 15200 6069 15209 6103
rect 15209 6069 15243 6103
rect 15243 6069 15252 6103
rect 15200 6060 15252 6069
rect 44548 6103 44600 6112
rect 44548 6069 44557 6103
rect 44557 6069 44591 6103
rect 44591 6069 44600 6103
rect 44548 6060 44600 6069
rect 45100 6103 45152 6112
rect 45100 6069 45109 6103
rect 45109 6069 45143 6103
rect 45143 6069 45152 6103
rect 45100 6060 45152 6069
rect 47400 6128 47452 6180
rect 47584 6060 47636 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1032 5856 1084 5908
rect 2136 5856 2188 5908
rect 7380 5899 7432 5908
rect 1124 5788 1176 5840
rect 1492 5652 1544 5704
rect 4160 5763 4212 5772
rect 4160 5729 4169 5763
rect 4169 5729 4203 5763
rect 4203 5729 4212 5763
rect 4160 5720 4212 5729
rect 5448 5720 5500 5772
rect 6736 5788 6788 5840
rect 7380 5865 7389 5899
rect 7389 5865 7423 5899
rect 7423 5865 7432 5899
rect 7380 5856 7432 5865
rect 8116 5856 8168 5908
rect 8208 5856 8260 5908
rect 9312 5856 9364 5908
rect 10232 5856 10284 5908
rect 12256 5856 12308 5908
rect 15292 5856 15344 5908
rect 15844 5899 15896 5908
rect 15844 5865 15853 5899
rect 15853 5865 15887 5899
rect 15887 5865 15896 5899
rect 15844 5856 15896 5865
rect 45008 5788 45060 5840
rect 45192 5788 45244 5840
rect 47400 5856 47452 5908
rect 46756 5788 46808 5840
rect 47216 5831 47268 5840
rect 47216 5797 47225 5831
rect 47225 5797 47259 5831
rect 47259 5797 47268 5831
rect 47216 5788 47268 5797
rect 47308 5788 47360 5840
rect 2596 5652 2648 5704
rect 4252 5652 4304 5704
rect 5724 5652 5776 5704
rect 6184 5652 6236 5704
rect 2136 5584 2188 5636
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 2964 5559 3016 5568
rect 2964 5525 2973 5559
rect 2973 5525 3007 5559
rect 3007 5525 3016 5559
rect 2964 5516 3016 5525
rect 3240 5584 3292 5636
rect 5448 5584 5500 5636
rect 6828 5652 6880 5704
rect 7380 5652 7432 5704
rect 8116 5652 8168 5704
rect 10968 5720 11020 5772
rect 12440 5763 12492 5772
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 10048 5652 10100 5704
rect 10232 5652 10284 5704
rect 12440 5729 12449 5763
rect 12449 5729 12483 5763
rect 12483 5729 12492 5763
rect 12440 5720 12492 5729
rect 14280 5720 14332 5772
rect 15200 5720 15252 5772
rect 44456 5720 44508 5772
rect 44548 5720 44600 5772
rect 11704 5695 11756 5704
rect 11704 5661 11713 5695
rect 11713 5661 11747 5695
rect 11747 5661 11756 5695
rect 11704 5652 11756 5661
rect 11980 5652 12032 5704
rect 17224 5652 17276 5704
rect 43628 5695 43680 5704
rect 43628 5661 43637 5695
rect 43637 5661 43671 5695
rect 43671 5661 43680 5695
rect 43628 5652 43680 5661
rect 44088 5652 44140 5704
rect 45836 5652 45888 5704
rect 47400 5695 47452 5704
rect 47400 5661 47409 5695
rect 47409 5661 47443 5695
rect 47443 5661 47452 5695
rect 47400 5652 47452 5661
rect 48044 5695 48096 5704
rect 48044 5661 48053 5695
rect 48053 5661 48087 5695
rect 48087 5661 48096 5695
rect 48044 5652 48096 5661
rect 4160 5516 4212 5568
rect 4620 5516 4672 5568
rect 4804 5516 4856 5568
rect 5724 5516 5776 5568
rect 8116 5516 8168 5568
rect 8300 5516 8352 5568
rect 10600 5584 10652 5636
rect 11244 5627 11296 5636
rect 11244 5593 11253 5627
rect 11253 5593 11287 5627
rect 11287 5593 11296 5627
rect 11244 5584 11296 5593
rect 14372 5584 14424 5636
rect 47492 5584 47544 5636
rect 12256 5516 12308 5568
rect 12900 5559 12952 5568
rect 12900 5525 12909 5559
rect 12909 5525 12943 5559
rect 12943 5525 12952 5559
rect 12900 5516 12952 5525
rect 12992 5516 13044 5568
rect 13636 5516 13688 5568
rect 15384 5516 15436 5568
rect 42064 5559 42116 5568
rect 42064 5525 42073 5559
rect 42073 5525 42107 5559
rect 42107 5525 42116 5559
rect 42064 5516 42116 5525
rect 42616 5559 42668 5568
rect 42616 5525 42625 5559
rect 42625 5525 42659 5559
rect 42659 5525 42668 5559
rect 42616 5516 42668 5525
rect 44272 5516 44324 5568
rect 45192 5516 45244 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1308 5244 1360 5296
rect 3240 5312 3292 5364
rect 3608 5312 3660 5364
rect 3700 5287 3752 5296
rect 3700 5253 3709 5287
rect 3709 5253 3743 5287
rect 3743 5253 3752 5287
rect 3700 5244 3752 5253
rect 4160 5244 4212 5296
rect 4528 5244 4580 5296
rect 1216 5176 1268 5228
rect 2136 5176 2188 5228
rect 2872 5176 2924 5228
rect 6920 5312 6972 5364
rect 7288 5244 7340 5296
rect 3700 5108 3752 5160
rect 4068 5108 4120 5160
rect 6184 5108 6236 5160
rect 7656 5312 7708 5364
rect 8484 5312 8536 5364
rect 9220 5312 9272 5364
rect 10140 5312 10192 5364
rect 10876 5312 10928 5364
rect 10232 5287 10284 5296
rect 7656 5176 7708 5228
rect 8024 5176 8076 5228
rect 204 4972 256 5024
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 5356 4972 5408 5024
rect 6828 5015 6880 5024
rect 6828 4981 6837 5015
rect 6837 4981 6871 5015
rect 6871 4981 6880 5015
rect 6828 4972 6880 4981
rect 7380 4972 7432 5024
rect 8024 5040 8076 5092
rect 10232 5253 10241 5287
rect 10241 5253 10275 5287
rect 10275 5253 10284 5287
rect 10232 5244 10284 5253
rect 10600 5244 10652 5296
rect 11336 5244 11388 5296
rect 8300 5108 8352 5160
rect 8484 5108 8536 5160
rect 14556 5244 14608 5296
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 15660 5312 15712 5364
rect 16120 5312 16172 5364
rect 44640 5312 44692 5364
rect 42616 5244 42668 5296
rect 44088 5244 44140 5296
rect 44180 5244 44232 5296
rect 13084 5176 13136 5185
rect 25228 5176 25280 5228
rect 43260 5219 43312 5228
rect 43260 5185 43269 5219
rect 43269 5185 43303 5219
rect 43303 5185 43312 5219
rect 43260 5176 43312 5185
rect 10600 5108 10652 5160
rect 11060 5108 11112 5160
rect 21364 5108 21416 5160
rect 44456 5176 44508 5228
rect 45100 5151 45152 5160
rect 45100 5117 45109 5151
rect 45109 5117 45143 5151
rect 45143 5117 45152 5151
rect 45100 5108 45152 5117
rect 8300 4972 8352 5024
rect 8484 4972 8536 5024
rect 8944 4972 8996 5024
rect 10508 5040 10560 5092
rect 9496 4972 9548 5024
rect 11336 4972 11388 5024
rect 47124 5176 47176 5228
rect 45376 5108 45428 5160
rect 45836 5108 45888 5160
rect 11888 4972 11940 5024
rect 12348 4972 12400 5024
rect 13176 4972 13228 5024
rect 14096 5015 14148 5024
rect 14096 4981 14105 5015
rect 14105 4981 14139 5015
rect 14139 4981 14148 5015
rect 14096 4972 14148 4981
rect 29092 5015 29144 5024
rect 29092 4981 29101 5015
rect 29101 4981 29135 5015
rect 29135 4981 29144 5015
rect 29092 4972 29144 4981
rect 30012 5015 30064 5024
rect 30012 4981 30021 5015
rect 30021 4981 30055 5015
rect 30055 4981 30064 5015
rect 30012 4972 30064 4981
rect 41328 5015 41380 5024
rect 41328 4981 41337 5015
rect 41337 4981 41371 5015
rect 41371 4981 41380 5015
rect 41328 4972 41380 4981
rect 45652 4972 45704 5024
rect 46296 4972 46348 5024
rect 46664 4972 46716 5024
rect 47032 4972 47084 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2320 4768 2372 4820
rect 2596 4768 2648 4820
rect 2872 4768 2924 4820
rect 664 4700 716 4752
rect 8484 4768 8536 4820
rect 8944 4811 8996 4820
rect 1032 4564 1084 4616
rect 1768 4564 1820 4616
rect 4068 4632 4120 4684
rect 8208 4700 8260 4752
rect 8576 4700 8628 4752
rect 8944 4777 8953 4811
rect 8953 4777 8987 4811
rect 8987 4777 8996 4811
rect 8944 4768 8996 4777
rect 9036 4768 9088 4820
rect 8852 4700 8904 4752
rect 4344 4564 4396 4616
rect 5816 4564 5868 4616
rect 6092 4564 6144 4616
rect 2044 4496 2096 4548
rect 3240 4496 3292 4548
rect 4436 4496 4488 4548
rect 8024 4632 8076 4684
rect 8300 4632 8352 4684
rect 9220 4700 9272 4752
rect 6920 4564 6972 4616
rect 7840 4564 7892 4616
rect 8852 4564 8904 4616
rect 9680 4768 9732 4820
rect 9496 4700 9548 4752
rect 17132 4768 17184 4820
rect 46388 4768 46440 4820
rect 9772 4564 9824 4616
rect 11428 4700 11480 4752
rect 11612 4700 11664 4752
rect 14372 4700 14424 4752
rect 11060 4675 11112 4684
rect 11060 4641 11069 4675
rect 11069 4641 11103 4675
rect 11103 4641 11112 4675
rect 11060 4632 11112 4641
rect 11244 4632 11296 4684
rect 11796 4632 11848 4684
rect 10784 4607 10836 4616
rect 10784 4573 10793 4607
rect 10793 4573 10827 4607
rect 10827 4573 10836 4607
rect 12808 4632 12860 4684
rect 16948 4675 17000 4684
rect 16948 4641 16957 4675
rect 16957 4641 16991 4675
rect 16991 4641 17000 4675
rect 16948 4632 17000 4641
rect 10784 4564 10836 4573
rect 10968 4496 11020 4548
rect 12440 4607 12492 4616
rect 12440 4573 12449 4607
rect 12449 4573 12483 4607
rect 12483 4573 12492 4607
rect 12440 4564 12492 4573
rect 13820 4564 13872 4616
rect 15200 4564 15252 4616
rect 29092 4564 29144 4616
rect 29920 4564 29972 4616
rect 30012 4564 30064 4616
rect 13636 4496 13688 4548
rect 37924 4564 37976 4616
rect 42064 4564 42116 4616
rect 42524 4607 42576 4616
rect 42524 4573 42533 4607
rect 42533 4573 42567 4607
rect 42567 4573 42576 4607
rect 42524 4564 42576 4573
rect 45376 4700 45428 4752
rect 45744 4700 45796 4752
rect 45100 4632 45152 4684
rect 45836 4632 45888 4684
rect 47400 4675 47452 4684
rect 47400 4641 47409 4675
rect 47409 4641 47443 4675
rect 47443 4641 47452 4675
rect 47400 4632 47452 4641
rect 45008 4607 45060 4616
rect 45008 4573 45017 4607
rect 45017 4573 45051 4607
rect 45051 4573 45060 4607
rect 45008 4564 45060 4573
rect 45652 4607 45704 4616
rect 45652 4573 45661 4607
rect 45661 4573 45695 4607
rect 45695 4573 45704 4607
rect 45652 4564 45704 4573
rect 7840 4428 7892 4480
rect 9036 4428 9088 4480
rect 9588 4428 9640 4480
rect 9680 4428 9732 4480
rect 10600 4428 10652 4480
rect 11060 4428 11112 4480
rect 12164 4428 12216 4480
rect 16304 4471 16356 4480
rect 16304 4437 16313 4471
rect 16313 4437 16347 4471
rect 16347 4437 16356 4471
rect 44180 4539 44232 4548
rect 44180 4505 44189 4539
rect 44189 4505 44223 4539
rect 44223 4505 44232 4539
rect 44180 4496 44232 4505
rect 28816 4471 28868 4480
rect 16304 4428 16356 4437
rect 28816 4437 28825 4471
rect 28825 4437 28859 4471
rect 28859 4437 28868 4471
rect 28816 4428 28868 4437
rect 29460 4428 29512 4480
rect 30564 4428 30616 4480
rect 30748 4471 30800 4480
rect 30748 4437 30757 4471
rect 30757 4437 30791 4471
rect 30791 4437 30800 4471
rect 30748 4428 30800 4437
rect 31392 4471 31444 4480
rect 31392 4437 31401 4471
rect 31401 4437 31435 4471
rect 31435 4437 31444 4471
rect 31392 4428 31444 4437
rect 40408 4471 40460 4480
rect 40408 4437 40417 4471
rect 40417 4437 40451 4471
rect 40451 4437 40460 4471
rect 40408 4428 40460 4437
rect 40868 4471 40920 4480
rect 40868 4437 40877 4471
rect 40877 4437 40911 4471
rect 40911 4437 40920 4471
rect 40868 4428 40920 4437
rect 41512 4471 41564 4480
rect 41512 4437 41521 4471
rect 41521 4437 41555 4471
rect 41555 4437 41564 4471
rect 41512 4428 41564 4437
rect 44640 4496 44692 4548
rect 46572 4564 46624 4616
rect 47768 4564 47820 4616
rect 48044 4607 48096 4616
rect 48044 4573 48053 4607
rect 48053 4573 48087 4607
rect 48087 4573 48096 4607
rect 48044 4564 48096 4573
rect 46940 4539 46992 4548
rect 46940 4505 46949 4539
rect 46949 4505 46983 4539
rect 46983 4505 46992 4539
rect 46940 4496 46992 4505
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 1860 4224 1912 4276
rect 1952 4199 2004 4208
rect 1952 4165 1961 4199
rect 1961 4165 1995 4199
rect 1995 4165 2004 4199
rect 1952 4156 2004 4165
rect 756 4088 808 4140
rect 1492 4088 1544 4140
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 3056 4224 3108 4276
rect 4436 4224 4488 4276
rect 5908 4224 5960 4276
rect 3700 4156 3752 4208
rect 3240 4088 3292 4140
rect 4344 4156 4396 4208
rect 6552 4156 6604 4208
rect 8484 4224 8536 4276
rect 8852 4224 8904 4276
rect 9588 4224 9640 4276
rect 9772 4224 9824 4276
rect 4068 4088 4120 4140
rect 4528 4131 4580 4140
rect 4528 4097 4562 4131
rect 4562 4097 4580 4131
rect 4528 4088 4580 4097
rect 5908 4088 5960 4140
rect 1492 3952 1544 4004
rect 2964 3952 3016 4004
rect 1124 3884 1176 3936
rect 3240 3927 3292 3936
rect 3240 3893 3249 3927
rect 3249 3893 3283 3927
rect 3283 3893 3292 3927
rect 3240 3884 3292 3893
rect 6552 4020 6604 4072
rect 7012 4156 7064 4208
rect 8116 4088 8168 4140
rect 8484 4088 8536 4140
rect 8392 4020 8444 4072
rect 9404 4088 9456 4140
rect 9588 4088 9640 4140
rect 10600 4224 10652 4276
rect 13084 4224 13136 4276
rect 41512 4224 41564 4276
rect 47768 4224 47820 4276
rect 10692 4156 10744 4208
rect 14004 4156 14056 4208
rect 9680 4063 9732 4072
rect 9680 4029 9689 4063
rect 9689 4029 9723 4063
rect 9723 4029 9732 4063
rect 9680 4020 9732 4029
rect 9956 4020 10008 4072
rect 10692 4063 10744 4072
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 10692 4020 10744 4029
rect 16948 4088 17000 4140
rect 20168 4088 20220 4140
rect 20352 4088 20404 4140
rect 30748 4131 30800 4140
rect 30748 4097 30757 4131
rect 30757 4097 30791 4131
rect 30791 4097 30800 4131
rect 31392 4131 31444 4140
rect 30748 4088 30800 4097
rect 31392 4097 31401 4131
rect 31401 4097 31435 4131
rect 31435 4097 31444 4131
rect 31392 4088 31444 4097
rect 41328 4156 41380 4208
rect 41696 4131 41748 4140
rect 41696 4097 41705 4131
rect 41705 4097 41739 4131
rect 41739 4097 41748 4131
rect 41696 4088 41748 4097
rect 45836 4156 45888 4208
rect 45192 4131 45244 4140
rect 45192 4097 45201 4131
rect 45201 4097 45235 4131
rect 45235 4097 45244 4131
rect 45192 4088 45244 4097
rect 45560 4131 45612 4140
rect 45560 4097 45569 4131
rect 45569 4097 45603 4131
rect 45603 4097 45612 4131
rect 45560 4088 45612 4097
rect 45652 4088 45704 4140
rect 48688 4088 48740 4140
rect 16304 4020 16356 4072
rect 17040 4020 17092 4072
rect 45100 4063 45152 4072
rect 45100 4029 45109 4063
rect 45109 4029 45143 4063
rect 45143 4029 45152 4063
rect 45100 4020 45152 4029
rect 45376 4020 45428 4072
rect 9404 3952 9456 4004
rect 7840 3884 7892 3936
rect 8392 3884 8444 3936
rect 9496 3884 9548 3936
rect 10324 3884 10376 3936
rect 10508 3884 10560 3936
rect 10968 3952 11020 4004
rect 11796 3884 11848 3936
rect 12716 3884 12768 3936
rect 13452 3884 13504 3936
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 14556 3952 14608 4004
rect 17132 3952 17184 4004
rect 22284 3952 22336 4004
rect 29736 3952 29788 4004
rect 30748 3952 30800 4004
rect 16396 3884 16448 3936
rect 17224 3884 17276 3936
rect 18420 3927 18472 3936
rect 18420 3893 18429 3927
rect 18429 3893 18463 3927
rect 18463 3893 18472 3927
rect 18420 3884 18472 3893
rect 27988 3927 28040 3936
rect 27988 3893 27997 3927
rect 27997 3893 28031 3927
rect 28031 3893 28040 3927
rect 27988 3884 28040 3893
rect 28632 3927 28684 3936
rect 28632 3893 28641 3927
rect 28641 3893 28675 3927
rect 28675 3893 28684 3927
rect 28632 3884 28684 3893
rect 28908 3884 28960 3936
rect 30104 3927 30156 3936
rect 30104 3893 30113 3927
rect 30113 3893 30147 3927
rect 30147 3893 30156 3927
rect 30104 3884 30156 3893
rect 30196 3884 30248 3936
rect 30656 3884 30708 3936
rect 45560 3952 45612 4004
rect 31208 3927 31260 3936
rect 31208 3893 31217 3927
rect 31217 3893 31251 3927
rect 31251 3893 31260 3927
rect 31208 3884 31260 3893
rect 40684 3927 40736 3936
rect 40684 3893 40693 3927
rect 40693 3893 40727 3927
rect 40727 3893 40736 3927
rect 40684 3884 40736 3893
rect 41880 3927 41932 3936
rect 41880 3893 41889 3927
rect 41889 3893 41923 3927
rect 41923 3893 41932 3927
rect 41880 3884 41932 3893
rect 42800 3927 42852 3936
rect 42800 3893 42809 3927
rect 42809 3893 42843 3927
rect 42843 3893 42852 3927
rect 42800 3884 42852 3893
rect 47216 4020 47268 4072
rect 46020 3952 46072 4004
rect 45744 3884 45796 3936
rect 46388 3884 46440 3936
rect 48136 3952 48188 4004
rect 49792 3884 49844 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 848 3680 900 3732
rect 3148 3680 3200 3732
rect 3240 3680 3292 3732
rect 1952 3612 2004 3664
rect 2872 3612 2924 3664
rect 664 3476 716 3528
rect 2136 3519 2188 3528
rect 2136 3485 2145 3519
rect 2145 3485 2179 3519
rect 2179 3485 2188 3519
rect 2136 3476 2188 3485
rect 3700 3612 3752 3664
rect 3700 3476 3752 3528
rect 4896 3680 4948 3732
rect 6184 3680 6236 3732
rect 6828 3680 6880 3732
rect 8300 3680 8352 3732
rect 9312 3680 9364 3732
rect 8392 3612 8444 3664
rect 8760 3612 8812 3664
rect 8852 3612 8904 3664
rect 11796 3680 11848 3732
rect 11980 3680 12032 3732
rect 12164 3680 12216 3732
rect 14372 3680 14424 3732
rect 14648 3680 14700 3732
rect 40684 3680 40736 3732
rect 44916 3680 44968 3732
rect 9864 3612 9916 3664
rect 10416 3612 10468 3664
rect 14832 3612 14884 3664
rect 23756 3655 23808 3664
rect 23756 3621 23765 3655
rect 23765 3621 23799 3655
rect 23799 3621 23808 3655
rect 23756 3612 23808 3621
rect 29552 3612 29604 3664
rect 30288 3612 30340 3664
rect 31392 3612 31444 3664
rect 39304 3612 39356 3664
rect 2964 3408 3016 3460
rect 3148 3340 3200 3392
rect 4344 3476 4396 3528
rect 4988 3476 5040 3528
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 4620 3408 4672 3460
rect 5356 3408 5408 3460
rect 4528 3340 4580 3392
rect 6644 3544 6696 3596
rect 6828 3544 6880 3596
rect 7932 3587 7984 3596
rect 7932 3553 7941 3587
rect 7941 3553 7975 3587
rect 7975 3553 7984 3587
rect 7932 3544 7984 3553
rect 9036 3544 9088 3596
rect 7104 3476 7156 3528
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 7472 3408 7524 3460
rect 8300 3476 8352 3528
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 9956 3544 10008 3596
rect 10508 3544 10560 3596
rect 9772 3476 9824 3528
rect 11428 3544 11480 3596
rect 11244 3476 11296 3528
rect 11060 3451 11112 3460
rect 11060 3417 11069 3451
rect 11069 3417 11103 3451
rect 11103 3417 11112 3451
rect 11060 3408 11112 3417
rect 12624 3544 12676 3596
rect 14280 3544 14332 3596
rect 13268 3476 13320 3528
rect 16028 3544 16080 3596
rect 14740 3476 14792 3528
rect 15016 3476 15068 3528
rect 16948 3476 17000 3528
rect 17868 3476 17920 3528
rect 19064 3476 19116 3528
rect 19432 3476 19484 3528
rect 20536 3519 20588 3528
rect 20536 3485 20545 3519
rect 20545 3485 20579 3519
rect 20579 3485 20588 3519
rect 20536 3476 20588 3485
rect 20812 3476 20864 3528
rect 21456 3476 21508 3528
rect 22376 3476 22428 3528
rect 23296 3519 23348 3528
rect 23296 3485 23305 3519
rect 23305 3485 23339 3519
rect 23339 3485 23348 3519
rect 23296 3476 23348 3485
rect 24124 3476 24176 3528
rect 25044 3519 25096 3528
rect 25044 3485 25053 3519
rect 25053 3485 25087 3519
rect 25087 3485 25096 3519
rect 25044 3476 25096 3485
rect 25964 3519 26016 3528
rect 25964 3485 25973 3519
rect 25973 3485 26007 3519
rect 26007 3485 26016 3519
rect 25964 3476 26016 3485
rect 26240 3476 26292 3528
rect 27436 3476 27488 3528
rect 28080 3476 28132 3528
rect 28356 3476 28408 3528
rect 29276 3476 29328 3528
rect 30472 3476 30524 3528
rect 31024 3476 31076 3528
rect 31944 3476 31996 3528
rect 33140 3476 33192 3528
rect 34612 3476 34664 3528
rect 35348 3519 35400 3528
rect 35348 3485 35357 3519
rect 35357 3485 35391 3519
rect 35391 3485 35400 3519
rect 35348 3476 35400 3485
rect 35808 3476 35860 3528
rect 36176 3476 36228 3528
rect 37004 3476 37056 3528
rect 38200 3519 38252 3528
rect 38200 3485 38209 3519
rect 38209 3485 38243 3519
rect 38243 3485 38252 3519
rect 38200 3476 38252 3485
rect 39120 3519 39172 3528
rect 39120 3485 39129 3519
rect 39129 3485 39163 3519
rect 39163 3485 39172 3519
rect 39120 3476 39172 3485
rect 40316 3519 40368 3528
rect 40316 3485 40325 3519
rect 40325 3485 40359 3519
rect 40359 3485 40368 3519
rect 40316 3476 40368 3485
rect 41236 3519 41288 3528
rect 41236 3485 41245 3519
rect 41245 3485 41279 3519
rect 41279 3485 41288 3519
rect 41236 3476 41288 3485
rect 35256 3408 35308 3460
rect 35900 3408 35952 3460
rect 40408 3408 40460 3460
rect 8024 3340 8076 3392
rect 9496 3340 9548 3392
rect 9772 3340 9824 3392
rect 10140 3340 10192 3392
rect 10508 3340 10560 3392
rect 24216 3340 24268 3392
rect 31116 3340 31168 3392
rect 36084 3340 36136 3392
rect 42156 3519 42208 3528
rect 42156 3485 42165 3519
rect 42165 3485 42199 3519
rect 42199 3485 42208 3519
rect 42156 3476 42208 3485
rect 43076 3476 43128 3528
rect 45008 3476 45060 3528
rect 45284 3519 45336 3528
rect 45284 3485 45288 3519
rect 45288 3485 45322 3519
rect 45322 3485 45336 3519
rect 45284 3476 45336 3485
rect 45468 3680 45520 3732
rect 45836 3680 45888 3732
rect 47492 3680 47544 3732
rect 49148 3612 49200 3664
rect 48964 3544 49016 3596
rect 45652 3519 45704 3528
rect 45652 3485 45661 3519
rect 45661 3485 45695 3519
rect 45695 3485 45704 3519
rect 45652 3476 45704 3485
rect 45836 3408 45888 3460
rect 45376 3340 45428 3392
rect 45560 3340 45612 3392
rect 49516 3340 49568 3392
rect 940 3272 992 3324
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 1400 3136 1452 3188
rect 2780 3136 2832 3188
rect 2872 3136 2924 3188
rect 3148 3136 3200 3188
rect 3700 3179 3752 3188
rect 3700 3145 3709 3179
rect 3709 3145 3743 3179
rect 3743 3145 3752 3179
rect 3700 3136 3752 3145
rect 3884 3136 3936 3188
rect 4436 3136 4488 3188
rect 6736 3136 6788 3188
rect 7288 3179 7340 3188
rect 7288 3145 7297 3179
rect 7297 3145 7331 3179
rect 7331 3145 7340 3179
rect 7288 3136 7340 3145
rect 9588 3136 9640 3188
rect 9680 3136 9732 3188
rect 10048 3136 10100 3188
rect 12348 3136 12400 3188
rect 1768 3068 1820 3120
rect 2136 3068 2188 3120
rect 2228 3068 2280 3120
rect 112 3000 164 3052
rect 1676 3000 1728 3052
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 4896 3068 4948 3120
rect 6368 3068 6420 3120
rect 2872 3000 2924 3009
rect 4252 3000 4304 3052
rect 5540 3043 5592 3052
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 5908 3000 5960 3052
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 1768 2932 1820 2984
rect 572 2864 624 2916
rect 3424 2932 3476 2984
rect 4160 2932 4212 2984
rect 4344 2932 4396 2984
rect 4896 2932 4948 2984
rect 5264 2932 5316 2984
rect 6460 2932 6512 2984
rect 6920 2932 6972 2984
rect 3700 2864 3752 2916
rect 3884 2864 3936 2916
rect 5172 2864 5224 2916
rect 2044 2796 2096 2848
rect 2688 2839 2740 2848
rect 2688 2805 2697 2839
rect 2697 2805 2731 2839
rect 2731 2805 2740 2839
rect 2688 2796 2740 2805
rect 3976 2839 4028 2848
rect 3976 2805 3985 2839
rect 3985 2805 4019 2839
rect 4019 2805 4028 2839
rect 3976 2796 4028 2805
rect 5632 2839 5684 2848
rect 5632 2805 5641 2839
rect 5641 2805 5675 2839
rect 5675 2805 5684 2839
rect 5632 2796 5684 2805
rect 6368 2839 6420 2848
rect 6368 2805 6377 2839
rect 6377 2805 6411 2839
rect 6411 2805 6420 2839
rect 6368 2796 6420 2805
rect 6460 2796 6512 2848
rect 8208 3000 8260 3052
rect 9036 3000 9088 3052
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 10048 3000 10100 3052
rect 7472 2932 7524 2984
rect 8116 2932 8168 2984
rect 8392 2932 8444 2984
rect 10140 2975 10192 2984
rect 10140 2941 10149 2975
rect 10149 2941 10183 2975
rect 10183 2941 10192 2975
rect 10140 2932 10192 2941
rect 7104 2864 7156 2916
rect 7564 2864 7616 2916
rect 8208 2864 8260 2916
rect 10600 3000 10652 3052
rect 10784 3000 10836 3052
rect 10876 3000 10928 3052
rect 11428 3000 11480 3052
rect 12348 3000 12400 3052
rect 12992 3136 13044 3188
rect 13268 3136 13320 3188
rect 14648 3136 14700 3188
rect 20352 3179 20404 3188
rect 20352 3145 20361 3179
rect 20361 3145 20395 3179
rect 20395 3145 20404 3179
rect 20352 3136 20404 3145
rect 24216 3179 24268 3188
rect 24216 3145 24225 3179
rect 24225 3145 24259 3179
rect 24259 3145 24268 3179
rect 24216 3136 24268 3145
rect 28540 3179 28592 3188
rect 28540 3145 28549 3179
rect 28549 3145 28583 3179
rect 28583 3145 28592 3179
rect 28540 3136 28592 3145
rect 30196 3136 30248 3188
rect 30564 3136 30616 3188
rect 31116 3136 31168 3188
rect 35900 3136 35952 3188
rect 36084 3179 36136 3188
rect 36084 3145 36093 3179
rect 36093 3145 36127 3179
rect 36127 3145 36136 3179
rect 36084 3136 36136 3145
rect 14464 3068 14516 3120
rect 18512 3111 18564 3120
rect 18512 3077 18521 3111
rect 18521 3077 18555 3111
rect 18555 3077 18564 3111
rect 18512 3068 18564 3077
rect 20168 3068 20220 3120
rect 22284 3111 22336 3120
rect 22284 3077 22293 3111
rect 22293 3077 22327 3111
rect 22327 3077 22336 3111
rect 22284 3068 22336 3077
rect 13268 3000 13320 3052
rect 15844 3000 15896 3052
rect 23756 3000 23808 3052
rect 27988 3068 28040 3120
rect 29828 3111 29880 3120
rect 29828 3077 29837 3111
rect 29837 3077 29871 3111
rect 29871 3077 29880 3111
rect 29828 3068 29880 3077
rect 35256 3068 35308 3120
rect 35716 3068 35768 3120
rect 11796 2975 11848 2984
rect 7012 2839 7064 2848
rect 7012 2805 7021 2839
rect 7021 2805 7055 2839
rect 7055 2805 7064 2839
rect 7012 2796 7064 2805
rect 9128 2796 9180 2848
rect 9312 2796 9364 2848
rect 9680 2796 9732 2848
rect 9956 2796 10008 2848
rect 11796 2941 11805 2975
rect 11805 2941 11839 2975
rect 11839 2941 11848 2975
rect 11796 2932 11848 2941
rect 14188 2932 14240 2984
rect 24492 2932 24544 2984
rect 11520 2864 11572 2916
rect 14740 2907 14792 2916
rect 14740 2873 14749 2907
rect 14749 2873 14783 2907
rect 14783 2873 14792 2907
rect 14740 2864 14792 2873
rect 10876 2796 10928 2848
rect 11244 2796 11296 2848
rect 12440 2796 12492 2848
rect 14280 2796 14332 2848
rect 14924 2796 14976 2848
rect 15752 2864 15804 2916
rect 18144 2864 18196 2916
rect 19984 2864 20036 2916
rect 21732 2864 21784 2916
rect 23572 2864 23624 2916
rect 25320 2864 25372 2916
rect 28816 2932 28868 2984
rect 30380 3000 30432 3052
rect 40684 3000 40736 3052
rect 47124 3136 47176 3188
rect 47308 3136 47360 3188
rect 48412 3136 48464 3188
rect 41696 3068 41748 3120
rect 45560 3068 45612 3120
rect 45468 3000 45520 3052
rect 49056 3068 49108 3120
rect 30656 2932 30708 2984
rect 31208 2932 31260 2984
rect 33416 2932 33468 2984
rect 37924 2932 37976 2984
rect 44180 2932 44232 2984
rect 40868 2864 40920 2916
rect 26516 2796 26568 2848
rect 27160 2796 27212 2848
rect 31392 2796 31444 2848
rect 32220 2796 32272 2848
rect 32864 2796 32916 2848
rect 34060 2796 34112 2848
rect 36452 2796 36504 2848
rect 37372 2796 37424 2848
rect 38568 2796 38620 2848
rect 39396 2796 39448 2848
rect 40040 2796 40092 2848
rect 40684 2796 40736 2848
rect 41880 2796 41932 2848
rect 42708 2796 42760 2848
rect 43352 2796 43404 2848
rect 43904 2796 43956 2848
rect 44548 2796 44600 2848
rect 49608 2864 49660 2916
rect 49332 2796 49384 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 1492 2592 1544 2644
rect 2504 2592 2556 2644
rect 2688 2592 2740 2644
rect 2872 2592 2924 2644
rect 3148 2635 3200 2644
rect 3148 2601 3157 2635
rect 3157 2601 3191 2635
rect 3191 2601 3200 2635
rect 3148 2592 3200 2601
rect 6736 2592 6788 2644
rect 7564 2592 7616 2644
rect 7932 2592 7984 2644
rect 8484 2524 8536 2576
rect 9404 2524 9456 2576
rect 10140 2592 10192 2644
rect 2044 2456 2096 2508
rect 2504 2456 2556 2508
rect 3056 2499 3108 2508
rect 3056 2465 3065 2499
rect 3065 2465 3099 2499
rect 3099 2465 3108 2499
rect 3056 2456 3108 2465
rect 7288 2456 7340 2508
rect 9680 2456 9732 2508
rect 9864 2456 9916 2508
rect 10324 2456 10376 2508
rect 11060 2524 11112 2576
rect 11980 2524 12032 2576
rect 29184 2592 29236 2644
rect 42524 2592 42576 2644
rect 46848 2592 46900 2644
rect 480 2388 532 2440
rect 848 2388 900 2440
rect 2320 2388 2372 2440
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 4344 2388 4396 2440
rect 6368 2388 6420 2440
rect 4160 2320 4212 2372
rect 4712 2320 4764 2372
rect 5632 2320 5684 2372
rect 6920 2388 6972 2440
rect 8116 2388 8168 2440
rect 9036 2388 9088 2440
rect 7012 2320 7064 2372
rect 2964 2252 3016 2304
rect 3700 2252 3752 2304
rect 4528 2295 4580 2304
rect 4528 2261 4537 2295
rect 4537 2261 4571 2295
rect 4571 2261 4580 2295
rect 4528 2252 4580 2261
rect 6920 2252 6972 2304
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 7380 2252 7432 2304
rect 10048 2320 10100 2372
rect 10324 2363 10376 2372
rect 10324 2329 10333 2363
rect 10333 2329 10367 2363
rect 10367 2329 10376 2363
rect 10324 2320 10376 2329
rect 10784 2388 10836 2440
rect 11152 2456 11204 2508
rect 11336 2388 11388 2440
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 14004 2524 14056 2576
rect 16672 2524 16724 2576
rect 23848 2524 23900 2576
rect 43260 2524 43312 2576
rect 46756 2524 46808 2576
rect 49424 2524 49476 2576
rect 12348 2388 12400 2440
rect 12532 2388 12584 2440
rect 15384 2456 15436 2508
rect 22928 2456 22980 2508
rect 24768 2456 24820 2508
rect 26884 2456 26936 2508
rect 12256 2320 12308 2372
rect 12716 2363 12768 2372
rect 12716 2329 12725 2363
rect 12725 2329 12759 2363
rect 12759 2329 12768 2363
rect 12716 2320 12768 2329
rect 9220 2252 9272 2304
rect 9680 2295 9732 2304
rect 9680 2261 9689 2295
rect 9689 2261 9723 2295
rect 9723 2261 9732 2295
rect 9680 2252 9732 2261
rect 12072 2252 12124 2304
rect 15476 2388 15528 2440
rect 15660 2388 15712 2440
rect 17592 2388 17644 2440
rect 18604 2431 18656 2440
rect 18604 2397 18613 2431
rect 18613 2397 18647 2431
rect 18647 2397 18656 2431
rect 18604 2388 18656 2397
rect 18788 2388 18840 2440
rect 19340 2388 19392 2440
rect 20260 2388 20312 2440
rect 21180 2388 21232 2440
rect 22100 2388 22152 2440
rect 22652 2388 22704 2440
rect 25780 2388 25832 2440
rect 27712 2388 27764 2440
rect 17408 2320 17460 2372
rect 30932 2456 30984 2508
rect 41328 2456 41380 2508
rect 29828 2388 29880 2440
rect 30748 2388 30800 2440
rect 31668 2388 31720 2440
rect 32588 2388 32640 2440
rect 33784 2431 33836 2440
rect 33784 2397 33793 2431
rect 33793 2397 33827 2431
rect 33827 2397 33836 2431
rect 33784 2388 33836 2397
rect 34336 2388 34388 2440
rect 34980 2388 35032 2440
rect 35532 2388 35584 2440
rect 36728 2388 36780 2440
rect 37648 2388 37700 2440
rect 38844 2431 38896 2440
rect 38844 2397 38853 2431
rect 38853 2397 38887 2431
rect 38887 2397 38896 2431
rect 38844 2388 38896 2397
rect 39764 2388 39816 2440
rect 40960 2431 41012 2440
rect 40960 2397 40969 2431
rect 40969 2397 41003 2431
rect 41003 2397 41012 2431
rect 40960 2388 41012 2397
rect 41512 2388 41564 2440
rect 42432 2431 42484 2440
rect 42432 2397 42441 2431
rect 42441 2397 42475 2431
rect 42475 2397 42484 2431
rect 42432 2388 42484 2397
rect 43628 2388 43680 2440
rect 44272 2388 44324 2440
rect 44824 2388 44876 2440
rect 29184 2320 29236 2372
rect 14188 2295 14240 2304
rect 14188 2261 14197 2295
rect 14197 2261 14231 2295
rect 14231 2261 14240 2295
rect 14188 2252 14240 2261
rect 17776 2252 17828 2304
rect 47124 2388 47176 2440
rect 49700 2320 49752 2372
rect 49240 2252 49292 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 20 2048 72 2100
rect 27896 2048 27948 2100
rect 5908 1980 5960 2032
rect 9404 1980 9456 2032
rect 10048 1980 10100 2032
rect 13912 1980 13964 2032
rect 7564 1912 7616 1964
rect 8300 1912 8352 1964
rect 8392 1912 8444 1964
rect 14188 1912 14240 1964
rect 12348 1844 12400 1896
rect 12716 1844 12768 1896
rect 17408 1844 17460 1896
rect 3148 1776 3200 1828
rect 3608 1776 3660 1828
rect 6920 1776 6972 1828
rect 13544 1776 13596 1828
rect 4712 1708 4764 1760
rect 5632 1708 5684 1760
rect 7104 1708 7156 1760
rect 15108 1708 15160 1760
rect 3608 1640 3660 1692
rect 3884 1640 3936 1692
rect 7288 1572 7340 1624
rect 8024 1572 8076 1624
rect 8300 1572 8352 1624
rect 9496 1572 9548 1624
rect 9680 1640 9732 1692
rect 20168 1640 20220 1692
rect 11980 1572 12032 1624
rect 13360 1572 13412 1624
rect 15016 1572 15068 1624
rect 4528 1504 4580 1556
rect 13268 1504 13320 1556
rect 4528 1300 4580 1352
rect 5172 1300 5224 1352
rect 7380 1436 7432 1488
rect 9220 1436 9272 1488
rect 18604 1436 18656 1488
rect 7012 1368 7064 1420
rect 7748 1368 7800 1420
rect 7380 1343 7432 1352
rect 7380 1309 7389 1343
rect 7389 1309 7423 1343
rect 7423 1309 7432 1343
rect 7380 1300 7432 1309
rect 7748 1232 7800 1284
rect 8392 1368 8444 1420
rect 9036 1368 9088 1420
rect 9312 1368 9364 1420
rect 9496 1368 9548 1420
rect 10048 1368 10100 1420
rect 10600 1368 10652 1420
rect 11336 1368 11388 1420
rect 17316 1368 17368 1420
rect 9220 1300 9272 1352
rect 9772 1300 9824 1352
rect 12348 1300 12400 1352
rect 12440 1300 12492 1352
rect 14648 1300 14700 1352
rect 44456 1300 44508 1352
rect 46480 1300 46532 1352
rect 10140 1232 10192 1284
rect 14740 1232 14792 1284
rect 4160 1164 4212 1216
rect 4804 1164 4856 1216
rect 5908 1164 5960 1216
rect 10324 1164 10376 1216
rect 10784 1164 10836 1216
rect 8392 1096 8444 1148
rect 11060 1096 11112 1148
rect 9680 1028 9732 1080
rect 11704 1028 11756 1080
rect 12808 1028 12860 1080
rect 14924 1028 14976 1080
rect 10692 960 10744 1012
rect 12624 960 12676 1012
rect 5264 892 5316 944
rect 6920 892 6972 944
rect 8852 935 8904 944
rect 8852 901 8861 935
rect 8861 901 8895 935
rect 8895 901 8904 935
rect 8852 892 8904 901
<< metal2 >>
rect 202 49200 258 50000
rect 570 49200 626 50000
rect 1030 49200 1086 50000
rect 1398 49200 1454 50000
rect 1858 49200 1914 50000
rect 2226 49200 2282 50000
rect 2686 49200 2742 50000
rect 3054 49200 3110 50000
rect 3514 49200 3570 50000
rect 3882 49200 3938 50000
rect 4342 49200 4398 50000
rect 4710 49200 4766 50000
rect 5170 49200 5226 50000
rect 5538 49200 5594 50000
rect 5998 49200 6054 50000
rect 6366 49200 6422 50000
rect 6826 49200 6882 50000
rect 7194 49200 7250 50000
rect 7654 49200 7710 50000
rect 8022 49200 8078 50000
rect 8482 49200 8538 50000
rect 8942 49200 8998 50000
rect 9310 49200 9366 50000
rect 9770 49200 9826 50000
rect 10138 49200 10194 50000
rect 10598 49200 10654 50000
rect 10966 49200 11022 50000
rect 11426 49200 11482 50000
rect 11794 49200 11850 50000
rect 12254 49200 12310 50000
rect 12622 49200 12678 50000
rect 13082 49200 13138 50000
rect 13450 49200 13506 50000
rect 13910 49200 13966 50000
rect 14278 49200 14334 50000
rect 14738 49200 14794 50000
rect 15106 49200 15162 50000
rect 15566 49200 15622 50000
rect 15934 49200 15990 50000
rect 16394 49200 16450 50000
rect 16854 49200 16910 50000
rect 17222 49200 17278 50000
rect 17682 49200 17738 50000
rect 18050 49200 18106 50000
rect 18510 49200 18566 50000
rect 18878 49200 18934 50000
rect 19338 49200 19394 50000
rect 19706 49200 19762 50000
rect 20166 49200 20222 50000
rect 20534 49200 20590 50000
rect 20994 49200 21050 50000
rect 21362 49200 21418 50000
rect 21822 49200 21878 50000
rect 22190 49200 22246 50000
rect 22650 49200 22706 50000
rect 23018 49200 23074 50000
rect 23478 49200 23534 50000
rect 23846 49200 23902 50000
rect 24306 49200 24362 50000
rect 24674 49200 24730 50000
rect 25134 49200 25190 50000
rect 25594 49200 25650 50000
rect 25962 49200 26018 50000
rect 26422 49200 26478 50000
rect 26790 49200 26846 50000
rect 27250 49200 27306 50000
rect 27618 49200 27674 50000
rect 28078 49200 28134 50000
rect 28446 49200 28502 50000
rect 28906 49200 28962 50000
rect 29274 49200 29330 50000
rect 29734 49200 29790 50000
rect 30102 49200 30158 50000
rect 30562 49200 30618 50000
rect 30930 49200 30986 50000
rect 31390 49200 31446 50000
rect 31758 49200 31814 50000
rect 32218 49200 32274 50000
rect 32586 49200 32642 50000
rect 33046 49200 33102 50000
rect 33506 49200 33562 50000
rect 33874 49200 33930 50000
rect 34334 49200 34390 50000
rect 34702 49200 34758 50000
rect 35162 49200 35218 50000
rect 35530 49200 35586 50000
rect 35990 49200 36046 50000
rect 36358 49200 36414 50000
rect 36818 49200 36874 50000
rect 37186 49200 37242 50000
rect 37646 49200 37702 50000
rect 38014 49200 38070 50000
rect 38474 49200 38530 50000
rect 38842 49200 38898 50000
rect 39302 49200 39358 50000
rect 39670 49200 39726 50000
rect 40130 49200 40186 50000
rect 40498 49200 40554 50000
rect 40958 49200 41014 50000
rect 41326 49200 41382 50000
rect 41786 49200 41842 50000
rect 42246 49200 42302 50000
rect 42614 49200 42670 50000
rect 43074 49200 43130 50000
rect 43442 49200 43498 50000
rect 43902 49200 43958 50000
rect 44270 49200 44326 50000
rect 44730 49200 44786 50000
rect 45098 49200 45154 50000
rect 45558 49200 45614 50000
rect 45926 49200 45982 50000
rect 46386 49200 46442 50000
rect 46478 49736 46534 49745
rect 46478 49671 46534 49680
rect 584 46714 612 49200
rect 1044 46918 1072 49200
rect 1490 47288 1546 47297
rect 1872 47258 1900 49200
rect 1490 47223 1492 47232
rect 1544 47223 1546 47232
rect 1860 47252 1912 47258
rect 1492 47194 1544 47200
rect 1860 47194 1912 47200
rect 1676 47048 1728 47054
rect 1676 46990 1728 46996
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 1032 46912 1084 46918
rect 1032 46854 1084 46860
rect 572 46708 624 46714
rect 572 46650 624 46656
rect 1688 46170 1716 46990
rect 1676 46164 1728 46170
rect 1676 46106 1728 46112
rect 1964 45354 1992 46990
rect 2240 46714 2268 49200
rect 3068 47258 3096 49200
rect 3056 47252 3108 47258
rect 3056 47194 3108 47200
rect 2872 47048 2924 47054
rect 2872 46990 2924 46996
rect 2228 46708 2280 46714
rect 2228 46650 2280 46656
rect 2504 46572 2556 46578
rect 2504 46514 2556 46520
rect 2596 46572 2648 46578
rect 2596 46514 2648 46520
rect 2516 46170 2544 46514
rect 2504 46164 2556 46170
rect 2504 46106 2556 46112
rect 2044 45960 2096 45966
rect 2044 45902 2096 45908
rect 1952 45348 2004 45354
rect 1952 45290 2004 45296
rect 2056 44742 2084 45902
rect 2504 45484 2556 45490
rect 2504 45426 2556 45432
rect 2516 45082 2544 45426
rect 2504 45076 2556 45082
rect 2504 45018 2556 45024
rect 2044 44736 2096 44742
rect 2044 44678 2096 44684
rect 2056 43790 2084 44678
rect 2044 43784 2096 43790
rect 2044 43726 2096 43732
rect 848 43104 900 43110
rect 848 43046 900 43052
rect 664 13864 716 13870
rect 664 13806 716 13812
rect 388 8968 440 8974
rect 388 8910 440 8916
rect 296 7880 348 7886
rect 296 7822 348 7828
rect 204 5024 256 5030
rect 204 4966 256 4972
rect 112 3052 164 3058
rect 112 2994 164 3000
rect 20 2100 72 2106
rect 20 2042 72 2048
rect 32 800 60 2042
rect 124 800 152 2994
rect 216 800 244 4966
rect 308 800 336 7822
rect 400 800 428 8910
rect 572 6928 624 6934
rect 572 6870 624 6876
rect 480 6792 532 6798
rect 480 6734 532 6740
rect 492 2774 520 6734
rect 584 2922 612 6870
rect 676 4758 704 13806
rect 756 9920 808 9926
rect 756 9862 808 9868
rect 768 7954 796 9862
rect 756 7948 808 7954
rect 756 7890 808 7896
rect 664 4752 716 4758
rect 664 4694 716 4700
rect 756 4140 808 4146
rect 756 4082 808 4088
rect 664 3528 716 3534
rect 664 3470 716 3476
rect 572 2916 624 2922
rect 572 2858 624 2864
rect 492 2746 612 2774
rect 480 2440 532 2446
rect 480 2382 532 2388
rect 492 800 520 2382
rect 584 800 612 2746
rect 676 800 704 3470
rect 768 800 796 4082
rect 860 3738 888 43046
rect 1952 42220 2004 42226
rect 1952 42162 2004 42168
rect 1492 42016 1544 42022
rect 1492 41958 1544 41964
rect 1504 41721 1532 41958
rect 1964 41818 1992 42162
rect 1952 41812 2004 41818
rect 1952 41754 2004 41760
rect 1490 41712 1546 41721
rect 1490 41647 1546 41656
rect 1490 36136 1546 36145
rect 1490 36071 1546 36080
rect 1504 36038 1532 36071
rect 1492 36032 1544 36038
rect 1492 35974 1544 35980
rect 1492 30592 1544 30598
rect 1490 30560 1492 30569
rect 1544 30560 1546 30569
rect 1490 30495 1546 30504
rect 1676 25288 1728 25294
rect 1676 25230 1728 25236
rect 1492 25152 1544 25158
rect 1492 25094 1544 25100
rect 1504 24993 1532 25094
rect 1490 24984 1546 24993
rect 1688 24954 1716 25230
rect 1490 24919 1546 24928
rect 1676 24948 1728 24954
rect 1676 24890 1728 24896
rect 1216 20596 1268 20602
rect 1216 20538 1268 20544
rect 1124 19304 1176 19310
rect 1124 19246 1176 19252
rect 940 9988 992 9994
rect 940 9930 992 9936
rect 848 3732 900 3738
rect 848 3674 900 3680
rect 952 3618 980 9930
rect 1136 6118 1164 19246
rect 1228 9926 1256 20538
rect 1952 19848 2004 19854
rect 1952 19790 2004 19796
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1504 19417 1532 19654
rect 1964 19514 1992 19790
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 1490 13832 1546 13841
rect 1490 13767 1492 13776
rect 1544 13767 1546 13776
rect 1492 13738 1544 13744
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1216 9920 1268 9926
rect 1216 9862 1268 9868
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1216 9716 1268 9722
rect 1216 9658 1268 9664
rect 1124 6112 1176 6118
rect 1124 6054 1176 6060
rect 1032 5908 1084 5914
rect 1032 5850 1084 5856
rect 1044 4706 1072 5850
rect 1124 5840 1176 5846
rect 1124 5782 1176 5788
rect 1136 5114 1164 5782
rect 1228 5234 1256 9658
rect 1308 9648 1360 9654
rect 1308 9590 1360 9596
rect 1320 5302 1348 9590
rect 1412 8974 1440 9862
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1504 8514 1532 9318
rect 1412 8486 1532 8514
rect 1412 7886 1440 8486
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 8265 1532 8298
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1504 7732 1532 8026
rect 1412 7704 1532 7732
rect 1412 7274 1440 7704
rect 1596 7290 1624 11018
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1400 7268 1452 7274
rect 1400 7210 1452 7216
rect 1504 7262 1624 7290
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 1308 5296 1360 5302
rect 1308 5238 1360 5244
rect 1216 5228 1268 5234
rect 1216 5170 1268 5176
rect 1136 5086 1348 5114
rect 1044 4678 1164 4706
rect 1032 4616 1084 4622
rect 1032 4558 1084 4564
rect 860 3590 980 3618
rect 860 2446 888 3590
rect 940 3324 992 3330
rect 940 3266 992 3272
rect 848 2440 900 2446
rect 848 2382 900 2388
rect 952 800 980 3266
rect 1044 800 1072 4558
rect 1136 3942 1164 4678
rect 1124 3936 1176 3942
rect 1124 3878 1176 3884
rect 1320 2774 1348 5086
rect 1412 3194 1440 6598
rect 1504 5710 1532 7262
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6254 1624 7142
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1504 4146 1532 5510
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1492 4004 1544 4010
rect 1492 3946 1544 3952
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 1504 2774 1532 3946
rect 1228 2746 1348 2774
rect 1412 2746 1532 2774
rect 1228 800 1256 2746
rect 1412 800 1440 2746
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 1504 800 1532 2586
rect 1596 800 1624 6054
rect 1688 3058 1716 10406
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1780 4622 1808 9318
rect 1872 6322 1900 11494
rect 2056 11121 2084 43726
rect 2320 43308 2372 43314
rect 2320 43250 2372 43256
rect 2332 42838 2360 43250
rect 2320 42832 2372 42838
rect 2320 42774 2372 42780
rect 2608 42702 2636 46514
rect 2780 45960 2832 45966
rect 2780 45902 2832 45908
rect 2792 45558 2820 45902
rect 2780 45552 2832 45558
rect 2780 45494 2832 45500
rect 2688 45280 2740 45286
rect 2688 45222 2740 45228
rect 2700 44878 2728 45222
rect 2688 44872 2740 44878
rect 2688 44814 2740 44820
rect 2688 44736 2740 44742
rect 2688 44678 2740 44684
rect 2700 43314 2728 44678
rect 2792 44334 2820 45494
rect 2780 44328 2832 44334
rect 2780 44270 2832 44276
rect 2780 44192 2832 44198
rect 2780 44134 2832 44140
rect 2688 43308 2740 43314
rect 2688 43250 2740 43256
rect 2700 42770 2728 43250
rect 2792 43178 2820 44134
rect 2884 43994 2912 46990
rect 3528 46714 3556 49200
rect 4356 48090 4384 49200
rect 4356 48062 4660 48090
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4632 47258 4660 48062
rect 4724 47258 4752 49200
rect 5552 47258 5580 49200
rect 4620 47252 4672 47258
rect 4620 47194 4672 47200
rect 4712 47252 4764 47258
rect 4712 47194 4764 47200
rect 5540 47252 5592 47258
rect 5540 47194 5592 47200
rect 3792 47048 3844 47054
rect 3792 46990 3844 46996
rect 4804 47048 4856 47054
rect 4804 46990 4856 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 3516 46708 3568 46714
rect 3516 46650 3568 46656
rect 3056 46572 3108 46578
rect 3056 46514 3108 46520
rect 3068 46034 3096 46514
rect 3608 46368 3660 46374
rect 3608 46310 3660 46316
rect 3056 46028 3108 46034
rect 3056 45970 3108 45976
rect 3068 44878 3096 45970
rect 3620 44878 3648 46310
rect 3804 46170 3832 46990
rect 4816 46714 4844 46990
rect 4804 46708 4856 46714
rect 4804 46650 4856 46656
rect 4160 46572 4212 46578
rect 4160 46514 4212 46520
rect 4172 46458 4200 46514
rect 4080 46430 4200 46458
rect 3792 46164 3844 46170
rect 4080 46152 4108 46430
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4080 46124 4200 46152
rect 3792 46106 3844 46112
rect 4172 45354 4200 46124
rect 5264 45892 5316 45898
rect 5264 45834 5316 45840
rect 4988 45824 5040 45830
rect 4988 45766 5040 45772
rect 4526 45520 4582 45529
rect 4894 45520 4950 45529
rect 4526 45455 4528 45464
rect 4580 45455 4582 45464
rect 4712 45484 4764 45490
rect 4528 45426 4580 45432
rect 4894 45455 4950 45464
rect 4712 45426 4764 45432
rect 4620 45416 4672 45422
rect 4620 45358 4672 45364
rect 4160 45348 4212 45354
rect 4160 45290 4212 45296
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4632 45082 4660 45358
rect 4620 45076 4672 45082
rect 4620 45018 4672 45024
rect 3056 44872 3108 44878
rect 3056 44814 3108 44820
rect 3608 44872 3660 44878
rect 3608 44814 3660 44820
rect 3068 44266 3096 44814
rect 4724 44810 4752 45426
rect 4804 45416 4856 45422
rect 4804 45358 4856 45364
rect 4816 44946 4844 45358
rect 4804 44940 4856 44946
rect 4804 44882 4856 44888
rect 4344 44804 4396 44810
rect 4344 44746 4396 44752
rect 4712 44804 4764 44810
rect 4712 44746 4764 44752
rect 3884 44736 3936 44742
rect 3884 44678 3936 44684
rect 3056 44260 3108 44266
rect 3056 44202 3108 44208
rect 2872 43988 2924 43994
rect 2872 43930 2924 43936
rect 2884 43314 2912 43930
rect 2964 43716 3016 43722
rect 2964 43658 3016 43664
rect 2976 43450 3004 43658
rect 2964 43444 3016 43450
rect 2964 43386 3016 43392
rect 2872 43308 2924 43314
rect 2872 43250 2924 43256
rect 2780 43172 2832 43178
rect 2780 43114 2832 43120
rect 2688 42764 2740 42770
rect 2688 42706 2740 42712
rect 2596 42696 2648 42702
rect 2792 42680 2820 43114
rect 2596 42638 2648 42644
rect 2780 42674 2832 42680
rect 2320 42560 2372 42566
rect 2320 42502 2372 42508
rect 2332 42294 2360 42502
rect 2320 42288 2372 42294
rect 2320 42230 2372 42236
rect 2608 42090 2636 42638
rect 2780 42616 2832 42622
rect 2596 42084 2648 42090
rect 2596 42026 2648 42032
rect 2792 41750 2820 42616
rect 2780 41744 2832 41750
rect 2780 41686 2832 41692
rect 2596 41608 2648 41614
rect 2596 41550 2648 41556
rect 2608 20602 2636 41550
rect 2872 30592 2924 30598
rect 2872 30534 2924 30540
rect 2688 24812 2740 24818
rect 2688 24754 2740 24760
rect 2700 24614 2728 24754
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2596 20596 2648 20602
rect 2596 20538 2648 20544
rect 2042 11112 2098 11121
rect 2042 11047 2098 11056
rect 2596 11076 2648 11082
rect 2596 11018 2648 11024
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2044 9988 2096 9994
rect 2044 9930 2096 9936
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1860 6180 1912 6186
rect 1860 6122 1912 6128
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1766 4448 1822 4457
rect 1766 4383 1822 4392
rect 1780 3126 1808 4383
rect 1872 4282 1900 6122
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1964 4214 1992 9454
rect 2056 8090 2084 9930
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 2056 6798 2084 7686
rect 2148 6866 2176 10406
rect 2240 7410 2268 10406
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2332 8498 2360 8774
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2332 8401 2360 8434
rect 2318 8392 2374 8401
rect 2318 8327 2374 8336
rect 2424 7834 2452 9862
rect 2516 7886 2544 9998
rect 2332 7806 2452 7834
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2332 7478 2360 7806
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2240 7274 2360 7290
rect 2240 7268 2372 7274
rect 2240 7262 2320 7268
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2056 4729 2084 6394
rect 2148 5914 2176 6598
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2136 5636 2188 5642
rect 2136 5578 2188 5584
rect 2148 5234 2176 5578
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2042 4720 2098 4729
rect 2042 4655 2098 4664
rect 2044 4548 2096 4554
rect 2044 4490 2096 4496
rect 1952 4208 2004 4214
rect 1872 4156 1952 4162
rect 1872 4150 2004 4156
rect 1872 4134 1992 4150
rect 1768 3120 1820 3126
rect 1768 3062 1820 3068
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1780 800 1808 2926
rect 1872 800 1900 4134
rect 1952 3664 2004 3670
rect 1952 3606 2004 3612
rect 1964 800 1992 3606
rect 2056 2961 2084 4490
rect 2148 3534 2176 4966
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 2240 3126 2268 7262
rect 2320 7210 2372 7216
rect 2424 7041 2452 7686
rect 2410 7032 2466 7041
rect 2410 6967 2466 6976
rect 2516 6882 2544 7822
rect 2424 6854 2544 6882
rect 2608 6866 2636 11018
rect 2700 9722 2728 24550
rect 2884 16574 2912 30534
rect 2884 16546 3004 16574
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2792 7886 2820 9862
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2596 6860 2648 6866
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2332 4826 2360 6734
rect 2424 6458 2452 6854
rect 2596 6802 2648 6808
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2318 4176 2374 4185
rect 2318 4111 2320 4120
rect 2372 4111 2374 4120
rect 2320 4082 2372 4088
rect 2318 4040 2374 4049
rect 2318 3975 2374 3984
rect 2136 3120 2188 3126
rect 2136 3062 2188 3068
rect 2228 3120 2280 3126
rect 2228 3062 2280 3068
rect 2042 2952 2098 2961
rect 2042 2887 2098 2896
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 2056 2514 2084 2790
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 2148 800 2176 3062
rect 2226 2680 2282 2689
rect 2226 2615 2282 2624
rect 2240 800 2268 2615
rect 2332 2446 2360 3975
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2424 800 2452 6054
rect 2516 2650 2544 6394
rect 2608 5710 2636 6802
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2516 800 2544 2450
rect 2608 800 2636 4762
rect 2700 2854 2728 7482
rect 2792 7313 2820 7822
rect 2778 7304 2834 7313
rect 2778 7239 2834 7248
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 6769 2820 7142
rect 2778 6760 2834 6769
rect 2778 6695 2834 6704
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2792 3369 2820 6598
rect 2884 5234 2912 9318
rect 2976 8945 3004 16546
rect 3068 12434 3096 44202
rect 3896 43926 3924 44678
rect 4356 44334 4384 44746
rect 4344 44328 4396 44334
rect 4344 44270 4396 44276
rect 4804 44328 4856 44334
rect 4804 44270 4856 44276
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 3884 43920 3936 43926
rect 3884 43862 3936 43868
rect 4620 43920 4672 43926
rect 4620 43862 4672 43868
rect 3516 43716 3568 43722
rect 3516 43658 3568 43664
rect 3528 43314 3556 43658
rect 3516 43308 3568 43314
rect 3516 43250 3568 43256
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4632 42838 4660 43862
rect 4816 43654 4844 44270
rect 4804 43648 4856 43654
rect 4804 43590 4856 43596
rect 4712 43308 4764 43314
rect 4712 43250 4764 43256
rect 4724 42906 4752 43250
rect 4816 43110 4844 43590
rect 4804 43104 4856 43110
rect 4804 43046 4856 43052
rect 4712 42900 4764 42906
rect 4712 42842 4764 42848
rect 4252 42832 4304 42838
rect 4252 42774 4304 42780
rect 4620 42832 4672 42838
rect 4620 42774 4672 42780
rect 3240 42560 3292 42566
rect 3240 42502 3292 42508
rect 3068 12406 3188 12434
rect 2962 8936 3018 8945
rect 2962 8871 3018 8880
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2976 5658 3004 8774
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3068 7041 3096 7686
rect 3054 7032 3110 7041
rect 3054 6967 3110 6976
rect 2976 5630 3096 5658
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2884 4826 2912 5170
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2976 4128 3004 5510
rect 3068 4282 3096 5630
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2884 4100 3004 4128
rect 2884 3670 2912 4100
rect 3054 4040 3110 4049
rect 2964 4004 3016 4010
rect 3054 3975 3110 3984
rect 2964 3946 3016 3952
rect 2872 3664 2924 3670
rect 2976 3641 3004 3946
rect 2872 3606 2924 3612
rect 2962 3632 3018 3641
rect 2962 3567 3018 3576
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2778 3360 2834 3369
rect 2778 3295 2834 3304
rect 2870 3224 2926 3233
rect 2780 3188 2832 3194
rect 2870 3159 2872 3168
rect 2780 3130 2832 3136
rect 2924 3159 2926 3168
rect 2872 3130 2924 3136
rect 2792 3040 2820 3130
rect 2872 3052 2924 3058
rect 2792 3012 2872 3040
rect 2872 2994 2924 3000
rect 2778 2952 2834 2961
rect 2976 2904 3004 3402
rect 2778 2887 2834 2896
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2700 800 2728 2586
rect 2792 800 2820 2887
rect 2884 2876 3004 2904
rect 2884 2650 2912 2876
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 3068 2514 3096 3975
rect 3160 3738 3188 12406
rect 3252 8294 3280 42502
rect 4264 42362 4292 42774
rect 4528 42764 4580 42770
rect 4528 42706 4580 42712
rect 4252 42356 4304 42362
rect 4252 42298 4304 42304
rect 4540 42242 4568 42706
rect 4712 42696 4764 42702
rect 4816 42684 4844 43046
rect 4908 42702 4936 45455
rect 5000 45422 5028 45766
rect 5276 45626 5304 45834
rect 5828 45830 5856 46990
rect 6012 46442 6040 49200
rect 6840 47274 6868 49200
rect 6840 47258 6960 47274
rect 6840 47252 6972 47258
rect 6840 47246 6920 47252
rect 6920 47194 6972 47200
rect 6368 47048 6420 47054
rect 6368 46990 6420 46996
rect 6380 46714 6408 46990
rect 7208 46714 7236 49200
rect 8036 48090 8064 49200
rect 8036 48062 8340 48090
rect 8312 47258 8340 48062
rect 8300 47252 8352 47258
rect 8300 47194 8352 47200
rect 7380 47048 7432 47054
rect 7380 46990 7432 46996
rect 8024 47048 8076 47054
rect 8024 46990 8076 46996
rect 6368 46708 6420 46714
rect 6368 46650 6420 46656
rect 7196 46708 7248 46714
rect 7196 46650 7248 46656
rect 6368 46572 6420 46578
rect 6368 46514 6420 46520
rect 6000 46436 6052 46442
rect 6000 46378 6052 46384
rect 5816 45824 5868 45830
rect 5816 45766 5868 45772
rect 5264 45620 5316 45626
rect 5264 45562 5316 45568
rect 5828 45490 5856 45766
rect 5816 45484 5868 45490
rect 5816 45426 5868 45432
rect 4988 45416 5040 45422
rect 4988 45358 5040 45364
rect 5000 45014 5028 45358
rect 5448 45076 5500 45082
rect 5448 45018 5500 45024
rect 4988 45008 5040 45014
rect 4988 44950 5040 44956
rect 5264 44804 5316 44810
rect 5264 44746 5316 44752
rect 4988 44192 5040 44198
rect 4988 44134 5040 44140
rect 5000 43858 5028 44134
rect 4988 43852 5040 43858
rect 4988 43794 5040 43800
rect 5000 43314 5028 43794
rect 4988 43308 5040 43314
rect 4988 43250 5040 43256
rect 4764 42656 4844 42684
rect 4896 42696 4948 42702
rect 4712 42638 4764 42644
rect 4896 42638 4948 42644
rect 4540 42214 4660 42242
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4632 13870 4660 42214
rect 4724 41818 4752 42638
rect 5000 42362 5028 43250
rect 4988 42356 5040 42362
rect 4988 42298 5040 42304
rect 4712 41812 4764 41818
rect 4712 41754 4764 41760
rect 5276 16574 5304 44746
rect 5460 43994 5488 45018
rect 5448 43988 5500 43994
rect 5448 43930 5500 43936
rect 5460 43382 5488 43930
rect 6380 43450 6408 46514
rect 7392 46170 7420 46990
rect 7748 46572 7800 46578
rect 7748 46514 7800 46520
rect 7380 46164 7432 46170
rect 7380 46106 7432 46112
rect 6920 45960 6972 45966
rect 6920 45902 6972 45908
rect 6460 45892 6512 45898
rect 6460 45834 6512 45840
rect 6472 45626 6500 45834
rect 6460 45620 6512 45626
rect 6460 45562 6512 45568
rect 6460 45416 6512 45422
rect 6460 45358 6512 45364
rect 6472 44742 6500 45358
rect 6736 45348 6788 45354
rect 6736 45290 6788 45296
rect 6460 44736 6512 44742
rect 6460 44678 6512 44684
rect 6472 44198 6500 44678
rect 6748 44470 6776 45290
rect 6932 45082 6960 45902
rect 7760 45830 7788 46514
rect 7748 45824 7800 45830
rect 7748 45766 7800 45772
rect 7760 45558 7788 45766
rect 7748 45552 7800 45558
rect 7194 45520 7250 45529
rect 7748 45494 7800 45500
rect 7194 45455 7196 45464
rect 7248 45455 7250 45464
rect 7196 45426 7248 45432
rect 8036 45354 8064 46990
rect 8496 46714 8524 49200
rect 9324 47258 9352 49200
rect 9312 47252 9364 47258
rect 9312 47194 9364 47200
rect 9784 47138 9812 49200
rect 10612 47258 10640 49200
rect 10600 47252 10652 47258
rect 10600 47194 10652 47200
rect 9784 47110 9904 47138
rect 9772 47048 9824 47054
rect 9772 46990 9824 46996
rect 8944 46980 8996 46986
rect 8944 46922 8996 46928
rect 8484 46708 8536 46714
rect 8484 46650 8536 46656
rect 8116 46572 8168 46578
rect 8116 46514 8168 46520
rect 7012 45348 7064 45354
rect 7012 45290 7064 45296
rect 8024 45348 8076 45354
rect 8024 45290 8076 45296
rect 6920 45076 6972 45082
rect 6920 45018 6972 45024
rect 6736 44464 6788 44470
rect 6736 44406 6788 44412
rect 6460 44192 6512 44198
rect 6460 44134 6512 44140
rect 5816 43444 5868 43450
rect 5816 43386 5868 43392
rect 6368 43444 6420 43450
rect 6368 43386 6420 43392
rect 5448 43376 5500 43382
rect 5448 43318 5500 43324
rect 5828 42702 5856 43386
rect 5816 42696 5868 42702
rect 5816 42638 5868 42644
rect 6368 42696 6420 42702
rect 6368 42638 6420 42644
rect 6380 42566 6408 42638
rect 6368 42560 6420 42566
rect 6368 42502 6420 42508
rect 6472 26234 6500 44134
rect 6748 42770 6776 44406
rect 6828 43308 6880 43314
rect 6932 43296 6960 45018
rect 7024 44946 7052 45290
rect 7012 44940 7064 44946
rect 7012 44882 7064 44888
rect 7024 43926 7052 44882
rect 7012 43920 7064 43926
rect 7012 43862 7064 43868
rect 7024 43466 7052 43862
rect 7024 43438 7144 43466
rect 8128 43450 8156 46514
rect 8956 46034 8984 46922
rect 9404 46368 9456 46374
rect 9404 46310 9456 46316
rect 8944 46028 8996 46034
rect 8944 45970 8996 45976
rect 8392 45960 8444 45966
rect 8392 45902 8444 45908
rect 8404 45558 8432 45902
rect 9416 45898 9444 46310
rect 9312 45892 9364 45898
rect 9312 45834 9364 45840
rect 9404 45892 9456 45898
rect 9404 45834 9456 45840
rect 9324 45626 9352 45834
rect 9312 45620 9364 45626
rect 9312 45562 9364 45568
rect 8392 45552 8444 45558
rect 8392 45494 8444 45500
rect 8300 45416 8352 45422
rect 8300 45358 8352 45364
rect 8312 44742 8340 45358
rect 8404 45082 8432 45494
rect 8852 45484 8904 45490
rect 8852 45426 8904 45432
rect 8392 45076 8444 45082
rect 8392 45018 8444 45024
rect 8300 44736 8352 44742
rect 8300 44678 8352 44684
rect 8208 43852 8260 43858
rect 8208 43794 8260 43800
rect 6880 43268 6960 43296
rect 6828 43250 6880 43256
rect 6736 42764 6788 42770
rect 6736 42706 6788 42712
rect 6552 42696 6604 42702
rect 6552 42638 6604 42644
rect 6564 42022 6592 42638
rect 6932 42362 6960 43268
rect 7012 43308 7064 43314
rect 7012 43250 7064 43256
rect 7024 42906 7052 43250
rect 7012 42900 7064 42906
rect 7012 42842 7064 42848
rect 7116 42634 7144 43438
rect 8116 43444 8168 43450
rect 8116 43386 8168 43392
rect 8128 42770 8156 43386
rect 8116 42764 8168 42770
rect 8116 42706 8168 42712
rect 8220 42702 8248 43794
rect 8208 42696 8260 42702
rect 8208 42638 8260 42644
rect 7104 42628 7156 42634
rect 7104 42570 7156 42576
rect 7748 42560 7800 42566
rect 7746 42528 7748 42537
rect 7800 42528 7802 42537
rect 7746 42463 7802 42472
rect 6920 42356 6972 42362
rect 6920 42298 6972 42304
rect 6552 42016 6604 42022
rect 6552 41958 6604 41964
rect 5000 16546 5304 16574
rect 6288 26206 6500 26234
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3252 6798 3280 8230
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3252 5642 3280 6258
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 3252 5545 3280 5578
rect 3238 5536 3294 5545
rect 3238 5471 3294 5480
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3252 4554 3280 5306
rect 3240 4548 3292 4554
rect 3240 4490 3292 4496
rect 3238 4448 3294 4457
rect 3238 4383 3294 4392
rect 3252 4146 3280 4383
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3252 3738 3280 3878
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3160 3194 3188 3334
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3146 3088 3202 3097
rect 3146 3023 3202 3032
rect 3160 2650 3188 3023
rect 3238 2952 3294 2961
rect 3238 2887 3294 2896
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3252 2446 3280 2887
rect 3240 2440 3292 2446
rect 3054 2408 3110 2417
rect 3240 2382 3292 2388
rect 3054 2343 3110 2352
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 2870 2000 2926 2009
rect 2870 1935 2926 1944
rect 2884 800 2912 1935
rect 2976 800 3004 2246
rect 3068 800 3096 2343
rect 3238 2272 3294 2281
rect 3238 2207 3294 2216
rect 3148 1828 3200 1834
rect 3148 1770 3200 1776
rect 3160 800 3188 1770
rect 3252 800 3280 2207
rect 3344 800 3372 8434
rect 3436 7002 3464 11018
rect 3884 10532 3936 10538
rect 3884 10474 3936 10480
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3528 7410 3556 10406
rect 3896 10062 3924 10474
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3528 6934 3556 7346
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3436 2990 3464 6666
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3528 2689 3556 6598
rect 3620 5370 3648 8774
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3712 5302 3740 9318
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3804 7041 3832 7686
rect 3790 7032 3846 7041
rect 3790 6967 3846 6976
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3804 6225 3832 6734
rect 3790 6216 3846 6225
rect 3790 6151 3846 6160
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3700 5296 3752 5302
rect 3620 5244 3700 5250
rect 3620 5238 3752 5244
rect 3620 5222 3740 5238
rect 3514 2680 3570 2689
rect 3514 2615 3570 2624
rect 3514 2544 3570 2553
rect 3514 2479 3570 2488
rect 3528 800 3556 2479
rect 3620 1834 3648 5222
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3712 4321 3740 5102
rect 3698 4312 3754 4321
rect 3698 4247 3754 4256
rect 3700 4208 3752 4214
rect 3700 4150 3752 4156
rect 3712 3670 3740 4150
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3712 3194 3740 3470
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3698 2952 3754 2961
rect 3698 2887 3700 2896
rect 3752 2887 3754 2896
rect 3700 2858 3752 2864
rect 3804 2496 3832 6054
rect 3896 3194 3924 8230
rect 3988 7449 4016 11018
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4080 7886 4108 10406
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4632 10146 4660 11018
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4540 10118 4660 10146
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9489 4200 9998
rect 4158 9480 4214 9489
rect 4540 9450 4568 10118
rect 4158 9415 4214 9424
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4344 8832 4396 8838
rect 4342 8800 4344 8809
rect 4396 8800 4398 8809
rect 4342 8735 4398 8744
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4068 7880 4120 7886
rect 4528 7880 4580 7886
rect 4068 7822 4120 7828
rect 4526 7848 4528 7857
rect 4580 7848 4582 7857
rect 3974 7440 4030 7449
rect 3974 7375 4030 7384
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3884 2916 3936 2922
rect 3884 2858 3936 2864
rect 3712 2468 3832 2496
rect 3712 2310 3740 2468
rect 3790 2408 3846 2417
rect 3790 2343 3846 2352
rect 3700 2304 3752 2310
rect 3700 2246 3752 2252
rect 3698 1864 3754 1873
rect 3608 1828 3660 1834
rect 3698 1799 3754 1808
rect 3608 1770 3660 1776
rect 3608 1692 3660 1698
rect 3608 1634 3660 1640
rect 3620 800 3648 1634
rect 3712 800 3740 1799
rect 3804 800 3832 2343
rect 3896 1698 3924 2858
rect 3988 2854 4016 7142
rect 4080 5166 4108 7822
rect 4526 7783 4582 7792
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 7313 4476 7686
rect 4434 7304 4490 7313
rect 4434 7239 4490 7248
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4160 6928 4212 6934
rect 4436 6928 4488 6934
rect 4160 6870 4212 6876
rect 4342 6896 4398 6905
rect 4172 6254 4200 6870
rect 4436 6870 4488 6876
rect 4342 6831 4398 6840
rect 4356 6390 4384 6831
rect 4448 6798 4476 6870
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 6390 4568 6734
rect 4344 6384 4396 6390
rect 4342 6352 4344 6361
rect 4528 6384 4580 6390
rect 4396 6352 4398 6361
rect 4252 6316 4304 6322
rect 4528 6326 4580 6332
rect 4342 6287 4398 6296
rect 4252 6258 4304 6264
rect 4160 6248 4212 6254
rect 4264 6225 4292 6258
rect 4160 6190 4212 6196
rect 4250 6216 4306 6225
rect 4250 6151 4306 6160
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4158 5808 4214 5817
rect 4158 5743 4160 5752
rect 4212 5743 4214 5752
rect 4160 5714 4212 5720
rect 4252 5704 4304 5710
rect 4632 5658 4660 9318
rect 4724 8498 4752 10406
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4710 8392 4766 8401
rect 4710 8327 4712 8336
rect 4764 8327 4766 8336
rect 4712 8298 4764 8304
rect 4712 7404 4764 7410
rect 4816 7392 4844 9318
rect 5000 8906 5028 16546
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4908 8673 4936 8774
rect 4894 8664 4950 8673
rect 5092 8634 5120 9386
rect 4894 8599 4950 8608
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5184 8566 5212 9862
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 4764 7364 4844 7392
rect 4712 7346 4764 7352
rect 4252 5646 4304 5652
rect 4160 5568 4212 5574
rect 4264 5545 4292 5646
rect 4540 5630 4660 5658
rect 4160 5510 4212 5516
rect 4250 5536 4306 5545
rect 4172 5409 4200 5510
rect 4250 5471 4306 5480
rect 4158 5400 4214 5409
rect 4158 5335 4214 5344
rect 4540 5302 4568 5630
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4528 5296 4580 5302
rect 4528 5238 4580 5244
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4172 5012 4200 5238
rect 4080 4984 4200 5012
rect 4080 4808 4108 4984
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4080 4780 4200 4808
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4080 4146 4108 4626
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4172 4026 4200 4780
rect 4526 4720 4582 4729
rect 4526 4655 4582 4664
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4434 4584 4490 4593
rect 4356 4457 4384 4558
rect 4434 4519 4436 4528
rect 4488 4519 4490 4528
rect 4436 4490 4488 4496
rect 4342 4448 4398 4457
rect 4540 4434 4568 4655
rect 4342 4383 4398 4392
rect 4448 4406 4568 4434
rect 4342 4312 4398 4321
rect 4448 4282 4476 4406
rect 4632 4298 4660 5510
rect 4342 4247 4398 4256
rect 4436 4276 4488 4282
rect 4356 4214 4384 4247
rect 4436 4218 4488 4224
rect 4540 4270 4660 4298
rect 4344 4208 4396 4214
rect 4448 4185 4476 4218
rect 4344 4150 4396 4156
rect 4434 4176 4490 4185
rect 4540 4146 4568 4270
rect 4724 4196 4752 7346
rect 4908 6934 4936 8502
rect 5000 7313 5028 8502
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4986 7304 5042 7313
rect 4986 7239 5042 7248
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4896 6928 4948 6934
rect 4802 6896 4858 6905
rect 4896 6870 4948 6876
rect 4802 6831 4858 6840
rect 4816 6322 4844 6831
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4632 4168 4752 4196
rect 4434 4111 4490 4120
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4080 3998 4200 4026
rect 4080 3913 4108 3998
rect 4632 3913 4660 4168
rect 4710 4040 4766 4049
rect 4710 3975 4766 3984
rect 4066 3904 4122 3913
rect 4618 3904 4674 3913
rect 4066 3839 4122 3848
rect 4214 3836 4522 3856
rect 4618 3839 4674 3848
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4526 3496 4582 3505
rect 4250 3360 4306 3369
rect 4250 3295 4306 3304
rect 4264 3058 4292 3295
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4356 2990 4384 3470
rect 4526 3431 4582 3440
rect 4620 3460 4672 3466
rect 4540 3398 4568 3431
rect 4620 3402 4672 3408
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4434 3224 4490 3233
rect 4434 3159 4436 3168
rect 4488 3159 4490 3168
rect 4436 3130 4488 3136
rect 4160 2984 4212 2990
rect 4080 2944 4160 2972
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 3884 1692 3936 1698
rect 3884 1634 3936 1640
rect 4080 1476 4108 2944
rect 4160 2926 4212 2932
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4250 2544 4306 2553
rect 4250 2479 4306 2488
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 3896 1448 4108 1476
rect 3896 800 3924 1448
rect 3974 1320 4030 1329
rect 4172 1306 4200 2314
rect 3974 1255 4030 1264
rect 4080 1278 4200 1306
rect 3988 800 4016 1255
rect 4080 800 4108 1278
rect 4160 1216 4212 1222
rect 4160 1158 4212 1164
rect 4172 800 4200 1158
rect 4264 800 4292 2479
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4356 800 4384 2382
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4540 1562 4568 2246
rect 4528 1556 4580 1562
rect 4528 1498 4580 1504
rect 4632 1442 4660 3402
rect 4724 2378 4752 3975
rect 4712 2372 4764 2378
rect 4712 2314 4764 2320
rect 4712 1760 4764 1766
rect 4712 1702 4764 1708
rect 4448 1414 4660 1442
rect 4448 800 4476 1414
rect 4528 1352 4580 1358
rect 4528 1294 4580 1300
rect 4540 800 4568 1294
rect 4724 800 4752 1702
rect 4816 1222 4844 5510
rect 4908 3738 4936 6598
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5000 3618 5028 7142
rect 5092 6225 5120 8434
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5078 6216 5134 6225
rect 5078 6151 5134 6160
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4908 3590 5028 3618
rect 4908 3126 4936 3590
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4896 3120 4948 3126
rect 4896 3062 4948 3068
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4804 1216 4856 1222
rect 4804 1158 4856 1164
rect 4802 1048 4858 1057
rect 4802 983 4858 992
rect 4816 800 4844 983
rect 4908 800 4936 2926
rect 5000 800 5028 3470
rect 5092 3346 5120 6054
rect 5184 3534 5212 8298
rect 5276 7410 5304 9318
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5092 3318 5212 3346
rect 5078 3224 5134 3233
rect 5078 3159 5134 3168
rect 5092 800 5120 3159
rect 5184 2922 5212 3318
rect 5276 2990 5304 7346
rect 5368 6905 5396 10406
rect 5354 6896 5410 6905
rect 5354 6831 5410 6840
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5368 5137 5396 6734
rect 5460 6254 5488 11018
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 6769 5580 9862
rect 6288 9654 6316 26206
rect 6564 19514 6592 41958
rect 8312 24818 8340 44678
rect 8864 44538 8892 45426
rect 9416 45422 9444 45834
rect 9404 45416 9456 45422
rect 9404 45358 9456 45364
rect 9784 45354 9812 46990
rect 9876 46714 9904 47110
rect 10600 47048 10652 47054
rect 10600 46990 10652 46996
rect 9864 46708 9916 46714
rect 9864 46650 9916 46656
rect 9864 46572 9916 46578
rect 9864 46514 9916 46520
rect 9876 45830 9904 46514
rect 9864 45824 9916 45830
rect 9864 45766 9916 45772
rect 9876 45490 9904 45766
rect 10048 45552 10100 45558
rect 10048 45494 10100 45500
rect 9864 45484 9916 45490
rect 9864 45426 9916 45432
rect 9772 45348 9824 45354
rect 9772 45290 9824 45296
rect 9680 44736 9732 44742
rect 9680 44678 9732 44684
rect 8852 44532 8904 44538
rect 8852 44474 8904 44480
rect 9692 44470 9720 44678
rect 9680 44464 9732 44470
rect 9680 44406 9732 44412
rect 9692 43450 9720 44406
rect 10060 43450 10088 45494
rect 10416 45484 10468 45490
rect 10416 45426 10468 45432
rect 10428 45014 10456 45426
rect 10612 45354 10640 46990
rect 10980 46714 11008 49200
rect 11808 47258 11836 49200
rect 11796 47252 11848 47258
rect 11796 47194 11848 47200
rect 12268 46730 12296 49200
rect 13096 47258 13124 49200
rect 13084 47252 13136 47258
rect 13084 47194 13136 47200
rect 12900 47048 12952 47054
rect 12900 46990 12952 46996
rect 13084 47048 13136 47054
rect 13084 46990 13136 46996
rect 12268 46714 12388 46730
rect 10968 46708 11020 46714
rect 12268 46708 12400 46714
rect 12268 46702 12348 46708
rect 10968 46650 11020 46656
rect 12348 46650 12400 46656
rect 11704 46572 11756 46578
rect 11704 46514 11756 46520
rect 12808 46572 12860 46578
rect 12808 46514 12860 46520
rect 11244 46368 11296 46374
rect 11244 46310 11296 46316
rect 11152 45960 11204 45966
rect 11152 45902 11204 45908
rect 10600 45348 10652 45354
rect 10600 45290 10652 45296
rect 10416 45008 10468 45014
rect 10416 44950 10468 44956
rect 10784 44736 10836 44742
rect 10784 44678 10836 44684
rect 10796 44470 10824 44678
rect 10784 44464 10836 44470
rect 10784 44406 10836 44412
rect 10232 44396 10284 44402
rect 10232 44338 10284 44344
rect 10244 43761 10272 44338
rect 10796 44198 10824 44406
rect 10784 44192 10836 44198
rect 10784 44134 10836 44140
rect 10230 43752 10286 43761
rect 10230 43687 10286 43696
rect 10244 43654 10272 43687
rect 10232 43648 10284 43654
rect 10232 43590 10284 43596
rect 9680 43444 9732 43450
rect 9680 43386 9732 43392
rect 10048 43444 10100 43450
rect 10048 43386 10100 43392
rect 8944 43308 8996 43314
rect 8944 43250 8996 43256
rect 10508 43308 10560 43314
rect 10508 43250 10560 43256
rect 8956 42906 8984 43250
rect 9220 43104 9272 43110
rect 9220 43046 9272 43052
rect 8944 42900 8996 42906
rect 8944 42842 8996 42848
rect 9232 42838 9260 43046
rect 10520 42906 10548 43250
rect 10508 42900 10560 42906
rect 10508 42842 10560 42848
rect 9220 42832 9272 42838
rect 9220 42774 9272 42780
rect 9128 42696 9180 42702
rect 9128 42638 9180 42644
rect 9140 42294 9168 42638
rect 9128 42288 9180 42294
rect 9128 42230 9180 42236
rect 9232 41614 9260 42774
rect 10508 42696 10560 42702
rect 10508 42638 10560 42644
rect 9680 42560 9732 42566
rect 9680 42502 9732 42508
rect 9692 41750 9720 42502
rect 10520 42362 10548 42638
rect 9956 42356 10008 42362
rect 9956 42298 10008 42304
rect 10140 42356 10192 42362
rect 10140 42298 10192 42304
rect 10508 42356 10560 42362
rect 10508 42298 10560 42304
rect 9680 41744 9732 41750
rect 9680 41686 9732 41692
rect 9220 41608 9272 41614
rect 9220 41550 9272 41556
rect 9968 36378 9996 42298
rect 9956 36372 10008 36378
rect 9956 36314 10008 36320
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 6552 19508 6604 19514
rect 6552 19450 6604 19456
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6472 9722 6500 9862
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5644 7410 5672 8910
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5644 7313 5672 7346
rect 5630 7304 5686 7313
rect 5630 7239 5686 7248
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5538 6760 5594 6769
rect 5538 6695 5594 6704
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5446 6080 5502 6089
rect 5446 6015 5502 6024
rect 5460 5778 5488 6015
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5354 5128 5410 5137
rect 5354 5063 5410 5072
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 3466 5396 4966
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5460 3312 5488 5578
rect 5368 3284 5488 3312
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5172 2916 5224 2922
rect 5172 2858 5224 2864
rect 5170 2816 5226 2825
rect 5170 2751 5226 2760
rect 5184 1358 5212 2751
rect 5172 1352 5224 1358
rect 5172 1294 5224 1300
rect 5170 1184 5226 1193
rect 5170 1119 5226 1128
rect 5184 800 5212 1119
rect 5264 944 5316 950
rect 5264 886 5316 892
rect 5276 800 5304 886
rect 5368 800 5396 3284
rect 5446 3224 5502 3233
rect 5446 3159 5502 3168
rect 5460 800 5488 3159
rect 5552 3058 5580 6598
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5644 2854 5672 7142
rect 5736 6322 5764 9114
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 5710 5764 6054
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5736 3369 5764 5510
rect 5828 4622 5856 8298
rect 5920 6798 5948 8774
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5920 4434 5948 6734
rect 5828 4406 5948 4434
rect 5722 3360 5778 3369
rect 5722 3295 5778 3304
rect 5828 3233 5856 4406
rect 5906 4312 5962 4321
rect 5906 4247 5908 4256
rect 5960 4247 5962 4256
rect 5908 4218 5960 4224
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5814 3224 5870 3233
rect 5814 3159 5870 3168
rect 5722 3088 5778 3097
rect 5920 3058 5948 4082
rect 6012 3516 6040 7346
rect 6104 4729 6132 8230
rect 6196 6730 6224 8774
rect 6380 7410 6408 9318
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6472 7290 6500 9658
rect 8312 9654 8340 12922
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6748 9178 6776 9318
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6288 7262 6500 7290
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 6288 6610 6316 7262
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6196 6582 6316 6610
rect 6196 6118 6224 6582
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6196 5545 6224 5646
rect 6182 5536 6238 5545
rect 6182 5471 6238 5480
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 6090 4720 6146 4729
rect 6090 4655 6146 4664
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6104 3618 6132 4558
rect 6196 3738 6224 5102
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6104 3590 6224 3618
rect 6012 3488 6132 3516
rect 5998 3360 6054 3369
rect 5998 3295 6054 3304
rect 5722 3023 5778 3032
rect 5908 3052 5960 3058
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5736 2666 5764 3023
rect 5908 2994 5960 3000
rect 6012 2904 6040 3295
rect 5552 2638 5764 2666
rect 5920 2876 6040 2904
rect 5552 800 5580 2638
rect 5814 2544 5870 2553
rect 5814 2479 5870 2488
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 5644 1766 5672 2314
rect 5632 1760 5684 1766
rect 5632 1702 5684 1708
rect 5828 1170 5856 2479
rect 5920 2038 5948 2876
rect 5998 2816 6054 2825
rect 5998 2751 6054 2760
rect 5908 2032 5960 2038
rect 5908 1974 5960 1980
rect 5736 1142 5856 1170
rect 5908 1216 5960 1222
rect 5908 1158 5960 1164
rect 5630 912 5686 921
rect 5630 847 5686 856
rect 5644 800 5672 847
rect 5736 800 5764 1142
rect 5920 800 5948 1158
rect 6012 800 6040 2751
rect 6104 800 6132 3488
rect 6196 800 6224 3590
rect 6288 800 6316 6054
rect 6380 3126 6408 7142
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6472 2990 6500 6598
rect 6564 4214 6592 7754
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6380 2446 6408 2790
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6366 2272 6422 2281
rect 6366 2207 6422 2216
rect 6380 800 6408 2207
rect 6472 800 6500 2790
rect 6564 800 6592 4014
rect 6656 3602 6684 7686
rect 6748 5846 6776 9114
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6840 5710 6868 7482
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6828 5704 6880 5710
rect 6748 5664 6828 5692
rect 6748 5137 6776 5664
rect 6828 5646 6880 5652
rect 6932 5522 6960 7142
rect 7024 6322 7052 9386
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7208 7410 7236 8774
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7208 7313 7236 7346
rect 7194 7304 7250 7313
rect 7194 7239 7250 7248
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 6840 5494 6960 5522
rect 6734 5128 6790 5137
rect 6840 5114 6868 5494
rect 6918 5400 6974 5409
rect 6918 5335 6920 5344
rect 6972 5335 6974 5344
rect 6920 5306 6972 5312
rect 6840 5086 6960 5114
rect 6734 5063 6790 5072
rect 6828 5024 6880 5030
rect 6748 4984 6828 5012
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6642 3224 6698 3233
rect 6748 3194 6776 4984
rect 6828 4966 6880 4972
rect 6932 4706 6960 5086
rect 6840 4678 6960 4706
rect 6840 3738 6868 4678
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6642 3159 6698 3168
rect 6736 3188 6788 3194
rect 6656 3058 6684 3159
rect 6736 3130 6788 3136
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6840 2836 6868 3538
rect 6932 2990 6960 4558
rect 7024 4214 7052 6054
rect 7012 4208 7064 4214
rect 7012 4150 7064 4156
rect 7010 4040 7066 4049
rect 7010 3975 7066 3984
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 7024 2854 7052 3975
rect 7116 3534 7144 6598
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7208 2961 7236 6734
rect 7300 6730 7328 8842
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7300 5545 7328 6666
rect 7392 6322 7420 9590
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7378 5944 7434 5953
rect 7378 5879 7380 5888
rect 7432 5879 7434 5888
rect 7380 5850 7432 5856
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7286 5536 7342 5545
rect 7286 5471 7342 5480
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7300 3194 7328 5238
rect 7392 5114 7420 5646
rect 7484 5273 7512 7686
rect 7576 6644 7604 7890
rect 7668 6798 7696 8298
rect 7760 7410 7788 8774
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7576 6616 7696 6644
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7470 5264 7526 5273
rect 7470 5199 7526 5208
rect 7392 5086 7512 5114
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 3534 7420 4966
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7484 3466 7512 5086
rect 7472 3460 7524 3466
rect 7472 3402 7524 3408
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7576 3074 7604 6054
rect 7668 5370 7696 6616
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7300 3046 7604 3074
rect 7194 2952 7250 2961
rect 7104 2916 7156 2922
rect 7194 2887 7250 2896
rect 7104 2858 7156 2864
rect 7012 2848 7064 2854
rect 6840 2808 6960 2836
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6642 2000 6698 2009
rect 6642 1935 6698 1944
rect 6656 800 6684 1935
rect 6748 800 6776 2586
rect 6932 2446 6960 2808
rect 7012 2790 7064 2796
rect 7116 2689 7144 2858
rect 7300 2774 7328 3046
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7208 2746 7328 2774
rect 7102 2680 7158 2689
rect 7102 2615 7158 2624
rect 6920 2440 6972 2446
rect 6826 2408 6882 2417
rect 6920 2382 6972 2388
rect 7010 2408 7066 2417
rect 6826 2343 6882 2352
rect 7010 2343 7012 2352
rect 6840 800 6868 2343
rect 7064 2343 7066 2352
rect 7012 2314 7064 2320
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 6932 1834 6960 2246
rect 6920 1828 6972 1834
rect 6920 1770 6972 1776
rect 7024 1714 7052 2314
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 1766 7144 2246
rect 6932 1686 7052 1714
rect 7104 1760 7156 1766
rect 7104 1702 7156 1708
rect 6932 950 6960 1686
rect 7102 1592 7158 1601
rect 7102 1527 7158 1536
rect 7012 1420 7064 1426
rect 7012 1362 7064 1368
rect 6920 944 6972 950
rect 6920 886 6972 892
rect 7024 800 7052 1362
rect 7116 800 7144 1527
rect 7208 800 7236 2746
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7300 1737 7328 2450
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7286 1728 7342 1737
rect 7286 1663 7342 1672
rect 7288 1624 7340 1630
rect 7288 1566 7340 1572
rect 7300 800 7328 1566
rect 7392 1494 7420 2246
rect 7380 1488 7432 1494
rect 7380 1430 7432 1436
rect 7380 1352 7432 1358
rect 7380 1294 7432 1300
rect 7392 800 7420 1294
rect 7484 800 7512 2926
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7576 2650 7604 2858
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7564 1964 7616 1970
rect 7564 1906 7616 1912
rect 7576 800 7604 1906
rect 7668 800 7696 5170
rect 7760 1426 7788 7346
rect 7852 4622 7880 8366
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7944 7041 7972 7142
rect 7930 7032 7986 7041
rect 7930 6967 7986 6976
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7852 4185 7880 4422
rect 7838 4176 7894 4185
rect 7838 4111 7894 4120
rect 7944 4128 7972 6598
rect 8036 5234 8064 7686
rect 8128 6644 8156 8842
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8220 6798 8248 8230
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8208 6792 8260 6798
rect 8206 6760 8208 6769
rect 8260 6760 8262 6769
rect 8206 6695 8262 6704
rect 8128 6616 8248 6644
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8128 5914 8156 6394
rect 8220 6118 8248 6616
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8206 5944 8262 5953
rect 8116 5908 8168 5914
rect 8206 5879 8208 5888
rect 8116 5850 8168 5856
rect 8260 5879 8262 5888
rect 8208 5850 8260 5856
rect 8312 5760 8340 7142
rect 8404 6322 8432 9454
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8956 8634 8984 8842
rect 9692 8838 9720 8910
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8680 7410 8708 8230
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8220 5732 8340 5760
rect 8116 5704 8168 5710
rect 8220 5692 8248 5732
rect 8168 5664 8248 5692
rect 8116 5646 8168 5652
rect 8116 5568 8168 5574
rect 8300 5568 8352 5574
rect 8116 5510 8168 5516
rect 8220 5516 8300 5522
rect 8220 5510 8352 5516
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8036 4690 8064 5034
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8128 4146 8156 5510
rect 8220 5494 8340 5510
rect 8220 5409 8248 5494
rect 8206 5400 8262 5409
rect 8206 5335 8262 5344
rect 8300 5160 8352 5166
rect 8220 5108 8300 5114
rect 8220 5102 8352 5108
rect 8220 5086 8340 5102
rect 8220 4758 8248 5086
rect 8300 5024 8352 5030
rect 8298 4992 8300 5001
rect 8352 4992 8354 5001
rect 8298 4927 8354 4936
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8300 4684 8352 4690
rect 8404 4672 8432 6054
rect 8496 5370 8524 6326
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8496 5166 8524 5306
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8496 4826 8524 4966
rect 8588 4865 8616 7278
rect 8574 4856 8630 4865
rect 8484 4820 8536 4826
rect 8574 4791 8630 4800
rect 8484 4762 8536 4768
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8352 4644 8432 4672
rect 8300 4626 8352 4632
rect 8206 4584 8262 4593
rect 8482 4584 8538 4593
rect 8262 4542 8340 4570
rect 8206 4519 8262 4528
rect 8206 4176 8262 4185
rect 8116 4140 8168 4146
rect 7944 4100 8064 4128
rect 7930 4040 7986 4049
rect 7930 3975 7986 3984
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7852 2904 7880 3878
rect 7944 3602 7972 3975
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7930 3496 7986 3505
rect 7930 3431 7986 3440
rect 7944 3210 7972 3431
rect 8036 3398 8064 4100
rect 8206 4111 8262 4120
rect 8116 4082 8168 4088
rect 8114 3768 8170 3777
rect 8114 3703 8170 3712
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 7944 3182 8064 3210
rect 7852 2876 7972 2904
rect 7838 2816 7894 2825
rect 7838 2751 7894 2760
rect 7748 1420 7800 1426
rect 7748 1362 7800 1368
rect 7748 1284 7800 1290
rect 7748 1226 7800 1232
rect 7760 800 7788 1226
rect 7852 800 7880 2751
rect 7944 2650 7972 2876
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 7930 2544 7986 2553
rect 7930 2479 7986 2488
rect 7944 800 7972 2479
rect 8036 1630 8064 3182
rect 8128 2990 8156 3703
rect 8220 3058 8248 4111
rect 8312 3738 8340 4542
rect 8482 4519 8538 4528
rect 8496 4282 8524 4519
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8482 4176 8538 4185
rect 8482 4111 8484 4120
rect 8536 4111 8538 4120
rect 8484 4082 8536 4088
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8404 3942 8432 4014
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8482 3904 8538 3913
rect 8482 3839 8538 3848
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8208 2916 8260 2922
rect 8312 2904 8340 3470
rect 8404 2990 8432 3606
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8260 2876 8340 2904
rect 8208 2858 8260 2864
rect 8496 2836 8524 3839
rect 8404 2808 8524 2836
rect 8298 2680 8354 2689
rect 8298 2615 8354 2624
rect 8312 2530 8340 2615
rect 8220 2502 8340 2530
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8024 1624 8076 1630
rect 8024 1566 8076 1572
rect 8128 1476 8156 2382
rect 8036 1448 8156 1476
rect 8036 800 8064 1448
rect 8220 800 8248 2502
rect 8404 2088 8432 2808
rect 8588 2774 8616 4694
rect 8680 3505 8708 7346
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8772 3670 8800 6802
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 8864 4758 8892 6734
rect 9036 6656 9088 6662
rect 9034 6624 9036 6633
rect 9128 6656 9180 6662
rect 9088 6624 9090 6633
rect 9128 6598 9180 6604
rect 9034 6559 9090 6568
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 9048 5409 9076 6054
rect 9034 5400 9090 5409
rect 9034 5335 9090 5344
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8956 4826 8984 4966
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 8942 4720 8998 4729
rect 9048 4706 9076 4762
rect 8998 4678 9076 4706
rect 8942 4655 8998 4664
rect 8852 4616 8904 4622
rect 8850 4584 8852 4593
rect 8904 4584 8906 4593
rect 8850 4519 8906 4528
rect 9036 4480 9088 4486
rect 8864 4428 9036 4434
rect 8864 4422 9088 4428
rect 8864 4406 9076 4422
rect 8864 4282 8892 4406
rect 8942 4312 8998 4321
rect 8852 4276 8904 4282
rect 8942 4247 8998 4256
rect 8852 4218 8904 4224
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8852 3664 8904 3670
rect 8852 3606 8904 3612
rect 8666 3496 8722 3505
rect 8864 3448 8892 3606
rect 8956 3534 8984 4247
rect 9034 3632 9090 3641
rect 9034 3567 9036 3576
rect 9088 3567 9090 3576
rect 9036 3538 9088 3544
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8666 3431 8722 3440
rect 8772 3420 8892 3448
rect 8772 3346 8800 3420
rect 8496 2746 8616 2774
rect 8680 3318 8800 3346
rect 8496 2582 8524 2746
rect 8574 2680 8630 2689
rect 8574 2615 8630 2624
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8482 2408 8538 2417
rect 8482 2343 8538 2352
rect 8312 2060 8432 2088
rect 8312 1970 8340 2060
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 8392 1964 8444 1970
rect 8392 1906 8444 1912
rect 8300 1624 8352 1630
rect 8300 1566 8352 1572
rect 8312 800 8340 1566
rect 8404 1426 8432 1906
rect 8392 1420 8444 1426
rect 8392 1362 8444 1368
rect 8392 1148 8444 1154
rect 8392 1090 8444 1096
rect 8404 800 8432 1090
rect 8496 800 8524 2343
rect 8588 800 8616 2615
rect 8680 800 8708 3318
rect 8758 3224 8814 3233
rect 8758 3159 8814 3168
rect 8772 800 8800 3159
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9048 2689 9076 2994
rect 9140 2854 9168 6598
rect 9232 5710 9260 8774
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9324 7410 9352 8230
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9508 6497 9536 7346
rect 9494 6488 9550 6497
rect 9494 6423 9550 6432
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9232 4758 9260 5306
rect 9220 4752 9272 4758
rect 9324 4729 9352 5850
rect 9416 4865 9444 6190
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9402 4856 9458 4865
rect 9402 4791 9458 4800
rect 9508 4758 9536 4966
rect 9496 4752 9548 4758
rect 9220 4694 9272 4700
rect 9310 4720 9366 4729
rect 9496 4694 9548 4700
rect 9310 4655 9366 4664
rect 9600 4604 9628 7686
rect 9692 6322 9720 8774
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9692 4826 9720 5646
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9784 4622 9812 7686
rect 9876 6798 9904 8230
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9876 5001 9904 6734
rect 9862 4992 9918 5001
rect 9862 4927 9918 4936
rect 9232 4576 9628 4604
rect 9772 4616 9824 4622
rect 9232 4321 9260 4576
rect 9772 4558 9824 4564
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9218 4312 9274 4321
rect 9600 4282 9628 4422
rect 9218 4247 9274 4256
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 9404 4140 9456 4146
rect 9588 4140 9640 4146
rect 9456 4100 9588 4128
rect 9404 4082 9456 4088
rect 9588 4082 9640 4088
rect 9416 4010 9444 4082
rect 9692 4078 9720 4422
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9784 4162 9812 4218
rect 9968 4162 9996 36314
rect 10152 12434 10180 42298
rect 10796 35894 10824 44134
rect 11164 43994 11192 45902
rect 11256 45422 11284 46310
rect 11520 45892 11572 45898
rect 11520 45834 11572 45840
rect 11532 45626 11560 45834
rect 11520 45620 11572 45626
rect 11520 45562 11572 45568
rect 11244 45416 11296 45422
rect 11244 45358 11296 45364
rect 11256 44742 11284 45358
rect 11244 44736 11296 44742
rect 11244 44678 11296 44684
rect 11152 43988 11204 43994
rect 11152 43930 11204 43936
rect 11152 36576 11204 36582
rect 11152 36518 11204 36524
rect 11164 36174 11192 36518
rect 11152 36168 11204 36174
rect 11152 36110 11204 36116
rect 10796 35866 10916 35894
rect 10152 12406 10364 12434
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10152 6322 10180 7686
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10244 6798 10272 7210
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10046 5944 10102 5953
rect 10046 5879 10102 5888
rect 10060 5710 10088 5879
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10152 5556 10180 6258
rect 10244 5914 10272 6734
rect 10336 6497 10364 12406
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10428 7410 10456 8230
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10600 6792 10652 6798
rect 10598 6760 10600 6769
rect 10652 6760 10654 6769
rect 10598 6695 10654 6704
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10598 6624 10654 6633
rect 10322 6488 10378 6497
rect 10322 6423 10378 6432
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 9784 4134 9996 4162
rect 10060 5528 10180 5556
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9496 3936 9548 3942
rect 9218 3904 9274 3913
rect 9274 3862 9444 3890
rect 9784 3890 9812 4134
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9496 3878 9548 3884
rect 9218 3839 9274 3848
rect 9416 3777 9444 3862
rect 9402 3768 9458 3777
rect 9312 3732 9364 3738
rect 9402 3703 9458 3712
rect 9312 3674 9364 3680
rect 9324 3176 9352 3674
rect 9508 3482 9536 3878
rect 9692 3862 9812 3890
rect 9692 3754 9720 3862
rect 9232 3148 9352 3176
rect 9416 3454 9536 3482
rect 9600 3726 9720 3754
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9034 2680 9090 2689
rect 9034 2615 9090 2624
rect 9036 2440 9088 2446
rect 9232 2394 9260 3148
rect 9310 3088 9366 3097
rect 9310 3023 9312 3032
rect 9364 3023 9366 3032
rect 9312 2994 9364 3000
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 9036 2382 9088 2388
rect 8942 2000 8998 2009
rect 8942 1935 8998 1944
rect 8852 944 8904 950
rect 8852 886 8904 892
rect 8864 800 8892 886
rect 8956 800 8984 1935
rect 9048 1426 9076 2382
rect 9140 2366 9260 2394
rect 9036 1420 9088 1426
rect 9036 1362 9088 1368
rect 9034 1320 9090 1329
rect 9034 1255 9090 1264
rect 9048 800 9076 1255
rect 9140 800 9168 2366
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9232 1494 9260 2246
rect 9220 1488 9272 1494
rect 9220 1430 9272 1436
rect 9324 1426 9352 2790
rect 9416 2582 9444 3454
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9404 2576 9456 2582
rect 9404 2518 9456 2524
rect 9404 2032 9456 2038
rect 9404 1974 9456 1980
rect 9312 1420 9364 1426
rect 9312 1362 9364 1368
rect 9220 1352 9272 1358
rect 9220 1294 9272 1300
rect 9232 800 9260 1294
rect 9416 800 9444 1974
rect 9508 1630 9536 3334
rect 9600 3194 9628 3726
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9784 3398 9812 3470
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9680 3188 9732 3194
rect 9876 3176 9904 3606
rect 9968 3602 9996 4014
rect 10060 3913 10088 5528
rect 10138 5400 10194 5409
rect 10138 5335 10140 5344
rect 10192 5335 10194 5344
rect 10140 5306 10192 5312
rect 10244 5302 10272 5646
rect 10232 5296 10284 5302
rect 10232 5238 10284 5244
rect 10230 4992 10286 5001
rect 10230 4927 10286 4936
rect 10244 4321 10272 4927
rect 10230 4312 10286 4321
rect 10230 4247 10286 4256
rect 10336 4026 10364 6054
rect 10244 3998 10364 4026
rect 10046 3904 10102 3913
rect 10046 3839 10102 3848
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9732 3148 9904 3176
rect 9680 3130 9732 3136
rect 9586 3088 9642 3097
rect 9586 3023 9642 3032
rect 9496 1624 9548 1630
rect 9496 1566 9548 1572
rect 9496 1420 9548 1426
rect 9496 1362 9548 1368
rect 9508 800 9536 1362
rect 9600 800 9628 3023
rect 9968 2854 9996 3538
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10152 3233 10180 3334
rect 10138 3224 10194 3233
rect 10048 3188 10100 3194
rect 10138 3159 10194 3168
rect 10048 3130 10100 3136
rect 10060 3058 10088 3130
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 9680 2848 9732 2854
rect 9678 2816 9680 2825
rect 9956 2848 10008 2854
rect 9732 2816 9734 2825
rect 9956 2790 10008 2796
rect 9678 2751 9734 2760
rect 10152 2650 10180 2926
rect 10244 2689 10272 3998
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10230 2680 10286 2689
rect 10140 2644 10192 2650
rect 10230 2615 10286 2624
rect 10140 2586 10192 2592
rect 9678 2544 9734 2553
rect 10336 2514 10364 3878
rect 10428 3670 10456 6598
rect 10598 6559 10654 6568
rect 10612 5642 10640 6559
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10600 5296 10652 5302
rect 10600 5238 10652 5244
rect 10612 5166 10640 5238
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10520 3942 10548 5034
rect 10612 4486 10640 5102
rect 10600 4480 10652 4486
rect 10704 4457 10732 7142
rect 10796 6322 10824 7686
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10888 5545 10916 35866
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10980 6186 11008 6802
rect 11072 6390 11100 7482
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 11058 6080 11114 6089
rect 11058 6015 11114 6024
rect 10966 5808 11022 5817
rect 10966 5743 10968 5752
rect 11020 5743 11022 5752
rect 10968 5714 11020 5720
rect 10874 5536 10930 5545
rect 10874 5471 10930 5480
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10600 4422 10652 4428
rect 10690 4448 10746 4457
rect 10690 4383 10746 4392
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10506 3768 10562 3777
rect 10506 3703 10562 3712
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10520 3602 10548 3703
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10612 3482 10640 4218
rect 10704 4214 10732 4383
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10692 4072 10744 4078
rect 10690 4040 10692 4049
rect 10744 4040 10746 4049
rect 10690 3975 10746 3984
rect 10428 3454 10640 3482
rect 9678 2479 9680 2488
rect 9732 2479 9734 2488
rect 9864 2508 9916 2514
rect 9680 2450 9732 2456
rect 9864 2450 9916 2456
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 1698 9720 2246
rect 9680 1692 9732 1698
rect 9680 1634 9732 1640
rect 9772 1352 9824 1358
rect 9772 1294 9824 1300
rect 9680 1080 9732 1086
rect 9680 1022 9732 1028
rect 9692 800 9720 1022
rect 9784 800 9812 1294
rect 9876 800 9904 2450
rect 9954 2408 10010 2417
rect 9954 2343 10010 2352
rect 10048 2372 10100 2378
rect 9968 800 9996 2343
rect 10048 2314 10100 2320
rect 10324 2372 10376 2378
rect 10324 2314 10376 2320
rect 10060 2038 10088 2314
rect 10336 2145 10364 2314
rect 10322 2136 10378 2145
rect 10322 2071 10378 2080
rect 10048 2032 10100 2038
rect 10048 1974 10100 1980
rect 10048 1420 10100 1426
rect 10048 1362 10100 1368
rect 10060 800 10088 1362
rect 10428 1306 10456 3454
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10140 1284 10192 1290
rect 10140 1226 10192 1232
rect 10244 1278 10456 1306
rect 10152 800 10180 1226
rect 10244 800 10272 1278
rect 10324 1216 10376 1222
rect 10324 1158 10376 1164
rect 10336 800 10364 1158
rect 10520 800 10548 3334
rect 10796 3058 10824 4558
rect 10888 3058 10916 5306
rect 11072 5250 11100 6015
rect 10980 5222 11100 5250
rect 10980 4554 11008 5222
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 11072 4690 11100 5102
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 11060 4480 11112 4486
rect 10966 4448 11022 4457
rect 11022 4428 11060 4434
rect 11022 4422 11112 4428
rect 11022 4406 11100 4422
rect 10966 4383 11022 4392
rect 11058 4312 11114 4321
rect 11058 4247 11114 4256
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10612 1426 10640 2994
rect 10876 2848 10928 2854
rect 10782 2816 10838 2825
rect 10876 2790 10928 2796
rect 10782 2751 10838 2760
rect 10796 2446 10824 2751
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10600 1420 10652 1426
rect 10600 1362 10652 1368
rect 10796 1222 10824 2382
rect 10888 2281 10916 2790
rect 10874 2272 10930 2281
rect 10874 2207 10930 2216
rect 10784 1216 10836 1222
rect 10784 1158 10836 1164
rect 10692 1012 10744 1018
rect 10692 954 10744 960
rect 10704 800 10732 954
rect 10980 800 11008 3946
rect 11072 3777 11100 4247
rect 11058 3768 11114 3777
rect 11058 3703 11114 3712
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 11072 3233 11100 3402
rect 11058 3224 11114 3233
rect 11058 3159 11114 3168
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11072 1154 11100 2518
rect 11164 2514 11192 36110
rect 11256 16574 11284 44678
rect 11716 44402 11744 46514
rect 12820 46170 12848 46514
rect 12912 46170 12940 46990
rect 12808 46164 12860 46170
rect 12808 46106 12860 46112
rect 12900 46164 12952 46170
rect 12900 46106 12952 46112
rect 12820 45558 12848 46106
rect 12900 45892 12952 45898
rect 12900 45834 12952 45840
rect 12808 45552 12860 45558
rect 12808 45494 12860 45500
rect 12912 45490 12940 45834
rect 12900 45484 12952 45490
rect 12900 45426 12952 45432
rect 11980 45416 12032 45422
rect 11980 45358 12032 45364
rect 12164 45416 12216 45422
rect 12164 45358 12216 45364
rect 11992 45286 12020 45358
rect 11980 45280 12032 45286
rect 11980 45222 12032 45228
rect 11992 44402 12020 45222
rect 12176 44402 12204 45358
rect 13096 45354 13124 46990
rect 13464 46714 13492 49200
rect 14292 47258 14320 49200
rect 14280 47252 14332 47258
rect 14280 47194 14332 47200
rect 14372 47048 14424 47054
rect 14372 46990 14424 46996
rect 13452 46708 13504 46714
rect 13452 46650 13504 46656
rect 13820 46572 13872 46578
rect 13820 46514 13872 46520
rect 13728 45484 13780 45490
rect 13728 45426 13780 45432
rect 12440 45348 12492 45354
rect 12440 45290 12492 45296
rect 13084 45348 13136 45354
rect 13084 45290 13136 45296
rect 11704 44396 11756 44402
rect 11704 44338 11756 44344
rect 11980 44396 12032 44402
rect 11980 44338 12032 44344
rect 12164 44396 12216 44402
rect 12164 44338 12216 44344
rect 11612 44192 11664 44198
rect 11612 44134 11664 44140
rect 11624 43790 11652 44134
rect 11612 43784 11664 43790
rect 11612 43726 11664 43732
rect 11716 43654 11744 44338
rect 11980 43852 12032 43858
rect 11980 43794 12032 43800
rect 11704 43648 11756 43654
rect 11704 43590 11756 43596
rect 11796 43648 11848 43654
rect 11796 43590 11848 43596
rect 11808 43382 11836 43590
rect 11796 43376 11848 43382
rect 11796 43318 11848 43324
rect 11992 43296 12020 43794
rect 12176 43790 12204 44338
rect 12452 44334 12480 45290
rect 12900 45280 12952 45286
rect 12900 45222 12952 45228
rect 12532 44940 12584 44946
rect 12584 44900 12664 44928
rect 12532 44882 12584 44888
rect 12636 44470 12664 44900
rect 12624 44464 12676 44470
rect 12624 44406 12676 44412
rect 12440 44328 12492 44334
rect 12440 44270 12492 44276
rect 12912 43858 12940 45222
rect 13740 45014 13768 45426
rect 13728 45008 13780 45014
rect 13728 44950 13780 44956
rect 13740 44742 13768 44950
rect 13728 44736 13780 44742
rect 13728 44678 13780 44684
rect 13176 44532 13228 44538
rect 13176 44474 13228 44480
rect 13188 44334 13216 44474
rect 13176 44328 13228 44334
rect 13176 44270 13228 44276
rect 13188 43858 13216 44270
rect 13268 44192 13320 44198
rect 13268 44134 13320 44140
rect 12900 43852 12952 43858
rect 12900 43794 12952 43800
rect 13176 43852 13228 43858
rect 13176 43794 13228 43800
rect 12164 43784 12216 43790
rect 12164 43726 12216 43732
rect 12176 43382 12204 43726
rect 13280 43722 13308 44134
rect 13268 43716 13320 43722
rect 13268 43658 13320 43664
rect 12164 43376 12216 43382
rect 12164 43318 12216 43324
rect 12072 43308 12124 43314
rect 11992 43268 12072 43296
rect 11992 42906 12020 43268
rect 12072 43250 12124 43256
rect 11980 42900 12032 42906
rect 11980 42842 12032 42848
rect 11992 40050 12020 42842
rect 12440 42152 12492 42158
rect 12440 42094 12492 42100
rect 12256 41812 12308 41818
rect 12256 41754 12308 41760
rect 11980 40044 12032 40050
rect 11980 39986 12032 39992
rect 11256 16546 11376 16574
rect 11348 12434 11376 16546
rect 11348 12406 11928 12434
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11348 6798 11376 7686
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11336 6792 11388 6798
rect 11612 6792 11664 6798
rect 11336 6734 11388 6740
rect 11610 6760 11612 6769
rect 11664 6760 11666 6769
rect 11610 6695 11666 6704
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11256 5642 11284 6258
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11348 5302 11376 6122
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11256 3534 11284 4626
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11256 2961 11284 3470
rect 11242 2952 11298 2961
rect 11242 2887 11298 2896
rect 11244 2848 11296 2854
rect 11348 2825 11376 4966
rect 11440 4758 11468 6394
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11426 4176 11482 4185
rect 11426 4111 11482 4120
rect 11440 3602 11468 4111
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11426 3360 11482 3369
rect 11426 3295 11482 3304
rect 11440 3058 11468 3295
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11532 2922 11560 6598
rect 11716 5710 11744 7142
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11612 4752 11664 4758
rect 11612 4694 11664 4700
rect 11520 2916 11572 2922
rect 11520 2858 11572 2864
rect 11244 2790 11296 2796
rect 11334 2816 11390 2825
rect 11152 2508 11204 2514
rect 11152 2450 11204 2456
rect 11060 1148 11112 1154
rect 11060 1090 11112 1096
rect 11256 800 11284 2790
rect 11624 2774 11652 4694
rect 11334 2751 11390 2760
rect 11532 2746 11652 2774
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11348 1426 11376 2382
rect 11336 1420 11388 1426
rect 11336 1362 11388 1368
rect 11532 800 11560 2746
rect 11716 1086 11744 5646
rect 11808 4690 11836 6598
rect 11900 5137 11928 12406
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 11980 7268 12032 7274
rect 12032 7228 12112 7256
rect 11980 7210 12032 7216
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11886 5128 11942 5137
rect 11886 5063 11942 5072
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 3738 11836 3878
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11808 2689 11836 2926
rect 11794 2680 11850 2689
rect 11794 2615 11850 2624
rect 11704 1080 11756 1086
rect 11704 1022 11756 1028
rect 11900 800 11928 4966
rect 11992 4321 12020 5646
rect 11978 4312 12034 4321
rect 11978 4247 12034 4256
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11992 2582 12020 3674
rect 11980 2576 12032 2582
rect 11980 2518 12032 2524
rect 11980 2440 12032 2446
rect 11978 2408 11980 2417
rect 12032 2408 12034 2417
rect 11978 2343 12034 2352
rect 11992 1630 12020 2343
rect 12084 2310 12112 7228
rect 12176 4593 12204 7346
rect 12268 6254 12296 41754
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12268 5817 12296 5850
rect 12254 5808 12310 5817
rect 12452 5778 12480 42094
rect 13280 35894 13308 43658
rect 13360 43648 13412 43654
rect 13360 43590 13412 43596
rect 13636 43648 13688 43654
rect 13636 43590 13688 43596
rect 13372 43314 13400 43590
rect 13648 43382 13676 43590
rect 13636 43376 13688 43382
rect 13636 43318 13688 43324
rect 13360 43308 13412 43314
rect 13360 43250 13412 43256
rect 13280 35866 13400 35894
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12254 5743 12310 5752
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 12162 4584 12218 4593
rect 12162 4519 12218 4528
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12176 3913 12204 4422
rect 12162 3904 12218 3913
rect 12162 3839 12218 3848
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 11980 1624 12032 1630
rect 11980 1566 12032 1572
rect 12176 800 12204 3674
rect 12268 2378 12296 5510
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12360 3194 12388 4966
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12360 2666 12388 2994
rect 12452 2854 12480 4558
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12360 2638 12480 2666
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12256 2372 12308 2378
rect 12256 2314 12308 2320
rect 12360 1902 12388 2382
rect 12348 1896 12400 1902
rect 12348 1838 12400 1844
rect 12452 1748 12480 2638
rect 12544 2446 12572 6054
rect 12820 4690 12848 7210
rect 13280 6798 13308 16186
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12360 1720 12480 1748
rect 12360 1358 12388 1720
rect 12348 1352 12400 1358
rect 12348 1294 12400 1300
rect 12440 1352 12492 1358
rect 12440 1294 12492 1300
rect 12452 800 12480 1294
rect 12636 1018 12664 3538
rect 12728 3097 12756 3878
rect 12806 3768 12862 3777
rect 12806 3703 12862 3712
rect 12820 3505 12848 3703
rect 12806 3496 12862 3505
rect 12806 3431 12862 3440
rect 12714 3088 12770 3097
rect 12714 3023 12770 3032
rect 12912 2553 12940 5510
rect 13004 3194 13032 5510
rect 13096 5234 13124 6054
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13096 4282 13124 5170
rect 13176 5024 13228 5030
rect 13176 4966 13228 4972
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13082 3768 13138 3777
rect 13082 3703 13138 3712
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 12898 2544 12954 2553
rect 12898 2479 12954 2488
rect 12716 2372 12768 2378
rect 12716 2314 12768 2320
rect 12728 1902 12756 2314
rect 12716 1896 12768 1902
rect 12716 1838 12768 1844
rect 12808 1080 12860 1086
rect 12808 1022 12860 1028
rect 12624 1012 12676 1018
rect 12624 954 12676 960
rect 12820 800 12848 1022
rect 13096 800 13124 3703
rect 13188 2417 13216 4966
rect 13280 3534 13308 6734
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13372 3346 13400 35866
rect 13740 12434 13768 44678
rect 13832 43790 13860 46514
rect 14188 46368 14240 46374
rect 14188 46310 14240 46316
rect 14200 45898 14228 46310
rect 14188 45892 14240 45898
rect 14188 45834 14240 45840
rect 14200 44878 14228 45834
rect 14280 45824 14332 45830
rect 14280 45766 14332 45772
rect 14292 45626 14320 45766
rect 14280 45620 14332 45626
rect 14280 45562 14332 45568
rect 14384 45082 14412 46990
rect 14752 46714 14780 49200
rect 15580 47258 15608 49200
rect 15568 47252 15620 47258
rect 15568 47194 15620 47200
rect 15660 47048 15712 47054
rect 15660 46990 15712 46996
rect 15200 46980 15252 46986
rect 15200 46922 15252 46928
rect 14740 46708 14792 46714
rect 14740 46650 14792 46656
rect 15108 46572 15160 46578
rect 15108 46514 15160 46520
rect 15120 45830 15148 46514
rect 15212 45966 15240 46922
rect 15200 45960 15252 45966
rect 15200 45902 15252 45908
rect 14740 45824 14792 45830
rect 14740 45766 14792 45772
rect 15108 45824 15160 45830
rect 15108 45766 15160 45772
rect 14752 45490 14780 45766
rect 14740 45484 14792 45490
rect 14740 45426 14792 45432
rect 15016 45484 15068 45490
rect 15016 45426 15068 45432
rect 14464 45348 14516 45354
rect 14464 45290 14516 45296
rect 14372 45076 14424 45082
rect 14372 45018 14424 45024
rect 14188 44872 14240 44878
rect 14188 44814 14240 44820
rect 14476 44538 14504 45290
rect 14924 44872 14976 44878
rect 14924 44814 14976 44820
rect 14936 44538 14964 44814
rect 15028 44742 15056 45426
rect 15108 45416 15160 45422
rect 15108 45358 15160 45364
rect 15016 44736 15068 44742
rect 15016 44678 15068 44684
rect 14464 44532 14516 44538
rect 14464 44474 14516 44480
rect 14924 44532 14976 44538
rect 14924 44474 14976 44480
rect 13820 43784 13872 43790
rect 13820 43726 13872 43732
rect 13832 43450 13860 43726
rect 13820 43444 13872 43450
rect 13820 43386 13872 43392
rect 14464 42220 14516 42226
rect 14464 42162 14516 42168
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 13556 12406 13768 12434
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13464 3777 13492 3878
rect 13450 3768 13506 3777
rect 13450 3703 13506 3712
rect 13280 3318 13400 3346
rect 13280 3194 13308 3318
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13280 3058 13308 3130
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13174 2408 13230 2417
rect 13174 2343 13230 2352
rect 13280 1562 13308 2994
rect 13556 1834 13584 12406
rect 14016 6390 14044 17206
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13648 4554 13676 5510
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 13832 2774 13860 4558
rect 14016 4214 14044 6326
rect 14384 6254 14412 6938
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14004 4208 14056 4214
rect 14108 4185 14136 4966
rect 14004 4150 14056 4156
rect 14094 4176 14150 4185
rect 14094 4111 14150 4120
rect 14292 3602 14320 5714
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 14384 4758 14412 5578
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14384 3738 14412 3878
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14476 3126 14504 42162
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 14568 6390 14596 19382
rect 15028 16574 15056 44678
rect 15120 43858 15148 45358
rect 15672 45082 15700 46990
rect 15948 46714 15976 49200
rect 16868 47258 16896 49200
rect 16856 47252 16908 47258
rect 16856 47194 16908 47200
rect 17236 46714 17264 49200
rect 18064 47258 18092 49200
rect 18052 47252 18104 47258
rect 18052 47194 18104 47200
rect 17776 47048 17828 47054
rect 17776 46990 17828 46996
rect 18420 47048 18472 47054
rect 18420 46990 18472 46996
rect 15936 46708 15988 46714
rect 15936 46650 15988 46656
rect 17224 46708 17276 46714
rect 17224 46650 17276 46656
rect 15936 46572 15988 46578
rect 15936 46514 15988 46520
rect 16672 46572 16724 46578
rect 16672 46514 16724 46520
rect 15844 45960 15896 45966
rect 15844 45902 15896 45908
rect 15660 45076 15712 45082
rect 15660 45018 15712 45024
rect 15856 44538 15884 45902
rect 15948 45830 15976 46514
rect 16684 46374 16712 46514
rect 16672 46368 16724 46374
rect 16672 46310 16724 46316
rect 16580 45892 16632 45898
rect 16580 45834 16632 45840
rect 15936 45824 15988 45830
rect 15936 45766 15988 45772
rect 15948 45490 15976 45766
rect 16592 45558 16620 45834
rect 16580 45552 16632 45558
rect 16580 45494 16632 45500
rect 15936 45484 15988 45490
rect 15936 45426 15988 45432
rect 16212 45280 16264 45286
rect 16212 45222 16264 45228
rect 16224 44878 16252 45222
rect 16684 45014 16712 46310
rect 17788 46170 17816 46990
rect 17960 46572 18012 46578
rect 17960 46514 18012 46520
rect 17776 46164 17828 46170
rect 17776 46106 17828 46112
rect 17408 45960 17460 45966
rect 17408 45902 17460 45908
rect 17420 45422 17448 45902
rect 17408 45416 17460 45422
rect 17408 45358 17460 45364
rect 17868 45280 17920 45286
rect 17868 45222 17920 45228
rect 16672 45008 16724 45014
rect 16672 44950 16724 44956
rect 17132 45008 17184 45014
rect 17132 44950 17184 44956
rect 16212 44872 16264 44878
rect 16212 44814 16264 44820
rect 16224 44742 16252 44814
rect 16212 44736 16264 44742
rect 16212 44678 16264 44684
rect 16224 44538 16252 44678
rect 15844 44532 15896 44538
rect 15844 44474 15896 44480
rect 16212 44532 16264 44538
rect 16212 44474 16264 44480
rect 15108 43852 15160 43858
rect 15108 43794 15160 43800
rect 15750 43752 15806 43761
rect 15750 43687 15752 43696
rect 15804 43687 15806 43696
rect 15752 43658 15804 43664
rect 15200 43648 15252 43654
rect 15200 43590 15252 43596
rect 15212 43450 15240 43590
rect 15856 43450 15884 44474
rect 15936 44328 15988 44334
rect 15936 44270 15988 44276
rect 15200 43444 15252 43450
rect 15200 43386 15252 43392
rect 15844 43444 15896 43450
rect 15844 43386 15896 43392
rect 15948 41414 15976 44270
rect 16672 43852 16724 43858
rect 16672 43794 16724 43800
rect 16684 43450 16712 43794
rect 17144 43790 17172 44950
rect 17880 44946 17908 45222
rect 17316 44940 17368 44946
rect 17316 44882 17368 44888
rect 17868 44940 17920 44946
rect 17868 44882 17920 44888
rect 17328 44742 17356 44882
rect 17316 44736 17368 44742
rect 17316 44678 17368 44684
rect 17224 44192 17276 44198
rect 17224 44134 17276 44140
rect 17236 43790 17264 44134
rect 16764 43784 16816 43790
rect 17132 43784 17184 43790
rect 16816 43744 17132 43772
rect 16764 43726 16816 43732
rect 17132 43726 17184 43732
rect 17224 43784 17276 43790
rect 17224 43726 17276 43732
rect 16948 43648 17000 43654
rect 16948 43590 17000 43596
rect 16672 43444 16724 43450
rect 16672 43386 16724 43392
rect 16960 43382 16988 43590
rect 16948 43376 17000 43382
rect 16948 43318 17000 43324
rect 17144 42770 17172 43726
rect 17132 42764 17184 42770
rect 17132 42706 17184 42712
rect 15856 41386 15976 41414
rect 15200 40112 15252 40118
rect 15200 40054 15252 40060
rect 15212 36106 15240 40054
rect 15200 36100 15252 36106
rect 15200 36042 15252 36048
rect 15212 31958 15240 36042
rect 15200 31952 15252 31958
rect 15200 31894 15252 31900
rect 15856 16574 15884 41386
rect 17236 30598 17264 43726
rect 17224 30592 17276 30598
rect 17224 30534 17276 30540
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 15028 16546 15148 16574
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14556 6384 14608 6390
rect 14556 6326 14608 6332
rect 14568 5302 14596 6326
rect 14556 5296 14608 5302
rect 14556 5238 14608 5244
rect 14844 4049 14872 7890
rect 14830 4040 14886 4049
rect 14556 4004 14608 4010
rect 14830 3975 14886 3984
rect 14556 3946 14608 3952
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14200 2774 14228 2926
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 13648 2746 13860 2774
rect 13924 2746 14228 2774
rect 13544 1828 13596 1834
rect 13544 1770 13596 1776
rect 13360 1624 13412 1630
rect 13360 1566 13412 1572
rect 13268 1556 13320 1562
rect 13268 1498 13320 1504
rect 13372 800 13400 1566
rect 13648 800 13676 2746
rect 13924 2038 13952 2746
rect 14004 2576 14056 2582
rect 14004 2518 14056 2524
rect 13912 2032 13964 2038
rect 13912 1974 13964 1980
rect 14016 800 14044 2518
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 1970 14228 2246
rect 14188 1964 14240 1970
rect 14188 1906 14240 1912
rect 14292 800 14320 2790
rect 14568 800 14596 3946
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14660 3194 14688 3674
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 14752 3040 14780 3470
rect 14660 3012 14780 3040
rect 14660 1358 14688 3012
rect 14740 2916 14792 2922
rect 14740 2858 14792 2864
rect 14648 1352 14700 1358
rect 14648 1294 14700 1300
rect 14752 1290 14780 2858
rect 14740 1284 14792 1290
rect 14740 1226 14792 1232
rect 14844 800 14872 3606
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14936 1086 14964 2790
rect 15028 1630 15056 3470
rect 15120 1766 15148 16546
rect 15764 16546 15884 16574
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15212 5778 15240 6054
rect 15304 5914 15332 11018
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15396 5574 15424 7822
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15108 1760 15160 1766
rect 15108 1702 15160 1708
rect 15016 1624 15068 1630
rect 15016 1566 15068 1572
rect 14924 1080 14976 1086
rect 14924 1022 14976 1028
rect 15212 800 15240 4558
rect 15396 2514 15424 5510
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15672 2802 15700 5306
rect 15764 4457 15792 16546
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15856 5914 15884 7754
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15750 4448 15806 4457
rect 15750 4383 15806 4392
rect 15856 3058 15884 5850
rect 16132 5370 16160 18362
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16776 5545 16804 7278
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 16762 5536 16818 5545
rect 16762 5471 16818 5480
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16946 4720 17002 4729
rect 16946 4655 16948 4664
rect 17000 4655 17002 4664
rect 16948 4626 17000 4632
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16316 4078 16344 4422
rect 16960 4146 16988 4626
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 17052 4078 17080 6598
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17236 5710 17264 6258
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 17144 4010 17172 4762
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 15488 2774 15700 2802
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 15488 2446 15516 2774
rect 15476 2440 15528 2446
rect 15660 2440 15712 2446
rect 15476 2382 15528 2388
rect 15580 2400 15660 2428
rect 15580 1306 15608 2400
rect 15660 2382 15712 2388
rect 15488 1278 15608 1306
rect 15488 800 15516 1278
rect 15764 800 15792 2858
rect 16040 800 16068 3538
rect 16408 800 16436 3878
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 16672 2576 16724 2582
rect 16672 2518 16724 2524
rect 16684 800 16712 2518
rect 16960 800 16988 3470
rect 17236 800 17264 3878
rect 17328 1426 17356 44678
rect 17408 43784 17460 43790
rect 17408 43726 17460 43732
rect 17498 43752 17554 43761
rect 17420 42702 17448 43726
rect 17498 43687 17500 43696
rect 17552 43687 17554 43696
rect 17500 43658 17552 43664
rect 17972 43450 18000 46514
rect 18432 46170 18460 46990
rect 18524 46714 18552 49200
rect 19352 47258 19380 49200
rect 19720 47818 19748 49200
rect 19720 47790 20024 47818
rect 19340 47252 19392 47258
rect 19340 47194 19392 47200
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19996 46714 20024 47790
rect 20548 47240 20576 49200
rect 20720 47252 20772 47258
rect 20548 47212 20720 47240
rect 20720 47194 20772 47200
rect 20444 47048 20496 47054
rect 20444 46990 20496 46996
rect 20628 47048 20680 47054
rect 20628 46990 20680 46996
rect 20456 46714 20484 46990
rect 18512 46708 18564 46714
rect 18512 46650 18564 46656
rect 19984 46708 20036 46714
rect 19984 46650 20036 46656
rect 20444 46708 20496 46714
rect 20444 46650 20496 46656
rect 18696 46572 18748 46578
rect 18696 46514 18748 46520
rect 19984 46572 20036 46578
rect 19984 46514 20036 46520
rect 18420 46164 18472 46170
rect 18420 46106 18472 46112
rect 18604 45484 18656 45490
rect 18604 45426 18656 45432
rect 18328 45416 18380 45422
rect 18328 45358 18380 45364
rect 18340 45082 18368 45358
rect 18328 45076 18380 45082
rect 18328 45018 18380 45024
rect 18616 45014 18644 45426
rect 18604 45008 18656 45014
rect 18604 44950 18656 44956
rect 18052 44872 18104 44878
rect 18052 44814 18104 44820
rect 18328 44872 18380 44878
rect 18328 44814 18380 44820
rect 18064 43790 18092 44814
rect 18340 44538 18368 44814
rect 18328 44532 18380 44538
rect 18328 44474 18380 44480
rect 18340 43858 18368 44474
rect 18328 43852 18380 43858
rect 18328 43794 18380 43800
rect 18604 43852 18656 43858
rect 18604 43794 18656 43800
rect 18052 43784 18104 43790
rect 18052 43726 18104 43732
rect 17960 43444 18012 43450
rect 17960 43386 18012 43392
rect 17408 42696 17460 42702
rect 17408 42638 17460 42644
rect 18340 42634 18368 43794
rect 18616 43314 18644 43794
rect 18708 43450 18736 46514
rect 19432 45892 19484 45898
rect 19432 45834 19484 45840
rect 19444 45354 19472 45834
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19432 45348 19484 45354
rect 19432 45290 19484 45296
rect 19996 45286 20024 46514
rect 20640 46170 20668 46990
rect 21008 46714 21036 49200
rect 21836 48090 21864 49200
rect 21836 48062 22140 48090
rect 22112 47258 22140 48062
rect 22100 47252 22152 47258
rect 22100 47194 22152 47200
rect 21916 47048 21968 47054
rect 21916 46990 21968 46996
rect 20996 46708 21048 46714
rect 20996 46650 21048 46656
rect 20720 46572 20772 46578
rect 20720 46514 20772 46520
rect 21088 46572 21140 46578
rect 21088 46514 21140 46520
rect 20628 46164 20680 46170
rect 20628 46106 20680 46112
rect 20732 45966 20760 46514
rect 20720 45960 20772 45966
rect 20720 45902 20772 45908
rect 20720 45348 20772 45354
rect 20720 45290 20772 45296
rect 19708 45280 19760 45286
rect 19708 45222 19760 45228
rect 19984 45280 20036 45286
rect 19984 45222 20036 45228
rect 18788 45008 18840 45014
rect 18788 44950 18840 44956
rect 18800 44198 18828 44950
rect 19720 44878 19748 45222
rect 20732 45082 20760 45290
rect 20720 45076 20772 45082
rect 20720 45018 20772 45024
rect 19708 44872 19760 44878
rect 19708 44814 19760 44820
rect 20352 44872 20404 44878
rect 20352 44814 20404 44820
rect 19432 44804 19484 44810
rect 19432 44746 19484 44752
rect 19444 44334 19472 44746
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19524 44396 19576 44402
rect 19524 44338 19576 44344
rect 20168 44396 20220 44402
rect 20168 44338 20220 44344
rect 20260 44396 20312 44402
rect 20260 44338 20312 44344
rect 19432 44328 19484 44334
rect 19432 44270 19484 44276
rect 19536 44198 19564 44338
rect 18788 44192 18840 44198
rect 18788 44134 18840 44140
rect 19524 44192 19576 44198
rect 19524 44134 19576 44140
rect 20180 43790 20208 44338
rect 20272 43790 20300 44338
rect 20168 43784 20220 43790
rect 20168 43726 20220 43732
rect 20260 43784 20312 43790
rect 20260 43726 20312 43732
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 18696 43444 18748 43450
rect 18696 43386 18748 43392
rect 18604 43308 18656 43314
rect 18604 43250 18656 43256
rect 18708 42702 18736 43386
rect 20180 43314 20208 43726
rect 19340 43308 19392 43314
rect 19340 43250 19392 43256
rect 20168 43308 20220 43314
rect 20168 43250 20220 43256
rect 19352 42770 19380 43250
rect 20364 43178 20392 44814
rect 20904 44804 20956 44810
rect 20904 44746 20956 44752
rect 20916 44538 20944 44746
rect 20996 44736 21048 44742
rect 20996 44678 21048 44684
rect 21008 44538 21036 44678
rect 20536 44532 20588 44538
rect 20536 44474 20588 44480
rect 20904 44532 20956 44538
rect 20904 44474 20956 44480
rect 20996 44532 21048 44538
rect 20996 44474 21048 44480
rect 20548 44334 20576 44474
rect 20536 44328 20588 44334
rect 20588 44288 20668 44316
rect 20536 44270 20588 44276
rect 20640 43382 20668 44288
rect 20628 43376 20680 43382
rect 20628 43318 20680 43324
rect 21100 43314 21128 46514
rect 21928 46170 21956 46990
rect 22204 46714 22232 49200
rect 23032 47258 23060 49200
rect 23020 47252 23072 47258
rect 23020 47194 23072 47200
rect 23112 47048 23164 47054
rect 23112 46990 23164 46996
rect 22192 46708 22244 46714
rect 22192 46650 22244 46656
rect 22560 46572 22612 46578
rect 22560 46514 22612 46520
rect 23020 46572 23072 46578
rect 23020 46514 23072 46520
rect 21916 46164 21968 46170
rect 21916 46106 21968 46112
rect 21548 45960 21600 45966
rect 21548 45902 21600 45908
rect 21560 45354 21588 45902
rect 21548 45348 21600 45354
rect 21548 45290 21600 45296
rect 21560 44946 21588 45290
rect 22572 45082 22600 46514
rect 22744 45892 22796 45898
rect 22744 45834 22796 45840
rect 22756 45626 22784 45834
rect 22744 45620 22796 45626
rect 22744 45562 22796 45568
rect 23032 45490 23060 46514
rect 23020 45484 23072 45490
rect 23020 45426 23072 45432
rect 22100 45076 22152 45082
rect 22100 45018 22152 45024
rect 22560 45076 22612 45082
rect 22560 45018 22612 45024
rect 21548 44940 21600 44946
rect 21548 44882 21600 44888
rect 22112 44402 22140 45018
rect 22100 44396 22152 44402
rect 22100 44338 22152 44344
rect 22284 44396 22336 44402
rect 22284 44338 22336 44344
rect 21272 44328 21324 44334
rect 21272 44270 21324 44276
rect 22192 44328 22244 44334
rect 22192 44270 22244 44276
rect 21284 43858 21312 44270
rect 22008 44192 22060 44198
rect 22204 44180 22232 44270
rect 22060 44152 22232 44180
rect 22008 44134 22060 44140
rect 21180 43852 21232 43858
rect 21180 43794 21232 43800
rect 21272 43852 21324 43858
rect 21272 43794 21324 43800
rect 21192 43314 21220 43794
rect 21284 43654 21312 43794
rect 22192 43784 22244 43790
rect 22192 43726 22244 43732
rect 21272 43648 21324 43654
rect 21272 43590 21324 43596
rect 20536 43308 20588 43314
rect 21088 43308 21140 43314
rect 20536 43250 20588 43256
rect 21008 43268 21088 43296
rect 20352 43172 20404 43178
rect 20352 43114 20404 43120
rect 19616 43104 19668 43110
rect 19616 43046 19668 43052
rect 19628 42770 19656 43046
rect 19340 42764 19392 42770
rect 19340 42706 19392 42712
rect 19616 42764 19668 42770
rect 19616 42706 19668 42712
rect 18696 42696 18748 42702
rect 18696 42638 18748 42644
rect 18328 42628 18380 42634
rect 18328 42570 18380 42576
rect 18512 42560 18564 42566
rect 18512 42502 18564 42508
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17774 2680 17830 2689
rect 17774 2615 17830 2624
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 17420 1902 17448 2314
rect 17408 1896 17460 1902
rect 17408 1838 17460 1844
rect 17316 1420 17368 1426
rect 17316 1362 17368 1368
rect 17604 800 17632 2382
rect 17788 2310 17816 2615
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17880 800 17908 3470
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 18156 800 18184 2858
rect 18432 800 18460 3878
rect 18524 3126 18552 42502
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 20548 42294 20576 43250
rect 20628 43240 20680 43246
rect 20628 43182 20680 43188
rect 20640 42906 20668 43182
rect 21008 42906 21036 43268
rect 21088 43250 21140 43256
rect 21180 43308 21232 43314
rect 21180 43250 21232 43256
rect 21916 43308 21968 43314
rect 21916 43250 21968 43256
rect 21088 43104 21140 43110
rect 21088 43046 21140 43052
rect 21364 43104 21416 43110
rect 21364 43046 21416 43052
rect 20628 42900 20680 42906
rect 20628 42842 20680 42848
rect 20996 42900 21048 42906
rect 20996 42842 21048 42848
rect 21100 42702 21128 43046
rect 21088 42696 21140 42702
rect 21088 42638 21140 42644
rect 20076 42288 20128 42294
rect 20076 42230 20128 42236
rect 20536 42288 20588 42294
rect 20536 42230 20588 42236
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 18604 40724 18656 40730
rect 18604 40666 18656 40672
rect 18616 5953 18644 40666
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19892 32428 19944 32434
rect 19892 32370 19944 32376
rect 19904 31822 19932 32370
rect 19892 31816 19944 31822
rect 19944 31764 20024 31770
rect 19892 31758 20024 31764
rect 19904 31742 20024 31758
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19996 25362 20024 31742
rect 19984 25356 20036 25362
rect 19984 25298 20036 25304
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 20088 16574 20116 42230
rect 20088 16546 20208 16574
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 18602 5944 18658 5953
rect 18602 5879 18658 5888
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 20180 4146 20208 16546
rect 21376 5166 21404 43046
rect 21928 42770 21956 43250
rect 21916 42764 21968 42770
rect 21916 42706 21968 42712
rect 22204 16574 22232 43726
rect 22296 43722 22324 44338
rect 22928 43784 22980 43790
rect 22926 43752 22928 43761
rect 22980 43752 22982 43761
rect 22284 43716 22336 43722
rect 22926 43687 22982 43696
rect 22284 43658 22336 43664
rect 22204 16546 22324 16574
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 19064 3528 19116 3534
rect 19064 3470 19116 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 18512 3120 18564 3126
rect 18512 3062 18564 3068
rect 18524 2774 18552 3062
rect 18524 2746 18644 2774
rect 18616 2446 18644 2746
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 18616 1494 18644 2382
rect 18604 1488 18656 1494
rect 18604 1430 18656 1436
rect 18800 800 18828 2382
rect 19076 800 19104 3470
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19352 800 19380 2382
rect 19444 1442 19472 3470
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 20180 3126 20208 4082
rect 20364 3194 20392 4082
rect 22296 4010 22324 16546
rect 23032 6458 23060 45426
rect 23124 45082 23152 46990
rect 23492 46714 23520 49200
rect 24320 47258 24348 49200
rect 24308 47252 24360 47258
rect 24308 47194 24360 47200
rect 24400 47048 24452 47054
rect 24400 46990 24452 46996
rect 23480 46708 23532 46714
rect 23480 46650 23532 46656
rect 23756 46572 23808 46578
rect 23756 46514 23808 46520
rect 23768 45830 23796 46514
rect 23756 45824 23808 45830
rect 23756 45766 23808 45772
rect 23768 45558 23796 45766
rect 23756 45552 23808 45558
rect 23756 45494 23808 45500
rect 23940 45552 23992 45558
rect 23940 45494 23992 45500
rect 23848 45484 23900 45490
rect 23848 45426 23900 45432
rect 23664 45416 23716 45422
rect 23664 45358 23716 45364
rect 23112 45076 23164 45082
rect 23112 45018 23164 45024
rect 23572 44804 23624 44810
rect 23572 44746 23624 44752
rect 23584 44402 23612 44746
rect 23572 44396 23624 44402
rect 23572 44338 23624 44344
rect 23480 44328 23532 44334
rect 23676 44282 23704 45358
rect 23756 45348 23808 45354
rect 23756 45290 23808 45296
rect 23768 44402 23796 45290
rect 23756 44396 23808 44402
rect 23756 44338 23808 44344
rect 23480 44270 23532 44276
rect 23492 44198 23520 44270
rect 23584 44254 23704 44282
rect 23480 44192 23532 44198
rect 23480 44134 23532 44140
rect 23584 43790 23612 44254
rect 23664 44192 23716 44198
rect 23664 44134 23716 44140
rect 23572 43784 23624 43790
rect 23386 43752 23442 43761
rect 23124 43710 23336 43738
rect 23124 43450 23152 43710
rect 23308 43654 23336 43710
rect 23572 43726 23624 43732
rect 23386 43687 23442 43696
rect 23204 43648 23256 43654
rect 23204 43590 23256 43596
rect 23296 43648 23348 43654
rect 23296 43590 23348 43596
rect 23112 43444 23164 43450
rect 23112 43386 23164 43392
rect 23216 43314 23244 43590
rect 23400 43450 23428 43687
rect 23388 43444 23440 43450
rect 23388 43386 23440 43392
rect 23296 43376 23348 43382
rect 23296 43318 23348 43324
rect 23204 43308 23256 43314
rect 23204 43250 23256 43256
rect 23308 42906 23336 43318
rect 23296 42900 23348 42906
rect 23296 42842 23348 42848
rect 23388 42628 23440 42634
rect 23388 42570 23440 42576
rect 23400 38282 23428 42570
rect 23584 42566 23612 43726
rect 23572 42560 23624 42566
rect 23572 42502 23624 42508
rect 23388 38276 23440 38282
rect 23388 38218 23440 38224
rect 23400 32502 23428 38218
rect 23388 32496 23440 32502
rect 23388 32438 23440 32444
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23676 6322 23704 44134
rect 23860 43790 23888 45426
rect 23952 44742 23980 45494
rect 24412 44742 24440 46990
rect 24688 46714 24716 49200
rect 25608 47258 25636 49200
rect 25596 47252 25648 47258
rect 25596 47194 25648 47200
rect 25688 47048 25740 47054
rect 25688 46990 25740 46996
rect 24676 46708 24728 46714
rect 24676 46650 24728 46656
rect 24952 46572 25004 46578
rect 24952 46514 25004 46520
rect 24768 46368 24820 46374
rect 24768 46310 24820 46316
rect 24584 45076 24636 45082
rect 24584 45018 24636 45024
rect 24596 44878 24624 45018
rect 24780 45014 24808 46310
rect 24860 45960 24912 45966
rect 24860 45902 24912 45908
rect 24768 45008 24820 45014
rect 24768 44950 24820 44956
rect 24584 44872 24636 44878
rect 24584 44814 24636 44820
rect 23940 44736 23992 44742
rect 23940 44678 23992 44684
rect 24400 44736 24452 44742
rect 24400 44678 24452 44684
rect 23952 44198 23980 44678
rect 24872 44402 24900 45902
rect 24768 44396 24820 44402
rect 24768 44338 24820 44344
rect 24860 44396 24912 44402
rect 24860 44338 24912 44344
rect 24676 44328 24728 44334
rect 24676 44270 24728 44276
rect 23940 44192 23992 44198
rect 23940 44134 23992 44140
rect 24584 44192 24636 44198
rect 24584 44134 24636 44140
rect 24596 43790 24624 44134
rect 24688 43790 24716 44270
rect 24780 43858 24808 44338
rect 24768 43852 24820 43858
rect 24768 43794 24820 43800
rect 23756 43784 23808 43790
rect 23756 43726 23808 43732
rect 23848 43784 23900 43790
rect 23848 43726 23900 43732
rect 24584 43784 24636 43790
rect 24584 43726 24636 43732
rect 24676 43784 24728 43790
rect 24676 43726 24728 43732
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20168 3120 20220 3126
rect 20168 3062 20220 3068
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19444 1414 19656 1442
rect 19628 800 19656 1414
rect 19996 800 20024 2858
rect 20180 1698 20208 3062
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20168 1692 20220 1698
rect 20168 1634 20220 1640
rect 20272 800 20300 2382
rect 20548 800 20576 3470
rect 20824 800 20852 3470
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 21192 800 21220 2382
rect 21468 800 21496 3470
rect 22296 3126 22324 3946
rect 23768 3670 23796 43726
rect 23860 42702 23888 43726
rect 23848 42696 23900 42702
rect 23848 42638 23900 42644
rect 24216 42628 24268 42634
rect 24216 42570 24268 42576
rect 24228 42022 24256 42570
rect 24216 42016 24268 42022
rect 24216 41958 24268 41964
rect 24228 36582 24256 41958
rect 24596 41478 24624 43726
rect 24780 42770 24808 43794
rect 24872 43382 24900 44338
rect 24964 43450 24992 46514
rect 25136 45892 25188 45898
rect 25136 45834 25188 45840
rect 25148 45626 25176 45834
rect 25136 45620 25188 45626
rect 25136 45562 25188 45568
rect 25700 45354 25728 46990
rect 25976 46714 26004 49200
rect 26804 47258 26832 49200
rect 26792 47252 26844 47258
rect 26792 47194 26844 47200
rect 26976 47048 27028 47054
rect 26976 46990 27028 46996
rect 25964 46708 26016 46714
rect 25964 46650 26016 46656
rect 26240 46572 26292 46578
rect 26240 46514 26292 46520
rect 26252 45830 26280 46514
rect 26988 46170 27016 46990
rect 27264 46714 27292 49200
rect 28092 47258 28120 49200
rect 28080 47252 28132 47258
rect 28080 47194 28132 47200
rect 28172 47048 28224 47054
rect 28172 46990 28224 46996
rect 27252 46708 27304 46714
rect 27252 46650 27304 46656
rect 27436 46572 27488 46578
rect 27436 46514 27488 46520
rect 27528 46572 27580 46578
rect 27528 46514 27580 46520
rect 26976 46164 27028 46170
rect 26976 46106 27028 46112
rect 26976 45960 27028 45966
rect 26976 45902 27028 45908
rect 26424 45892 26476 45898
rect 26424 45834 26476 45840
rect 26240 45824 26292 45830
rect 26240 45766 26292 45772
rect 26252 45558 26280 45766
rect 26240 45552 26292 45558
rect 26240 45494 26292 45500
rect 26332 45484 26384 45490
rect 26332 45426 26384 45432
rect 25688 45348 25740 45354
rect 25688 45290 25740 45296
rect 26344 45286 26372 45426
rect 26332 45280 26384 45286
rect 26332 45222 26384 45228
rect 25136 44396 25188 44402
rect 25136 44338 25188 44344
rect 25148 43858 25176 44338
rect 26436 44198 26464 45834
rect 26988 45286 27016 45902
rect 27448 45422 27476 46514
rect 27436 45416 27488 45422
rect 27436 45358 27488 45364
rect 26976 45280 27028 45286
rect 26976 45222 27028 45228
rect 26988 45082 27016 45222
rect 26976 45076 27028 45082
rect 26976 45018 27028 45024
rect 27344 44804 27396 44810
rect 27344 44746 27396 44752
rect 27356 44402 27384 44746
rect 27344 44396 27396 44402
rect 27344 44338 27396 44344
rect 26424 44192 26476 44198
rect 26424 44134 26476 44140
rect 25136 43852 25188 43858
rect 25136 43794 25188 43800
rect 26436 43790 26464 44134
rect 27356 43858 27384 44338
rect 27344 43852 27396 43858
rect 27344 43794 27396 43800
rect 26424 43784 26476 43790
rect 26424 43726 26476 43732
rect 27540 43450 27568 46514
rect 28184 46170 28212 46990
rect 28460 46170 28488 49200
rect 29288 47258 29316 49200
rect 29276 47252 29328 47258
rect 29276 47194 29328 47200
rect 29552 47048 29604 47054
rect 29552 46990 29604 46996
rect 28816 46912 28868 46918
rect 28816 46854 28868 46860
rect 28828 46578 28856 46854
rect 28816 46572 28868 46578
rect 28816 46514 28868 46520
rect 28172 46164 28224 46170
rect 28172 46106 28224 46112
rect 28448 46164 28500 46170
rect 28448 46106 28500 46112
rect 28448 45620 28500 45626
rect 28448 45562 28500 45568
rect 28264 45484 28316 45490
rect 28264 45426 28316 45432
rect 27988 45416 28040 45422
rect 27988 45358 28040 45364
rect 24952 43444 25004 43450
rect 24952 43386 25004 43392
rect 26332 43444 26384 43450
rect 26332 43386 26384 43392
rect 27528 43444 27580 43450
rect 27528 43386 27580 43392
rect 24860 43376 24912 43382
rect 24860 43318 24912 43324
rect 25228 43308 25280 43314
rect 25228 43250 25280 43256
rect 25240 42906 25268 43250
rect 25228 42900 25280 42906
rect 25228 42842 25280 42848
rect 24768 42764 24820 42770
rect 24768 42706 24820 42712
rect 26344 42702 26372 43386
rect 28000 43246 28028 45358
rect 28276 45082 28304 45426
rect 28264 45076 28316 45082
rect 28264 45018 28316 45024
rect 28356 45076 28408 45082
rect 28356 45018 28408 45024
rect 28368 44946 28396 45018
rect 28356 44940 28408 44946
rect 28356 44882 28408 44888
rect 28460 44878 28488 45562
rect 28540 45552 28592 45558
rect 28540 45494 28592 45500
rect 28552 44962 28580 45494
rect 28828 45082 28856 46514
rect 29000 46368 29052 46374
rect 29000 46310 29052 46316
rect 29012 46102 29040 46310
rect 29564 46170 29592 46990
rect 29748 46714 29776 49200
rect 30576 47258 30604 49200
rect 30564 47252 30616 47258
rect 30564 47194 30616 47200
rect 30656 47048 30708 47054
rect 30656 46990 30708 46996
rect 29736 46708 29788 46714
rect 29736 46650 29788 46656
rect 29828 46572 29880 46578
rect 29828 46514 29880 46520
rect 29552 46164 29604 46170
rect 29552 46106 29604 46112
rect 29000 46096 29052 46102
rect 29000 46038 29052 46044
rect 29736 45960 29788 45966
rect 29736 45902 29788 45908
rect 29748 45830 29776 45902
rect 29736 45824 29788 45830
rect 29736 45766 29788 45772
rect 29000 45484 29052 45490
rect 29000 45426 29052 45432
rect 28816 45076 28868 45082
rect 28816 45018 28868 45024
rect 28552 44946 28764 44962
rect 28540 44940 28764 44946
rect 28592 44934 28764 44940
rect 28540 44882 28592 44888
rect 28448 44872 28500 44878
rect 28448 44814 28500 44820
rect 28540 44736 28592 44742
rect 28540 44678 28592 44684
rect 28080 44328 28132 44334
rect 28080 44270 28132 44276
rect 28092 44198 28120 44270
rect 28080 44192 28132 44198
rect 28080 44134 28132 44140
rect 28092 43654 28120 44134
rect 28552 43722 28580 44678
rect 28736 44470 28764 44934
rect 28828 44878 28856 45018
rect 29012 44878 29040 45426
rect 28816 44872 28868 44878
rect 28816 44814 28868 44820
rect 29000 44872 29052 44878
rect 29000 44814 29052 44820
rect 28908 44804 28960 44810
rect 28908 44746 28960 44752
rect 28724 44464 28776 44470
rect 28724 44406 28776 44412
rect 28736 44180 28764 44406
rect 28644 44152 28764 44180
rect 28644 43790 28672 44152
rect 28632 43784 28684 43790
rect 28632 43726 28684 43732
rect 28540 43716 28592 43722
rect 28540 43658 28592 43664
rect 28080 43648 28132 43654
rect 28080 43590 28132 43596
rect 28264 43648 28316 43654
rect 28264 43590 28316 43596
rect 28276 43382 28304 43590
rect 28264 43376 28316 43382
rect 28264 43318 28316 43324
rect 28920 43314 28948 44746
rect 29012 44334 29040 44814
rect 29748 44810 29776 45766
rect 29736 44804 29788 44810
rect 29736 44746 29788 44752
rect 29090 44432 29146 44441
rect 29090 44367 29092 44376
rect 29144 44367 29146 44376
rect 29092 44338 29144 44344
rect 29000 44328 29052 44334
rect 29000 44270 29052 44276
rect 29012 43790 29040 44270
rect 29000 43784 29052 43790
rect 29000 43726 29052 43732
rect 29276 43648 29328 43654
rect 29276 43590 29328 43596
rect 28908 43308 28960 43314
rect 28908 43250 28960 43256
rect 27988 43240 28040 43246
rect 27988 43182 28040 43188
rect 26332 42696 26384 42702
rect 26332 42638 26384 42644
rect 26792 42696 26844 42702
rect 26792 42638 26844 42644
rect 26804 42362 26832 42638
rect 26792 42356 26844 42362
rect 26792 42298 26844 42304
rect 28000 42226 28028 43182
rect 27988 42220 28040 42226
rect 27988 42162 28040 42168
rect 24584 41472 24636 41478
rect 24584 41414 24636 41420
rect 28000 38486 28028 42162
rect 27988 38480 28040 38486
rect 27988 38422 28040 38428
rect 24216 36576 24268 36582
rect 24216 36518 24268 36524
rect 28540 25152 28592 25158
rect 28540 25094 28592 25100
rect 27344 14340 27396 14346
rect 27344 14282 27396 14288
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 25240 5234 25268 11834
rect 27356 9518 27384 14282
rect 27344 9512 27396 9518
rect 27344 9454 27396 9460
rect 25228 5228 25280 5234
rect 25228 5170 25280 5176
rect 27988 3936 28040 3942
rect 27988 3878 28040 3884
rect 23756 3664 23808 3670
rect 23754 3632 23756 3641
rect 23808 3632 23810 3641
rect 23754 3567 23810 3576
rect 22376 3528 22428 3534
rect 22376 3470 22428 3476
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 22284 3120 22336 3126
rect 22284 3062 22336 3068
rect 21732 2916 21784 2922
rect 21732 2858 21784 2864
rect 21744 800 21772 2858
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22112 800 22140 2382
rect 22388 800 22416 3470
rect 22928 2508 22980 2514
rect 22928 2450 22980 2456
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22664 800 22692 2382
rect 22940 800 22968 2450
rect 23308 800 23336 3470
rect 23768 3058 23796 3567
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 25044 3528 25096 3534
rect 25044 3470 25096 3476
rect 25964 3528 26016 3534
rect 25964 3470 26016 3476
rect 26240 3528 26292 3534
rect 26240 3470 26292 3476
rect 27436 3528 27488 3534
rect 27436 3470 27488 3476
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 23572 2916 23624 2922
rect 23572 2858 23624 2864
rect 23584 800 23612 2858
rect 23848 2576 23900 2582
rect 23848 2518 23900 2524
rect 23860 800 23888 2518
rect 24136 800 24164 3470
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24228 3194 24256 3334
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 24504 800 24532 2926
rect 24768 2508 24820 2514
rect 24768 2450 24820 2456
rect 24780 800 24808 2450
rect 25056 800 25084 3470
rect 25320 2916 25372 2922
rect 25320 2858 25372 2864
rect 25332 800 25360 2858
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 25792 1306 25820 2382
rect 25700 1278 25820 1306
rect 25700 800 25728 1278
rect 25976 800 26004 3470
rect 26252 800 26280 3470
rect 26516 2848 26568 2854
rect 26516 2790 26568 2796
rect 27160 2848 27212 2854
rect 27160 2790 27212 2796
rect 26528 800 26556 2790
rect 26884 2508 26936 2514
rect 26884 2450 26936 2456
rect 26896 800 26924 2450
rect 27172 800 27200 2790
rect 27448 800 27476 3470
rect 28000 3126 28028 3878
rect 28080 3528 28132 3534
rect 28080 3470 28132 3476
rect 28356 3528 28408 3534
rect 28356 3470 28408 3476
rect 27988 3120 28040 3126
rect 27988 3062 28040 3068
rect 28000 2774 28028 3062
rect 27908 2746 28028 2774
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 27724 800 27752 2382
rect 27908 2106 27936 2746
rect 27896 2100 27948 2106
rect 27896 2042 27948 2048
rect 28092 800 28120 3470
rect 28368 800 28396 3470
rect 28552 3194 28580 25094
rect 29288 12434 29316 43590
rect 29748 41414 29776 44746
rect 29840 43858 29868 46514
rect 30668 46170 30696 46990
rect 30944 46170 30972 49200
rect 31772 47258 31800 49200
rect 31760 47252 31812 47258
rect 31760 47194 31812 47200
rect 31300 46912 31352 46918
rect 31300 46854 31352 46860
rect 31312 46578 31340 46854
rect 32036 46640 32088 46646
rect 32036 46582 32088 46588
rect 31300 46572 31352 46578
rect 31300 46514 31352 46520
rect 31760 46572 31812 46578
rect 31760 46514 31812 46520
rect 30656 46164 30708 46170
rect 30656 46106 30708 46112
rect 30932 46164 30984 46170
rect 30932 46106 30984 46112
rect 30472 45960 30524 45966
rect 30472 45902 30524 45908
rect 30484 45626 30512 45902
rect 30472 45620 30524 45626
rect 30472 45562 30524 45568
rect 31208 45552 31260 45558
rect 30930 45520 30986 45529
rect 31208 45494 31260 45500
rect 30930 45455 30932 45464
rect 30984 45455 30986 45464
rect 30932 45426 30984 45432
rect 30944 45370 30972 45426
rect 31116 45416 31168 45422
rect 30196 45348 30248 45354
rect 30196 45290 30248 45296
rect 30852 45342 30972 45370
rect 31036 45376 31116 45404
rect 30208 44334 30236 45290
rect 30472 44804 30524 44810
rect 30472 44746 30524 44752
rect 30484 44470 30512 44746
rect 30472 44464 30524 44470
rect 30472 44406 30524 44412
rect 30196 44328 30248 44334
rect 30196 44270 30248 44276
rect 30746 44296 30802 44305
rect 30746 44231 30748 44240
rect 30800 44231 30802 44240
rect 30748 44202 30800 44208
rect 30104 44192 30156 44198
rect 30104 44134 30156 44140
rect 29828 43852 29880 43858
rect 29828 43794 29880 43800
rect 29840 43450 29868 43794
rect 29828 43444 29880 43450
rect 29828 43386 29880 43392
rect 30116 43382 30144 44134
rect 30380 43648 30432 43654
rect 30380 43590 30432 43596
rect 30104 43376 30156 43382
rect 30104 43318 30156 43324
rect 30116 42906 30144 43318
rect 30104 42900 30156 42906
rect 30104 42842 30156 42848
rect 29748 41386 29868 41414
rect 29196 12406 29316 12434
rect 29092 5024 29144 5030
rect 29092 4966 29144 4972
rect 29104 4622 29132 4966
rect 29092 4616 29144 4622
rect 29092 4558 29144 4564
rect 28816 4480 28868 4486
rect 28816 4422 28868 4428
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 28540 3188 28592 3194
rect 28540 3130 28592 3136
rect 28644 800 28672 3878
rect 28828 2990 28856 4422
rect 28908 3936 28960 3942
rect 28908 3878 28960 3884
rect 28816 2984 28868 2990
rect 28816 2926 28868 2932
rect 28920 800 28948 3878
rect 29196 2650 29224 12406
rect 29460 4480 29512 4486
rect 29460 4422 29512 4428
rect 29276 3528 29328 3534
rect 29472 3505 29500 4422
rect 29736 4004 29788 4010
rect 29736 3946 29788 3952
rect 29552 3664 29604 3670
rect 29552 3606 29604 3612
rect 29276 3470 29328 3476
rect 29458 3496 29514 3505
rect 29184 2644 29236 2650
rect 29184 2586 29236 2592
rect 29196 2378 29224 2586
rect 29184 2372 29236 2378
rect 29184 2314 29236 2320
rect 29288 800 29316 3470
rect 29458 3431 29514 3440
rect 29564 800 29592 3606
rect 29748 800 29776 3946
rect 29840 3126 29868 41386
rect 30392 7954 30420 43590
rect 30472 42560 30524 42566
rect 30472 42502 30524 42508
rect 30484 42226 30512 42502
rect 30472 42220 30524 42226
rect 30472 42162 30524 42168
rect 30748 41608 30800 41614
rect 30748 41550 30800 41556
rect 30760 41274 30788 41550
rect 30852 41414 30880 45342
rect 31036 44742 31064 45376
rect 31116 45358 31168 45364
rect 31220 44878 31248 45494
rect 31208 44872 31260 44878
rect 31208 44814 31260 44820
rect 31024 44736 31076 44742
rect 31024 44678 31076 44684
rect 30932 44396 30984 44402
rect 31036 44384 31064 44678
rect 31220 44402 31248 44814
rect 30984 44356 31064 44384
rect 31208 44396 31260 44402
rect 30932 44338 30984 44344
rect 31208 44338 31260 44344
rect 31312 44334 31340 46514
rect 31392 45892 31444 45898
rect 31392 45834 31444 45840
rect 31404 45626 31432 45834
rect 31392 45620 31444 45626
rect 31392 45562 31444 45568
rect 31772 45014 31800 46514
rect 32048 46170 32076 46582
rect 32232 46442 32260 49200
rect 33060 47240 33088 49200
rect 33520 47258 33548 49200
rect 33140 47252 33192 47258
rect 33060 47212 33140 47240
rect 33140 47194 33192 47200
rect 33508 47252 33560 47258
rect 34348 47240 34376 49200
rect 34520 47252 34572 47258
rect 34348 47212 34520 47240
rect 33508 47194 33560 47200
rect 34520 47194 34572 47200
rect 34716 47138 34744 49200
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 35544 47258 35572 49200
rect 35532 47252 35584 47258
rect 35532 47194 35584 47200
rect 34716 47110 34836 47138
rect 32404 47048 32456 47054
rect 32404 46990 32456 46996
rect 33416 47048 33468 47054
rect 33416 46990 33468 46996
rect 34704 47048 34756 47054
rect 34704 46990 34756 46996
rect 32416 46714 32444 46990
rect 33140 46980 33192 46986
rect 33140 46922 33192 46928
rect 32404 46708 32456 46714
rect 32404 46650 32456 46656
rect 32220 46436 32272 46442
rect 32220 46378 32272 46384
rect 32036 46164 32088 46170
rect 32036 46106 32088 46112
rect 31852 46096 31904 46102
rect 31904 46044 32168 46050
rect 31852 46038 32168 46044
rect 31864 46022 32168 46038
rect 31944 45892 31996 45898
rect 31944 45834 31996 45840
rect 31956 45558 31984 45834
rect 32140 45626 32168 46022
rect 33152 45830 33180 46922
rect 33428 46714 33456 46990
rect 34612 46980 34664 46986
rect 34612 46922 34664 46928
rect 33416 46708 33468 46714
rect 33416 46650 33468 46656
rect 34336 46572 34388 46578
rect 34336 46514 34388 46520
rect 34348 45966 34376 46514
rect 33232 45960 33284 45966
rect 33232 45902 33284 45908
rect 33324 45960 33376 45966
rect 33324 45902 33376 45908
rect 34336 45960 34388 45966
rect 34336 45902 34388 45908
rect 33140 45824 33192 45830
rect 33140 45766 33192 45772
rect 32128 45620 32180 45626
rect 32128 45562 32180 45568
rect 31944 45552 31996 45558
rect 31944 45494 31996 45500
rect 33152 45490 33180 45766
rect 33244 45490 33272 45902
rect 33336 45558 33364 45902
rect 33324 45552 33376 45558
rect 33324 45494 33376 45500
rect 33140 45484 33192 45490
rect 33140 45426 33192 45432
rect 33232 45484 33284 45490
rect 33232 45426 33284 45432
rect 33508 45484 33560 45490
rect 33508 45426 33560 45432
rect 33140 45348 33192 45354
rect 33140 45290 33192 45296
rect 31760 45008 31812 45014
rect 31760 44950 31812 44956
rect 31772 44470 31800 44950
rect 33152 44946 33180 45290
rect 33244 45082 33272 45426
rect 33520 45082 33548 45426
rect 34348 45082 34376 45902
rect 34624 45286 34652 46922
rect 34716 46714 34744 46990
rect 34808 46918 34836 47110
rect 35624 47048 35676 47054
rect 35624 46990 35676 46996
rect 34796 46912 34848 46918
rect 34796 46854 34848 46860
rect 34704 46708 34756 46714
rect 34704 46650 34756 46656
rect 34796 46572 34848 46578
rect 34796 46514 34848 46520
rect 34808 45830 34836 46514
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 35636 46170 35664 46990
rect 36004 46714 36032 49200
rect 36832 46918 36860 49200
rect 36820 46912 36872 46918
rect 36820 46854 36872 46860
rect 37200 46714 37228 49200
rect 38028 47258 38056 49200
rect 38016 47252 38068 47258
rect 38488 47240 38516 49200
rect 39316 47258 39344 49200
rect 38660 47252 38712 47258
rect 38488 47212 38660 47240
rect 38016 47194 38068 47200
rect 38660 47194 38712 47200
rect 39304 47252 39356 47258
rect 39304 47194 39356 47200
rect 37556 47048 37608 47054
rect 37556 46990 37608 46996
rect 38660 47048 38712 47054
rect 38660 46990 38712 46996
rect 38752 47048 38804 47054
rect 38752 46990 38804 46996
rect 37568 46714 37596 46990
rect 38672 46714 38700 46990
rect 35992 46708 36044 46714
rect 35992 46650 36044 46656
rect 37188 46708 37240 46714
rect 37188 46650 37240 46656
rect 37556 46708 37608 46714
rect 37556 46650 37608 46656
rect 38660 46708 38712 46714
rect 38660 46650 38712 46656
rect 36268 46572 36320 46578
rect 36268 46514 36320 46520
rect 37372 46572 37424 46578
rect 37372 46514 37424 46520
rect 35440 46164 35492 46170
rect 35440 46106 35492 46112
rect 35624 46164 35676 46170
rect 35624 46106 35676 46112
rect 35452 45830 35480 46106
rect 35992 45960 36044 45966
rect 35992 45902 36044 45908
rect 34796 45824 34848 45830
rect 34796 45766 34848 45772
rect 35440 45824 35492 45830
rect 35440 45766 35492 45772
rect 34612 45280 34664 45286
rect 34612 45222 34664 45228
rect 33232 45076 33284 45082
rect 33232 45018 33284 45024
rect 33508 45076 33560 45082
rect 33508 45018 33560 45024
rect 34336 45076 34388 45082
rect 34336 45018 34388 45024
rect 32220 44940 32272 44946
rect 32220 44882 32272 44888
rect 33140 44940 33192 44946
rect 33140 44882 33192 44888
rect 32232 44742 32260 44882
rect 33232 44872 33284 44878
rect 33232 44814 33284 44820
rect 32220 44736 32272 44742
rect 32220 44678 32272 44684
rect 31760 44464 31812 44470
rect 31390 44432 31446 44441
rect 31760 44406 31812 44412
rect 31390 44367 31392 44376
rect 31444 44367 31446 44376
rect 31392 44338 31444 44344
rect 31116 44328 31168 44334
rect 31300 44328 31352 44334
rect 31116 44270 31168 44276
rect 31206 44296 31262 44305
rect 31128 43654 31156 44270
rect 31300 44270 31352 44276
rect 31206 44231 31208 44240
rect 31260 44231 31262 44240
rect 31208 44202 31260 44208
rect 31576 43784 31628 43790
rect 31576 43726 31628 43732
rect 31116 43648 31168 43654
rect 31116 43590 31168 43596
rect 31588 43314 31616 43726
rect 31852 43648 31904 43654
rect 31852 43590 31904 43596
rect 31576 43308 31628 43314
rect 31576 43250 31628 43256
rect 31300 43104 31352 43110
rect 31300 43046 31352 43052
rect 31116 42696 31168 42702
rect 31116 42638 31168 42644
rect 31128 41750 31156 42638
rect 31116 41744 31168 41750
rect 31116 41686 31168 41692
rect 31312 41614 31340 43046
rect 31588 42022 31616 43250
rect 31576 42016 31628 42022
rect 31628 41964 31708 41970
rect 31576 41958 31708 41964
rect 31588 41942 31708 41958
rect 31680 41614 31708 41942
rect 31864 41682 31892 43590
rect 31944 43240 31996 43246
rect 31944 43182 31996 43188
rect 31956 42566 31984 43182
rect 31944 42560 31996 42566
rect 31944 42502 31996 42508
rect 31852 41676 31904 41682
rect 31852 41618 31904 41624
rect 31300 41608 31352 41614
rect 31300 41550 31352 41556
rect 31668 41608 31720 41614
rect 31668 41550 31720 41556
rect 31956 41546 31984 42502
rect 31944 41540 31996 41546
rect 31944 41482 31996 41488
rect 30852 41386 31248 41414
rect 30748 41268 30800 41274
rect 30748 41210 30800 41216
rect 31220 26234 31248 41386
rect 30944 26206 31248 26234
rect 30380 7948 30432 7954
rect 30380 7890 30432 7896
rect 30012 5024 30064 5030
rect 30012 4966 30064 4972
rect 30024 4622 30052 4966
rect 29920 4616 29972 4622
rect 29920 4558 29972 4564
rect 30012 4616 30064 4622
rect 30012 4558 30064 4564
rect 29828 3120 29880 3126
rect 29826 3088 29828 3097
rect 29880 3088 29882 3097
rect 29826 3023 29882 3032
rect 29828 2440 29880 2446
rect 29828 2382 29880 2388
rect 29840 800 29868 2382
rect 29932 800 29960 4558
rect 30024 800 30052 4558
rect 30564 4480 30616 4486
rect 30564 4422 30616 4428
rect 30748 4480 30800 4486
rect 30748 4422 30800 4428
rect 30104 3936 30156 3942
rect 30104 3878 30156 3884
rect 30196 3936 30248 3942
rect 30196 3878 30248 3884
rect 30116 800 30144 3878
rect 30208 3194 30236 3878
rect 30288 3664 30340 3670
rect 30288 3606 30340 3612
rect 30196 3188 30248 3194
rect 30196 3130 30248 3136
rect 30300 800 30328 3606
rect 30472 3528 30524 3534
rect 30378 3496 30434 3505
rect 30472 3470 30524 3476
rect 30378 3431 30434 3440
rect 30392 3058 30420 3431
rect 30380 3052 30432 3058
rect 30380 2994 30432 3000
rect 30484 800 30512 3470
rect 30576 3194 30604 4422
rect 30760 4146 30788 4422
rect 30748 4140 30800 4146
rect 30748 4082 30800 4088
rect 30760 4010 30788 4082
rect 30748 4004 30800 4010
rect 30748 3946 30800 3952
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 30564 3188 30616 3194
rect 30564 3130 30616 3136
rect 30668 2990 30696 3878
rect 30656 2984 30708 2990
rect 30656 2926 30708 2932
rect 30944 2514 30972 26206
rect 32232 6089 32260 44678
rect 33244 43874 33272 44814
rect 34348 44470 34376 45018
rect 34624 44878 34652 45222
rect 34808 45014 34836 45766
rect 36004 45558 36032 45902
rect 35992 45552 36044 45558
rect 36176 45552 36228 45558
rect 35992 45494 36044 45500
rect 36096 45500 36176 45506
rect 36096 45494 36228 45500
rect 35716 45484 35768 45490
rect 35716 45426 35768 45432
rect 35348 45416 35400 45422
rect 35348 45358 35400 45364
rect 35360 45286 35388 45358
rect 35348 45280 35400 45286
rect 35348 45222 35400 45228
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 35360 45082 35388 45222
rect 35348 45076 35400 45082
rect 35348 45018 35400 45024
rect 34796 45008 34848 45014
rect 34796 44950 34848 44956
rect 34612 44872 34664 44878
rect 34612 44814 34664 44820
rect 34704 44736 34756 44742
rect 34704 44678 34756 44684
rect 34336 44464 34388 44470
rect 34336 44406 34388 44412
rect 33244 43858 33364 43874
rect 32404 43852 32456 43858
rect 32404 43794 32456 43800
rect 33244 43852 33376 43858
rect 33244 43846 33324 43852
rect 32416 43314 32444 43794
rect 32864 43784 32916 43790
rect 32864 43726 32916 43732
rect 33140 43784 33192 43790
rect 33140 43726 33192 43732
rect 32496 43648 32548 43654
rect 32496 43590 32548 43596
rect 32404 43308 32456 43314
rect 32404 43250 32456 43256
rect 32508 42634 32536 43590
rect 32876 43382 32904 43726
rect 33152 43450 33180 43726
rect 33244 43450 33272 43846
rect 33324 43794 33376 43800
rect 34060 43716 34112 43722
rect 34060 43658 34112 43664
rect 33140 43444 33192 43450
rect 33140 43386 33192 43392
rect 33232 43444 33284 43450
rect 33232 43386 33284 43392
rect 32864 43376 32916 43382
rect 32864 43318 32916 43324
rect 33152 43314 33180 43386
rect 33140 43308 33192 43314
rect 33140 43250 33192 43256
rect 34072 42906 34100 43658
rect 34060 42900 34112 42906
rect 34060 42842 34112 42848
rect 32680 42696 32732 42702
rect 32680 42638 32732 42644
rect 32496 42628 32548 42634
rect 32496 42570 32548 42576
rect 32692 42294 32720 42638
rect 32680 42288 32732 42294
rect 32680 42230 32732 42236
rect 34716 42022 34744 44678
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 35072 43920 35124 43926
rect 35072 43862 35124 43868
rect 34796 43648 34848 43654
rect 34796 43590 34848 43596
rect 34808 42634 34836 43590
rect 35084 43450 35112 43862
rect 35256 43784 35308 43790
rect 35256 43726 35308 43732
rect 35072 43444 35124 43450
rect 35072 43386 35124 43392
rect 35268 43246 35296 43726
rect 35256 43240 35308 43246
rect 35256 43182 35308 43188
rect 35360 43178 35388 45018
rect 35728 44878 35756 45426
rect 36004 45354 36032 45494
rect 36096 45478 36216 45494
rect 35992 45348 36044 45354
rect 35992 45290 36044 45296
rect 35900 45008 35952 45014
rect 35900 44950 35952 44956
rect 35716 44872 35768 44878
rect 35716 44814 35768 44820
rect 35808 44872 35860 44878
rect 35808 44814 35860 44820
rect 35624 44192 35676 44198
rect 35624 44134 35676 44140
rect 35636 43790 35664 44134
rect 35728 43790 35756 44814
rect 35820 44742 35848 44814
rect 35808 44736 35860 44742
rect 35808 44678 35860 44684
rect 35912 43858 35940 44950
rect 36004 43858 36032 45290
rect 36096 44878 36124 45478
rect 36176 45416 36228 45422
rect 36176 45358 36228 45364
rect 36188 44946 36216 45358
rect 36176 44940 36228 44946
rect 36176 44882 36228 44888
rect 36084 44872 36136 44878
rect 36084 44814 36136 44820
rect 35900 43852 35952 43858
rect 35900 43794 35952 43800
rect 35992 43852 36044 43858
rect 35992 43794 36044 43800
rect 35624 43784 35676 43790
rect 35624 43726 35676 43732
rect 35716 43784 35768 43790
rect 35716 43726 35768 43732
rect 35348 43172 35400 43178
rect 35348 43114 35400 43120
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34796 42628 34848 42634
rect 34796 42570 34848 42576
rect 34704 42016 34756 42022
rect 34704 41958 34756 41964
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 35636 35894 35664 43726
rect 35728 43314 35756 43726
rect 35912 43314 35940 43794
rect 35716 43308 35768 43314
rect 35716 43250 35768 43256
rect 35900 43308 35952 43314
rect 35900 43250 35952 43256
rect 36096 43246 36124 44814
rect 36280 43722 36308 46514
rect 36452 45892 36504 45898
rect 36452 45834 36504 45840
rect 36464 45082 36492 45834
rect 37384 45830 37412 46514
rect 37372 45824 37424 45830
rect 37372 45766 37424 45772
rect 36452 45076 36504 45082
rect 36452 45018 36504 45024
rect 37384 44878 37412 45766
rect 38660 45484 38712 45490
rect 38764 45472 38792 46990
rect 39684 46714 39712 49200
rect 40512 47258 40540 49200
rect 40500 47252 40552 47258
rect 40500 47194 40552 47200
rect 40224 47116 40276 47122
rect 40224 47058 40276 47064
rect 39856 47048 39908 47054
rect 39856 46990 39908 46996
rect 39672 46708 39724 46714
rect 39672 46650 39724 46656
rect 39120 46572 39172 46578
rect 39120 46514 39172 46520
rect 39764 46572 39816 46578
rect 39764 46514 39816 46520
rect 39132 46170 39160 46514
rect 39120 46164 39172 46170
rect 39120 46106 39172 46112
rect 39132 45966 39160 46106
rect 39120 45960 39172 45966
rect 39120 45902 39172 45908
rect 39672 45960 39724 45966
rect 39672 45902 39724 45908
rect 39132 45558 39160 45902
rect 39120 45552 39172 45558
rect 39120 45494 39172 45500
rect 38712 45444 38792 45472
rect 38660 45426 38712 45432
rect 38672 45286 38700 45426
rect 38660 45280 38712 45286
rect 38660 45222 38712 45228
rect 39132 45082 39160 45494
rect 39684 45286 39712 45902
rect 39672 45280 39724 45286
rect 39672 45222 39724 45228
rect 39120 45076 39172 45082
rect 39120 45018 39172 45024
rect 39684 45014 39712 45222
rect 39672 45008 39724 45014
rect 39672 44950 39724 44956
rect 37372 44872 37424 44878
rect 37372 44814 37424 44820
rect 39776 43926 39804 46514
rect 39868 46170 39896 46990
rect 40132 46504 40184 46510
rect 39946 46472 40002 46481
rect 40132 46446 40184 46452
rect 39946 46407 40002 46416
rect 39856 46164 39908 46170
rect 39856 46106 39908 46112
rect 39960 46102 39988 46407
rect 40040 46368 40092 46374
rect 40040 46310 40092 46316
rect 39948 46096 40000 46102
rect 39948 46038 40000 46044
rect 40052 45422 40080 46310
rect 40144 46102 40172 46446
rect 40132 46096 40184 46102
rect 40132 46038 40184 46044
rect 40236 45626 40264 47058
rect 40972 46918 41000 49200
rect 41800 47258 41828 49200
rect 41788 47252 41840 47258
rect 41788 47194 41840 47200
rect 41052 47184 41104 47190
rect 41052 47126 41104 47132
rect 40960 46912 41012 46918
rect 40960 46854 41012 46860
rect 41064 46646 41092 47126
rect 41144 47048 41196 47054
rect 41144 46990 41196 46996
rect 41328 47048 41380 47054
rect 41328 46990 41380 46996
rect 41880 47048 41932 47054
rect 41880 46990 41932 46996
rect 41156 46646 41184 46990
rect 41052 46640 41104 46646
rect 40498 46608 40554 46617
rect 41052 46582 41104 46588
rect 41144 46640 41196 46646
rect 41144 46582 41196 46588
rect 40498 46543 40500 46552
rect 40552 46543 40554 46552
rect 41236 46572 41288 46578
rect 40500 46514 40552 46520
rect 41236 46514 41288 46520
rect 40224 45620 40276 45626
rect 40224 45562 40276 45568
rect 40040 45416 40092 45422
rect 40040 45358 40092 45364
rect 40512 44742 40540 46514
rect 41052 46436 41104 46442
rect 41052 46378 41104 46384
rect 41064 46345 41092 46378
rect 41050 46336 41106 46345
rect 41050 46271 41106 46280
rect 41248 45626 41276 46514
rect 41340 46170 41368 46990
rect 41786 46608 41842 46617
rect 41786 46543 41788 46552
rect 41840 46543 41842 46552
rect 41788 46514 41840 46520
rect 41892 46170 41920 46990
rect 42260 46714 42288 49200
rect 43088 47258 43116 49200
rect 43076 47252 43128 47258
rect 43076 47194 43128 47200
rect 43168 47048 43220 47054
rect 43168 46990 43220 46996
rect 42708 46980 42760 46986
rect 42708 46922 42760 46928
rect 42248 46708 42300 46714
rect 42248 46650 42300 46656
rect 42432 46572 42484 46578
rect 42432 46514 42484 46520
rect 41328 46164 41380 46170
rect 41328 46106 41380 46112
rect 41880 46164 41932 46170
rect 41880 46106 41932 46112
rect 41512 45960 41564 45966
rect 41512 45902 41564 45908
rect 41696 45960 41748 45966
rect 41696 45902 41748 45908
rect 41236 45620 41288 45626
rect 41236 45562 41288 45568
rect 41524 45490 41552 45902
rect 41708 45626 41736 45902
rect 42444 45626 42472 46514
rect 42720 46374 42748 46922
rect 42708 46368 42760 46374
rect 42708 46310 42760 46316
rect 43180 46170 43208 46990
rect 43456 46714 43484 49200
rect 44284 47258 44312 49200
rect 44272 47252 44324 47258
rect 44272 47194 44324 47200
rect 44180 47048 44232 47054
rect 44180 46990 44232 46996
rect 43444 46708 43496 46714
rect 43444 46650 43496 46656
rect 43536 46572 43588 46578
rect 43536 46514 43588 46520
rect 43168 46164 43220 46170
rect 43168 46106 43220 46112
rect 43548 45626 43576 46514
rect 44192 46170 44220 46990
rect 44744 46714 44772 49200
rect 44732 46708 44784 46714
rect 44732 46650 44784 46656
rect 44548 46572 44600 46578
rect 44548 46514 44600 46520
rect 45284 46572 45336 46578
rect 45284 46514 45336 46520
rect 44180 46164 44232 46170
rect 44180 46106 44232 46112
rect 43904 45960 43956 45966
rect 43904 45902 43956 45908
rect 43916 45626 43944 45902
rect 44560 45626 44588 46514
rect 45100 46368 45152 46374
rect 45100 46310 45152 46316
rect 45112 46102 45140 46310
rect 45100 46096 45152 46102
rect 45100 46038 45152 46044
rect 45296 45898 45324 46514
rect 45572 46170 45600 49200
rect 45650 49056 45706 49065
rect 45650 48991 45706 49000
rect 45664 47258 45692 48991
rect 45652 47252 45704 47258
rect 45652 47194 45704 47200
rect 45744 46980 45796 46986
rect 45744 46922 45796 46928
rect 45560 46164 45612 46170
rect 45560 46106 45612 46112
rect 44732 45892 44784 45898
rect 44732 45834 44784 45840
rect 45284 45892 45336 45898
rect 45284 45834 45336 45840
rect 41696 45620 41748 45626
rect 41696 45562 41748 45568
rect 42432 45620 42484 45626
rect 42432 45562 42484 45568
rect 43536 45620 43588 45626
rect 43536 45562 43588 45568
rect 43904 45620 43956 45626
rect 43904 45562 43956 45568
rect 44548 45620 44600 45626
rect 44548 45562 44600 45568
rect 41512 45484 41564 45490
rect 41512 45426 41564 45432
rect 40500 44736 40552 44742
rect 40500 44678 40552 44684
rect 38660 43920 38712 43926
rect 38660 43862 38712 43868
rect 39764 43920 39816 43926
rect 39764 43862 39816 43868
rect 36268 43716 36320 43722
rect 36268 43658 36320 43664
rect 36360 43716 36412 43722
rect 36360 43658 36412 43664
rect 36084 43240 36136 43246
rect 36084 43182 36136 43188
rect 36280 42838 36308 43658
rect 36372 43450 36400 43658
rect 36360 43444 36412 43450
rect 36360 43386 36412 43392
rect 38672 43314 38700 43862
rect 38660 43308 38712 43314
rect 38660 43250 38712 43256
rect 41524 42906 41552 45426
rect 43916 45082 43944 45562
rect 44456 45484 44508 45490
rect 44456 45426 44508 45432
rect 43904 45076 43956 45082
rect 43904 45018 43956 45024
rect 44468 44946 44496 45426
rect 44456 44940 44508 44946
rect 44456 44882 44508 44888
rect 44364 44736 44416 44742
rect 44364 44678 44416 44684
rect 44376 44266 44404 44678
rect 44744 44470 44772 45834
rect 45098 45520 45154 45529
rect 45098 45455 45100 45464
rect 45152 45455 45154 45464
rect 45100 45426 45152 45432
rect 45112 45082 45140 45426
rect 45652 45416 45704 45422
rect 45652 45358 45704 45364
rect 45100 45076 45152 45082
rect 45100 45018 45152 45024
rect 45664 44538 45692 45358
rect 45756 44878 45784 46922
rect 45940 45354 45968 49200
rect 46202 48376 46258 48385
rect 46202 48311 46258 48320
rect 46216 46714 46244 48311
rect 46204 46708 46256 46714
rect 46204 46650 46256 46656
rect 46020 46572 46072 46578
rect 46020 46514 46072 46520
rect 46032 46345 46060 46514
rect 46204 46368 46256 46374
rect 46018 46336 46074 46345
rect 46204 46310 46256 46316
rect 46018 46271 46074 46280
rect 46020 45484 46072 45490
rect 46020 45426 46072 45432
rect 45836 45348 45888 45354
rect 45836 45290 45888 45296
rect 45928 45348 45980 45354
rect 45928 45290 45980 45296
rect 45744 44872 45796 44878
rect 45744 44814 45796 44820
rect 45652 44532 45704 44538
rect 45652 44474 45704 44480
rect 44732 44464 44784 44470
rect 44732 44406 44784 44412
rect 44364 44260 44416 44266
rect 44364 44202 44416 44208
rect 45664 43926 45692 44474
rect 45756 44402 45784 44814
rect 45848 44538 45876 45290
rect 46032 45082 46060 45426
rect 46020 45076 46072 45082
rect 46020 45018 46072 45024
rect 45836 44532 45888 44538
rect 45836 44474 45888 44480
rect 45744 44396 45796 44402
rect 45744 44338 45796 44344
rect 46216 43926 46244 46310
rect 46492 46170 46520 49671
rect 46754 49200 46810 50000
rect 47214 49200 47270 50000
rect 47582 49200 47638 50000
rect 48042 49200 48098 50000
rect 48410 49200 48466 50000
rect 48870 49200 48926 50000
rect 49238 49200 49294 50000
rect 49698 49200 49754 50000
rect 46662 46472 46718 46481
rect 46662 46407 46718 46416
rect 46480 46164 46532 46170
rect 46480 46106 46532 46112
rect 46480 45960 46532 45966
rect 46480 45902 46532 45908
rect 46492 45286 46520 45902
rect 46480 45280 46532 45286
rect 46480 45222 46532 45228
rect 46676 43926 46704 46407
rect 46768 46102 46796 49200
rect 46848 47184 46900 47190
rect 46846 47152 46848 47161
rect 46900 47152 46902 47161
rect 46846 47087 46902 47096
rect 46756 46096 46808 46102
rect 46756 46038 46808 46044
rect 46848 45280 46900 45286
rect 46848 45222 46900 45228
rect 46860 45121 46888 45222
rect 46846 45112 46902 45121
rect 46846 45047 46902 45056
rect 46848 44736 46900 44742
rect 46848 44678 46900 44684
rect 46860 44441 46888 44678
rect 46846 44432 46902 44441
rect 46846 44367 46902 44376
rect 46940 44396 46992 44402
rect 46940 44338 46992 44344
rect 46952 44198 46980 44338
rect 46940 44192 46992 44198
rect 46940 44134 46992 44140
rect 46952 43994 46980 44134
rect 47228 43994 47256 49200
rect 47306 47696 47362 47705
rect 47306 47631 47362 47640
rect 47320 46170 47348 47631
rect 47308 46164 47360 46170
rect 47308 46106 47360 46112
rect 47596 45082 47624 49200
rect 47952 47048 48004 47054
rect 47952 46990 48004 46996
rect 47860 46572 47912 46578
rect 47860 46514 47912 46520
rect 47872 46481 47900 46514
rect 47858 46472 47914 46481
rect 47858 46407 47914 46416
rect 47860 45960 47912 45966
rect 47860 45902 47912 45908
rect 47584 45076 47636 45082
rect 47584 45018 47636 45024
rect 47308 44940 47360 44946
rect 47308 44882 47360 44888
rect 46940 43988 46992 43994
rect 46940 43930 46992 43936
rect 47216 43988 47268 43994
rect 47216 43930 47268 43936
rect 45652 43920 45704 43926
rect 45652 43862 45704 43868
rect 46204 43920 46256 43926
rect 46204 43862 46256 43868
rect 46664 43920 46716 43926
rect 46664 43862 46716 43868
rect 47320 43790 47348 44882
rect 47676 44872 47728 44878
rect 47676 44814 47728 44820
rect 47688 44470 47716 44814
rect 47872 44538 47900 45902
rect 47860 44532 47912 44538
rect 47860 44474 47912 44480
rect 47676 44464 47728 44470
rect 47676 44406 47728 44412
rect 47964 43994 47992 46990
rect 48056 46646 48084 49200
rect 48424 47258 48452 49200
rect 48412 47252 48464 47258
rect 48412 47194 48464 47200
rect 48884 46714 48912 49200
rect 49252 47190 49280 49200
rect 49240 47184 49292 47190
rect 49240 47126 49292 47132
rect 48872 46708 48924 46714
rect 48872 46650 48924 46656
rect 48044 46640 48096 46646
rect 48044 46582 48096 46588
rect 48042 46472 48098 46481
rect 48042 46407 48044 46416
rect 48096 46407 48098 46416
rect 48044 46378 48096 46384
rect 48044 45824 48096 45830
rect 48042 45792 48044 45801
rect 48096 45792 48098 45801
rect 48042 45727 48098 45736
rect 49712 45626 49740 49200
rect 49700 45620 49752 45626
rect 49700 45562 49752 45568
rect 48044 44192 48096 44198
rect 48044 44134 48096 44140
rect 47952 43988 48004 43994
rect 47952 43930 48004 43936
rect 48056 43897 48084 44134
rect 48042 43888 48098 43897
rect 48042 43823 48098 43832
rect 47308 43784 47360 43790
rect 47308 43726 47360 43732
rect 46940 43308 46992 43314
rect 46940 43250 46992 43256
rect 46952 43110 46980 43250
rect 48042 43208 48098 43217
rect 48042 43143 48044 43152
rect 48096 43143 48098 43152
rect 48044 43114 48096 43120
rect 46940 43104 46992 43110
rect 46940 43046 46992 43052
rect 41512 42900 41564 42906
rect 41512 42842 41564 42848
rect 36268 42832 36320 42838
rect 36268 42774 36320 42780
rect 46296 41540 46348 41546
rect 46296 41482 46348 41488
rect 45560 39296 45612 39302
rect 45560 39238 45612 39244
rect 35636 35866 35756 35894
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 33140 15564 33192 15570
rect 33140 15506 33192 15512
rect 33152 8974 33180 15506
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 33140 8968 33192 8974
rect 33140 8910 33192 8916
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 32218 6080 32274 6089
rect 32218 6015 32274 6024
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 31392 4480 31444 4486
rect 31392 4422 31444 4428
rect 31404 4146 31432 4422
rect 31392 4140 31444 4146
rect 31392 4082 31444 4088
rect 31208 3936 31260 3942
rect 31208 3878 31260 3884
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 30932 2508 30984 2514
rect 30932 2450 30984 2456
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 30760 800 30788 2382
rect 31036 800 31064 3470
rect 31116 3392 31168 3398
rect 31116 3334 31168 3340
rect 31128 3194 31156 3334
rect 31116 3188 31168 3194
rect 31116 3130 31168 3136
rect 31220 2990 31248 3878
rect 31404 3670 31432 4082
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 31392 3664 31444 3670
rect 31392 3606 31444 3612
rect 31944 3528 31996 3534
rect 31944 3470 31996 3476
rect 33140 3528 33192 3534
rect 33140 3470 33192 3476
rect 34612 3528 34664 3534
rect 34612 3470 34664 3476
rect 35348 3528 35400 3534
rect 35348 3470 35400 3476
rect 31208 2984 31260 2990
rect 31208 2926 31260 2932
rect 31392 2848 31444 2854
rect 31392 2790 31444 2796
rect 31404 800 31432 2790
rect 31668 2440 31720 2446
rect 31668 2382 31720 2388
rect 31680 800 31708 2382
rect 31956 800 31984 3470
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 32864 2848 32916 2854
rect 32864 2790 32916 2796
rect 32232 800 32260 2790
rect 32588 2440 32640 2446
rect 32588 2382 32640 2388
rect 32600 800 32628 2382
rect 32876 800 32904 2790
rect 33152 800 33180 3470
rect 33416 2984 33468 2990
rect 33416 2926 33468 2932
rect 33428 800 33456 2926
rect 34060 2848 34112 2854
rect 34060 2790 34112 2796
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 33796 800 33824 2382
rect 34072 800 34100 2790
rect 34336 2440 34388 2446
rect 34336 2382 34388 2388
rect 34348 800 34376 2382
rect 34624 800 34652 3470
rect 35256 3460 35308 3466
rect 35256 3402 35308 3408
rect 35268 3126 35296 3402
rect 35256 3120 35308 3126
rect 35256 3062 35308 3068
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 34980 2440 35032 2446
rect 34980 2382 35032 2388
rect 34992 800 35020 2382
rect 35360 1850 35388 3470
rect 35728 3126 35756 35866
rect 44640 28416 44692 28422
rect 44640 28358 44692 28364
rect 44272 22976 44324 22982
rect 44272 22918 44324 22924
rect 40684 19984 40736 19990
rect 40684 19926 40736 19932
rect 40696 19446 40724 19926
rect 40684 19440 40736 19446
rect 40684 19382 40736 19388
rect 39304 19372 39356 19378
rect 39304 19314 39356 19320
rect 37924 14952 37976 14958
rect 37924 14894 37976 14900
rect 36636 13864 36688 13870
rect 36636 13806 36688 13812
rect 36648 7886 36676 13806
rect 37648 8900 37700 8906
rect 37648 8842 37700 8848
rect 37660 8566 37688 8842
rect 37648 8560 37700 8566
rect 37648 8502 37700 8508
rect 36636 7880 36688 7886
rect 36636 7822 36688 7828
rect 37936 4622 37964 14894
rect 39316 7818 39344 19314
rect 44284 12434 44312 22918
rect 44284 12406 44404 12434
rect 39304 7812 39356 7818
rect 39304 7754 39356 7760
rect 43076 7744 43128 7750
rect 43076 7686 43128 7692
rect 44272 7744 44324 7750
rect 44272 7686 44324 7692
rect 43088 7410 43116 7686
rect 44284 7478 44312 7686
rect 44272 7472 44324 7478
rect 44272 7414 44324 7420
rect 43076 7404 43128 7410
rect 43076 7346 43128 7352
rect 43168 7404 43220 7410
rect 43168 7346 43220 7352
rect 44088 7404 44140 7410
rect 44088 7346 44140 7352
rect 43180 7206 43208 7346
rect 44100 7274 44128 7346
rect 44088 7268 44140 7274
rect 44088 7210 44140 7216
rect 42800 7200 42852 7206
rect 42800 7142 42852 7148
rect 43168 7200 43220 7206
rect 43168 7142 43220 7148
rect 42812 6798 42840 7142
rect 42800 6792 42852 6798
rect 42800 6734 42852 6740
rect 43180 6254 43208 7142
rect 44180 6860 44232 6866
rect 44180 6802 44232 6808
rect 43258 6760 43314 6769
rect 43258 6695 43260 6704
rect 43312 6695 43314 6704
rect 43260 6666 43312 6672
rect 44086 6488 44142 6497
rect 44086 6423 44088 6432
rect 44140 6423 44142 6432
rect 44088 6394 44140 6400
rect 39304 6248 39356 6254
rect 39304 6190 39356 6196
rect 43168 6248 43220 6254
rect 43168 6190 43220 6196
rect 37924 4616 37976 4622
rect 37924 4558 37976 4564
rect 39316 3670 39344 6190
rect 43260 6180 43312 6186
rect 43260 6122 43312 6128
rect 42064 5568 42116 5574
rect 42064 5510 42116 5516
rect 42616 5568 42668 5574
rect 42616 5510 42668 5516
rect 41328 5024 41380 5030
rect 41328 4966 41380 4972
rect 40408 4480 40460 4486
rect 40408 4422 40460 4428
rect 40868 4480 40920 4486
rect 40868 4422 40920 4428
rect 40420 4049 40448 4422
rect 40406 4040 40462 4049
rect 40406 3975 40462 3984
rect 39304 3664 39356 3670
rect 39304 3606 39356 3612
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 36176 3528 36228 3534
rect 36176 3470 36228 3476
rect 37004 3528 37056 3534
rect 37004 3470 37056 3476
rect 38200 3528 38252 3534
rect 38200 3470 38252 3476
rect 39120 3528 39172 3534
rect 39120 3470 39172 3476
rect 40316 3528 40368 3534
rect 40316 3470 40368 3476
rect 35716 3120 35768 3126
rect 35716 3062 35768 3068
rect 35532 2440 35584 2446
rect 35532 2382 35584 2388
rect 35268 1822 35388 1850
rect 35268 800 35296 1822
rect 35544 800 35572 2382
rect 35820 800 35848 3470
rect 35900 3460 35952 3466
rect 35900 3402 35952 3408
rect 35912 3194 35940 3402
rect 36084 3392 36136 3398
rect 36084 3334 36136 3340
rect 36096 3194 36124 3334
rect 35900 3188 35952 3194
rect 35900 3130 35952 3136
rect 36084 3188 36136 3194
rect 36084 3130 36136 3136
rect 36188 800 36216 3470
rect 36452 2848 36504 2854
rect 36452 2790 36504 2796
rect 36464 800 36492 2790
rect 36728 2440 36780 2446
rect 36728 2382 36780 2388
rect 36740 800 36768 2382
rect 37016 800 37044 3470
rect 37924 2984 37976 2990
rect 37924 2926 37976 2932
rect 37372 2848 37424 2854
rect 37372 2790 37424 2796
rect 37384 800 37412 2790
rect 37648 2440 37700 2446
rect 37648 2382 37700 2388
rect 37660 800 37688 2382
rect 37936 800 37964 2926
rect 38212 800 38240 3470
rect 38568 2848 38620 2854
rect 38568 2790 38620 2796
rect 38580 800 38608 2790
rect 38844 2440 38896 2446
rect 38844 2382 38896 2388
rect 38856 800 38884 2382
rect 39132 800 39160 3470
rect 39396 2848 39448 2854
rect 39396 2790 39448 2796
rect 40040 2848 40092 2854
rect 40040 2790 40092 2796
rect 39408 800 39436 2790
rect 39764 2440 39816 2446
rect 39764 2382 39816 2388
rect 39776 800 39804 2382
rect 40052 800 40080 2790
rect 40328 800 40356 3470
rect 40420 3466 40448 3975
rect 40684 3936 40736 3942
rect 40684 3878 40736 3884
rect 40696 3738 40724 3878
rect 40684 3732 40736 3738
rect 40684 3674 40736 3680
rect 40408 3460 40460 3466
rect 40408 3402 40460 3408
rect 40696 3058 40724 3674
rect 40684 3052 40736 3058
rect 40684 2994 40736 3000
rect 40880 2922 40908 4422
rect 41340 4214 41368 4966
rect 42076 4622 42104 5510
rect 42628 5302 42656 5510
rect 42616 5296 42668 5302
rect 42616 5238 42668 5244
rect 42064 4616 42116 4622
rect 42064 4558 42116 4564
rect 42524 4616 42576 4622
rect 42524 4558 42576 4564
rect 41512 4480 41564 4486
rect 41512 4422 41564 4428
rect 41524 4282 41552 4422
rect 41512 4276 41564 4282
rect 41512 4218 41564 4224
rect 41328 4208 41380 4214
rect 41328 4150 41380 4156
rect 41236 3528 41288 3534
rect 41236 3470 41288 3476
rect 40868 2916 40920 2922
rect 40868 2858 40920 2864
rect 40684 2848 40736 2854
rect 40684 2790 40736 2796
rect 40696 800 40724 2790
rect 40960 2440 41012 2446
rect 40960 2382 41012 2388
rect 40972 800 41000 2382
rect 41248 800 41276 3470
rect 41340 2514 41368 4150
rect 41696 4140 41748 4146
rect 41696 4082 41748 4088
rect 41708 3126 41736 4082
rect 41880 3936 41932 3942
rect 41880 3878 41932 3884
rect 41892 3641 41920 3878
rect 41878 3632 41934 3641
rect 41878 3567 41934 3576
rect 42156 3528 42208 3534
rect 42156 3470 42208 3476
rect 41696 3120 41748 3126
rect 41696 3062 41748 3068
rect 41880 2848 41932 2854
rect 41880 2790 41932 2796
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 41512 2440 41564 2446
rect 41512 2382 41564 2388
rect 41524 800 41552 2382
rect 41892 800 41920 2790
rect 42168 800 42196 3470
rect 42536 2650 42564 4558
rect 42524 2644 42576 2650
rect 42524 2586 42576 2592
rect 42432 2440 42484 2446
rect 42432 2382 42484 2388
rect 42444 800 42472 2382
rect 42628 921 42656 5238
rect 43272 5234 43300 6122
rect 43628 5704 43680 5710
rect 43628 5646 43680 5652
rect 44088 5704 44140 5710
rect 44088 5646 44140 5652
rect 43260 5228 43312 5234
rect 43260 5170 43312 5176
rect 42800 3936 42852 3942
rect 42800 3878 42852 3884
rect 42812 3369 42840 3878
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 42798 3360 42854 3369
rect 42798 3295 42854 3304
rect 42708 2848 42760 2854
rect 42708 2790 42760 2796
rect 42614 912 42670 921
rect 42614 847 42670 856
rect 42720 800 42748 2790
rect 43088 800 43116 3470
rect 43272 2582 43300 5170
rect 43640 4865 43668 5646
rect 44100 5302 44128 5646
rect 44192 5302 44220 6802
rect 44272 6452 44324 6458
rect 44272 6394 44324 6400
rect 44284 5574 44312 6394
rect 44272 5568 44324 5574
rect 44272 5510 44324 5516
rect 44088 5296 44140 5302
rect 44088 5238 44140 5244
rect 44180 5296 44232 5302
rect 44180 5238 44232 5244
rect 43626 4856 43682 4865
rect 43626 4791 43682 4800
rect 44376 4570 44404 12406
rect 44652 8634 44680 28358
rect 45376 24064 45428 24070
rect 45376 24006 45428 24012
rect 44824 19780 44876 19786
rect 44824 19722 44876 19728
rect 44836 12434 44864 19722
rect 45192 12912 45244 12918
rect 45192 12854 45244 12860
rect 44744 12406 44864 12434
rect 44640 8628 44692 8634
rect 44640 8570 44692 8576
rect 44652 7818 44680 8570
rect 44548 7812 44600 7818
rect 44548 7754 44600 7760
rect 44640 7812 44692 7818
rect 44640 7754 44692 7760
rect 44456 6928 44508 6934
rect 44456 6870 44508 6876
rect 44468 6390 44496 6870
rect 44456 6384 44508 6390
rect 44456 6326 44508 6332
rect 44560 6322 44588 7754
rect 44548 6316 44600 6322
rect 44548 6258 44600 6264
rect 44744 6202 44772 12406
rect 45204 11014 45232 12854
rect 45284 12436 45336 12442
rect 45284 12378 45336 12384
rect 45296 11762 45324 12378
rect 45284 11756 45336 11762
rect 45284 11698 45336 11704
rect 45192 11008 45244 11014
rect 45192 10950 45244 10956
rect 45388 9674 45416 24006
rect 45468 21888 45520 21894
rect 45468 21830 45520 21836
rect 45296 9646 45416 9674
rect 45192 8968 45244 8974
rect 45192 8910 45244 8916
rect 45100 7404 45152 7410
rect 45100 7346 45152 7352
rect 45112 7274 45140 7346
rect 45204 7274 45232 8910
rect 45100 7268 45152 7274
rect 45100 7210 45152 7216
rect 45192 7268 45244 7274
rect 45192 7210 45244 7216
rect 44824 6792 44876 6798
rect 44822 6760 44824 6769
rect 44876 6760 44878 6769
rect 44822 6695 44878 6704
rect 44468 6174 44772 6202
rect 44468 5778 44496 6174
rect 44548 6112 44600 6118
rect 44548 6054 44600 6060
rect 44560 5778 44588 6054
rect 44456 5772 44508 5778
rect 44456 5714 44508 5720
rect 44548 5772 44600 5778
rect 44548 5714 44600 5720
rect 44640 5364 44692 5370
rect 44640 5306 44692 5312
rect 44456 5228 44508 5234
rect 44456 5170 44508 5176
rect 44192 4554 44404 4570
rect 44180 4548 44404 4554
rect 44232 4542 44404 4548
rect 44180 4490 44232 4496
rect 44178 4040 44234 4049
rect 44178 3975 44234 3984
rect 44192 2990 44220 3975
rect 44180 2984 44232 2990
rect 44180 2926 44232 2932
rect 43352 2848 43404 2854
rect 43352 2790 43404 2796
rect 43904 2848 43956 2854
rect 43904 2790 43956 2796
rect 43260 2576 43312 2582
rect 43260 2518 43312 2524
rect 43364 800 43392 2790
rect 43628 2440 43680 2446
rect 43628 2382 43680 2388
rect 43640 800 43668 2382
rect 43916 800 43944 2790
rect 44272 2440 44324 2446
rect 44272 2382 44324 2388
rect 44284 800 44312 2382
rect 44468 1358 44496 5170
rect 44652 4554 44680 5306
rect 44640 4548 44692 4554
rect 44640 4490 44692 4496
rect 44836 3505 44864 6695
rect 45204 6322 45232 7210
rect 44916 6316 44968 6322
rect 44916 6258 44968 6264
rect 45192 6316 45244 6322
rect 45192 6258 45244 6264
rect 44928 4321 44956 6258
rect 45100 6112 45152 6118
rect 45100 6054 45152 6060
rect 45008 5840 45060 5846
rect 45008 5782 45060 5788
rect 45020 4622 45048 5782
rect 45112 5166 45140 6054
rect 45204 5846 45232 6258
rect 45192 5840 45244 5846
rect 45192 5782 45244 5788
rect 45192 5568 45244 5574
rect 45192 5510 45244 5516
rect 45100 5160 45152 5166
rect 45100 5102 45152 5108
rect 45112 4690 45140 5102
rect 45100 4684 45152 4690
rect 45100 4626 45152 4632
rect 45008 4616 45060 4622
rect 45008 4558 45060 4564
rect 44914 4312 44970 4321
rect 44914 4247 44970 4256
rect 45112 4078 45140 4626
rect 45204 4146 45232 5510
rect 45296 5284 45324 9646
rect 45480 7970 45508 21830
rect 45572 18290 45600 39238
rect 45836 36644 45888 36650
rect 45836 36586 45888 36592
rect 45652 31204 45704 31210
rect 45652 31146 45704 31152
rect 45560 18284 45612 18290
rect 45560 18226 45612 18232
rect 45560 17604 45612 17610
rect 45560 17546 45612 17552
rect 45572 15162 45600 17546
rect 45664 17218 45692 31146
rect 45744 29504 45796 29510
rect 45744 29446 45796 29452
rect 45756 17354 45784 29446
rect 45848 21350 45876 36586
rect 45928 35556 45980 35562
rect 45928 35498 45980 35504
rect 45836 21344 45888 21350
rect 45836 21286 45888 21292
rect 45940 21162 45968 35498
rect 46020 32292 46072 32298
rect 46020 32234 46072 32240
rect 45848 21134 45968 21162
rect 45848 17610 45876 21134
rect 45928 21072 45980 21078
rect 45928 21014 45980 21020
rect 45940 19854 45968 21014
rect 45928 19848 45980 19854
rect 45928 19790 45980 19796
rect 45928 18828 45980 18834
rect 45928 18770 45980 18776
rect 45940 18222 45968 18770
rect 45928 18216 45980 18222
rect 45928 18158 45980 18164
rect 45836 17604 45888 17610
rect 45836 17546 45888 17552
rect 45928 17536 45980 17542
rect 45928 17478 45980 17484
rect 45756 17326 45876 17354
rect 45940 17338 45968 17478
rect 45664 17190 45784 17218
rect 45652 17128 45704 17134
rect 45652 17070 45704 17076
rect 45560 15156 45612 15162
rect 45560 15098 45612 15104
rect 45560 15020 45612 15026
rect 45560 14962 45612 14968
rect 45572 14657 45600 14962
rect 45558 14648 45614 14657
rect 45558 14583 45614 14592
rect 45664 14498 45692 17070
rect 45572 14470 45692 14498
rect 45572 12102 45600 14470
rect 45652 12776 45704 12782
rect 45652 12718 45704 12724
rect 45560 12096 45612 12102
rect 45560 12038 45612 12044
rect 45560 11688 45612 11694
rect 45560 11630 45612 11636
rect 45572 9450 45600 11630
rect 45560 9444 45612 9450
rect 45560 9386 45612 9392
rect 45664 9110 45692 12718
rect 45756 11218 45784 17190
rect 45848 12918 45876 17326
rect 45928 17332 45980 17338
rect 45928 17274 45980 17280
rect 45928 17128 45980 17134
rect 45928 17070 45980 17076
rect 45940 16522 45968 17070
rect 45928 16516 45980 16522
rect 45928 16458 45980 16464
rect 45928 16108 45980 16114
rect 45928 16050 45980 16056
rect 45940 15881 45968 16050
rect 45926 15872 45982 15881
rect 45926 15807 45982 15816
rect 46032 15722 46060 32234
rect 46112 21344 46164 21350
rect 46112 21286 46164 21292
rect 46124 18290 46152 21286
rect 46308 20602 46336 41482
rect 46952 40730 46980 43046
rect 47308 42560 47360 42566
rect 48044 42560 48096 42566
rect 47308 42502 47360 42508
rect 48042 42528 48044 42537
rect 48096 42528 48098 42537
rect 47320 41818 47348 42502
rect 48042 42463 48098 42472
rect 48044 42016 48096 42022
rect 48044 41958 48096 41964
rect 48056 41857 48084 41958
rect 48042 41848 48098 41857
rect 47308 41812 47360 41818
rect 48042 41783 48098 41792
rect 47308 41754 47360 41760
rect 48044 41608 48096 41614
rect 48044 41550 48096 41556
rect 48056 41313 48084 41550
rect 48042 41304 48098 41313
rect 48042 41239 48098 41248
rect 48044 41132 48096 41138
rect 48044 41074 48096 41080
rect 47032 40996 47084 41002
rect 47032 40938 47084 40944
rect 46940 40724 46992 40730
rect 46940 40666 46992 40672
rect 46572 38208 46624 38214
rect 46572 38150 46624 38156
rect 46480 20868 46532 20874
rect 46480 20810 46532 20816
rect 46296 20596 46348 20602
rect 46296 20538 46348 20544
rect 46308 19854 46336 20538
rect 46296 19848 46348 19854
rect 46296 19790 46348 19796
rect 46388 19848 46440 19854
rect 46388 19790 46440 19796
rect 46204 19780 46256 19786
rect 46204 19722 46256 19728
rect 46216 19378 46244 19722
rect 46400 19446 46428 19790
rect 46388 19440 46440 19446
rect 46388 19382 46440 19388
rect 46204 19372 46256 19378
rect 46204 19314 46256 19320
rect 46112 18284 46164 18290
rect 46112 18226 46164 18232
rect 46112 18080 46164 18086
rect 46112 18022 46164 18028
rect 45940 15694 46060 15722
rect 45836 12912 45888 12918
rect 45836 12854 45888 12860
rect 45834 12744 45890 12753
rect 45834 12679 45890 12688
rect 45744 11212 45796 11218
rect 45744 11154 45796 11160
rect 45848 11150 45876 12679
rect 45940 11830 45968 15694
rect 46020 15632 46072 15638
rect 46020 15574 46072 15580
rect 46032 14414 46060 15574
rect 46020 14408 46072 14414
rect 46020 14350 46072 14356
rect 46032 12646 46060 14350
rect 46020 12640 46072 12646
rect 46020 12582 46072 12588
rect 46018 12472 46074 12481
rect 46018 12407 46074 12416
rect 46032 12306 46060 12407
rect 46020 12300 46072 12306
rect 46020 12242 46072 12248
rect 46124 12209 46152 18022
rect 46110 12200 46166 12209
rect 46110 12135 46166 12144
rect 46020 12096 46072 12102
rect 46020 12038 46072 12044
rect 46112 12096 46164 12102
rect 46112 12038 46164 12044
rect 45928 11824 45980 11830
rect 45928 11766 45980 11772
rect 45928 11280 45980 11286
rect 45928 11222 45980 11228
rect 45836 11144 45888 11150
rect 45836 11086 45888 11092
rect 45744 11008 45796 11014
rect 45744 10950 45796 10956
rect 45756 10266 45784 10950
rect 45940 10826 45968 11222
rect 45848 10798 45968 10826
rect 45744 10260 45796 10266
rect 45744 10202 45796 10208
rect 45848 9674 45876 10798
rect 45928 10668 45980 10674
rect 45928 10610 45980 10616
rect 45756 9646 45876 9674
rect 45652 9104 45704 9110
rect 45652 9046 45704 9052
rect 45756 8362 45784 9646
rect 45836 9512 45888 9518
rect 45836 9454 45888 9460
rect 45848 9178 45876 9454
rect 45836 9172 45888 9178
rect 45836 9114 45888 9120
rect 45560 8356 45612 8362
rect 45560 8298 45612 8304
rect 45744 8356 45796 8362
rect 45744 8298 45796 8304
rect 45572 8129 45600 8298
rect 45558 8120 45614 8129
rect 45756 8090 45784 8298
rect 45558 8055 45614 8064
rect 45744 8084 45796 8090
rect 45744 8026 45796 8032
rect 45388 7942 45508 7970
rect 45388 7018 45416 7942
rect 45652 7880 45704 7886
rect 45652 7822 45704 7828
rect 45468 7812 45520 7818
rect 45468 7754 45520 7760
rect 45480 7274 45508 7754
rect 45664 7478 45692 7822
rect 45652 7472 45704 7478
rect 45652 7414 45704 7420
rect 45940 7410 45968 10610
rect 45928 7404 45980 7410
rect 45928 7346 45980 7352
rect 45468 7268 45520 7274
rect 45468 7210 45520 7216
rect 46032 7206 46060 12038
rect 46124 11286 46152 12038
rect 46112 11280 46164 11286
rect 46112 11222 46164 11228
rect 46112 11144 46164 11150
rect 46112 11086 46164 11092
rect 46124 7886 46152 11086
rect 46216 8974 46244 19314
rect 46296 18760 46348 18766
rect 46296 18702 46348 18708
rect 46308 18465 46336 18702
rect 46294 18456 46350 18465
rect 46294 18391 46350 18400
rect 46296 18284 46348 18290
rect 46296 18226 46348 18232
rect 46308 16794 46336 18226
rect 46296 16788 46348 16794
rect 46296 16730 46348 16736
rect 46296 16584 46348 16590
rect 46294 16552 46296 16561
rect 46348 16552 46350 16561
rect 46294 16487 46350 16496
rect 46296 15904 46348 15910
rect 46296 15846 46348 15852
rect 46308 15502 46336 15846
rect 46296 15496 46348 15502
rect 46296 15438 46348 15444
rect 46308 13977 46336 15438
rect 46294 13968 46350 13977
rect 46294 13903 46350 13912
rect 46296 13320 46348 13326
rect 46296 13262 46348 13268
rect 46308 12617 46336 13262
rect 46400 12730 46428 19382
rect 46492 19378 46520 20810
rect 46480 19372 46532 19378
rect 46480 19314 46532 19320
rect 46480 18624 46532 18630
rect 46480 18566 46532 18572
rect 46492 18290 46520 18566
rect 46480 18284 46532 18290
rect 46480 18226 46532 18232
rect 46480 17604 46532 17610
rect 46480 17546 46532 17552
rect 46492 16794 46520 17546
rect 46584 17542 46612 38150
rect 47044 35894 47072 40938
rect 48056 40730 48084 41074
rect 48044 40724 48096 40730
rect 48044 40666 48096 40672
rect 48056 40633 48084 40666
rect 48042 40624 48098 40633
rect 48042 40559 48098 40568
rect 48044 40384 48096 40390
rect 48044 40326 48096 40332
rect 48056 40118 48084 40326
rect 48044 40112 48096 40118
rect 48044 40054 48096 40060
rect 48056 39953 48084 40054
rect 48042 39944 48098 39953
rect 48042 39879 48098 39888
rect 48136 39840 48188 39846
rect 48136 39782 48188 39788
rect 48044 39364 48096 39370
rect 48044 39306 48096 39312
rect 48056 39273 48084 39306
rect 48042 39264 48098 39273
rect 48042 39199 48098 39208
rect 48044 38956 48096 38962
rect 48044 38898 48096 38904
rect 47768 38820 47820 38826
rect 47768 38762 47820 38768
rect 46952 35866 47072 35894
rect 46664 29028 46716 29034
rect 46664 28970 46716 28976
rect 46572 17536 46624 17542
rect 46572 17478 46624 17484
rect 46572 16992 46624 16998
rect 46572 16934 46624 16940
rect 46480 16788 46532 16794
rect 46480 16730 46532 16736
rect 46480 16108 46532 16114
rect 46480 16050 46532 16056
rect 46492 15638 46520 16050
rect 46480 15632 46532 15638
rect 46480 15574 46532 15580
rect 46584 15026 46612 16934
rect 46572 15020 46624 15026
rect 46572 14962 46624 14968
rect 46480 14816 46532 14822
rect 46480 14758 46532 14764
rect 46492 13938 46520 14758
rect 46480 13932 46532 13938
rect 46480 13874 46532 13880
rect 46572 13320 46624 13326
rect 46572 13262 46624 13268
rect 46480 13184 46532 13190
rect 46480 13126 46532 13132
rect 46492 12850 46520 13126
rect 46480 12844 46532 12850
rect 46480 12786 46532 12792
rect 46584 12782 46612 13262
rect 46572 12776 46624 12782
rect 46400 12702 46520 12730
rect 46572 12718 46624 12724
rect 46388 12640 46440 12646
rect 46294 12608 46350 12617
rect 46388 12582 46440 12588
rect 46294 12543 46350 12552
rect 46296 12232 46348 12238
rect 46296 12174 46348 12180
rect 46308 11393 46336 12174
rect 46294 11384 46350 11393
rect 46294 11319 46350 11328
rect 46400 10674 46428 12582
rect 46492 12238 46520 12702
rect 46572 12300 46624 12306
rect 46572 12242 46624 12248
rect 46480 12232 46532 12238
rect 46480 12174 46532 12180
rect 46478 11656 46534 11665
rect 46478 11591 46534 11600
rect 46388 10668 46440 10674
rect 46388 10610 46440 10616
rect 46296 10056 46348 10062
rect 46492 10010 46520 11591
rect 46296 9998 46348 10004
rect 46308 9353 46336 9998
rect 46400 9982 46520 10010
rect 46294 9344 46350 9353
rect 46400 9330 46428 9982
rect 46480 9920 46532 9926
rect 46480 9862 46532 9868
rect 46492 9586 46520 9862
rect 46480 9580 46532 9586
rect 46480 9522 46532 9528
rect 46400 9302 46520 9330
rect 46294 9279 46350 9288
rect 46388 9172 46440 9178
rect 46388 9114 46440 9120
rect 46204 8968 46256 8974
rect 46204 8910 46256 8916
rect 46296 8968 46348 8974
rect 46296 8910 46348 8916
rect 46112 7880 46164 7886
rect 46112 7822 46164 7828
rect 46020 7200 46072 7206
rect 46020 7142 46072 7148
rect 45388 6990 45508 7018
rect 45376 6860 45428 6866
rect 45376 6802 45428 6808
rect 45388 5545 45416 6802
rect 45480 6458 45508 6990
rect 45926 6896 45982 6905
rect 45926 6831 45982 6840
rect 45652 6792 45704 6798
rect 45650 6760 45652 6769
rect 45704 6760 45706 6769
rect 45650 6695 45706 6704
rect 45744 6656 45796 6662
rect 45744 6598 45796 6604
rect 45468 6452 45520 6458
rect 45468 6394 45520 6400
rect 45480 6066 45508 6394
rect 45560 6248 45612 6254
rect 45558 6216 45560 6225
rect 45612 6216 45614 6225
rect 45558 6151 45614 6160
rect 45480 6038 45600 6066
rect 45374 5536 45430 5545
rect 45374 5471 45430 5480
rect 45296 5256 45508 5284
rect 45376 5160 45428 5166
rect 45376 5102 45428 5108
rect 45388 4758 45416 5102
rect 45376 4752 45428 4758
rect 45376 4694 45428 4700
rect 45192 4140 45244 4146
rect 45192 4082 45244 4088
rect 45388 4078 45416 4694
rect 45100 4072 45152 4078
rect 45100 4014 45152 4020
rect 45376 4072 45428 4078
rect 45376 4014 45428 4020
rect 44914 3768 44970 3777
rect 44914 3703 44916 3712
rect 44968 3703 44970 3712
rect 44916 3674 44968 3680
rect 45008 3528 45060 3534
rect 44822 3496 44878 3505
rect 45008 3470 45060 3476
rect 44822 3431 44878 3440
rect 44548 2848 44600 2854
rect 44548 2790 44600 2796
rect 45020 2802 45048 3470
rect 45112 3233 45140 4014
rect 45284 3528 45336 3534
rect 45388 3516 45416 4014
rect 45480 3738 45508 5256
rect 45572 4146 45600 6038
rect 45652 5024 45704 5030
rect 45652 4966 45704 4972
rect 45664 4622 45692 4966
rect 45756 4758 45784 6598
rect 45940 6458 45968 6831
rect 46308 6662 46336 8910
rect 46400 8430 46428 9114
rect 46388 8424 46440 8430
rect 46388 8366 46440 8372
rect 46400 7342 46428 8366
rect 46388 7336 46440 7342
rect 46388 7278 46440 7284
rect 46296 6656 46348 6662
rect 46296 6598 46348 6604
rect 45928 6452 45980 6458
rect 45928 6394 45980 6400
rect 45836 5704 45888 5710
rect 45836 5646 45888 5652
rect 45848 5166 45876 5646
rect 45836 5160 45888 5166
rect 45836 5102 45888 5108
rect 45744 4752 45796 4758
rect 45744 4694 45796 4700
rect 45848 4690 45876 5102
rect 46296 5024 46348 5030
rect 46296 4966 46348 4972
rect 45836 4684 45888 4690
rect 45836 4626 45888 4632
rect 45652 4616 45704 4622
rect 45652 4558 45704 4564
rect 45836 4208 45888 4214
rect 45836 4150 45888 4156
rect 45560 4140 45612 4146
rect 45560 4082 45612 4088
rect 45652 4140 45704 4146
rect 45652 4082 45704 4088
rect 45560 4004 45612 4010
rect 45560 3946 45612 3952
rect 45468 3732 45520 3738
rect 45468 3674 45520 3680
rect 45336 3488 45416 3516
rect 45284 3470 45336 3476
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45098 3224 45154 3233
rect 45098 3159 45154 3168
rect 44456 1352 44508 1358
rect 44456 1294 44508 1300
rect 44560 800 44588 2790
rect 45020 2774 45140 2802
rect 44824 2440 44876 2446
rect 44824 2382 44876 2388
rect 44836 800 44864 2382
rect 45112 800 45140 2774
rect 45388 1850 45416 3334
rect 45480 3058 45508 3674
rect 45572 3398 45600 3946
rect 45664 3777 45692 4082
rect 45744 3936 45796 3942
rect 45744 3878 45796 3884
rect 45650 3768 45706 3777
rect 45650 3703 45706 3712
rect 45652 3528 45704 3534
rect 45652 3470 45704 3476
rect 45560 3392 45612 3398
rect 45560 3334 45612 3340
rect 45664 3233 45692 3470
rect 45650 3224 45706 3233
rect 45650 3159 45706 3168
rect 45560 3120 45612 3126
rect 45560 3062 45612 3068
rect 45468 3052 45520 3058
rect 45468 2994 45520 3000
rect 45572 2961 45600 3062
rect 45558 2952 45614 2961
rect 45558 2887 45614 2896
rect 45388 1822 45508 1850
rect 45480 800 45508 1822
rect 45756 800 45784 3878
rect 45848 3738 45876 4150
rect 46020 4004 46072 4010
rect 46020 3946 46072 3952
rect 45836 3732 45888 3738
rect 45836 3674 45888 3680
rect 45834 3632 45890 3641
rect 45834 3567 45890 3576
rect 45848 3466 45876 3567
rect 45836 3460 45888 3466
rect 45836 3402 45888 3408
rect 46032 800 46060 3946
rect 46308 800 46336 4966
rect 46388 4820 46440 4826
rect 46388 4762 46440 4768
rect 46400 3942 46428 4762
rect 46492 4729 46520 9302
rect 46478 4720 46534 4729
rect 46478 4655 46534 4664
rect 46584 4622 46612 12242
rect 46676 9654 46704 28970
rect 46756 21344 46808 21350
rect 46756 21286 46808 21292
rect 46768 18057 46796 21286
rect 46848 20800 46900 20806
rect 46848 20742 46900 20748
rect 46860 20466 46888 20742
rect 46848 20460 46900 20466
rect 46848 20402 46900 20408
rect 46848 19848 46900 19854
rect 46848 19790 46900 19796
rect 46860 18834 46888 19790
rect 46952 19378 46980 35866
rect 47124 34944 47176 34950
rect 47124 34886 47176 34892
rect 47032 26852 47084 26858
rect 47032 26794 47084 26800
rect 46940 19372 46992 19378
rect 46940 19314 46992 19320
rect 46848 18828 46900 18834
rect 46848 18770 46900 18776
rect 46754 18048 46810 18057
rect 46754 17983 46810 17992
rect 46860 17746 46888 18770
rect 47044 18714 47072 26794
rect 47136 18970 47164 34886
rect 47584 34536 47636 34542
rect 47584 34478 47636 34484
rect 47400 33380 47452 33386
rect 47400 33322 47452 33328
rect 47216 32768 47268 32774
rect 47216 32710 47268 32716
rect 47228 21321 47256 32710
rect 47308 26920 47360 26926
rect 47308 26862 47360 26868
rect 47214 21312 47270 21321
rect 47214 21247 47270 21256
rect 47320 21162 47348 26862
rect 47228 21134 47348 21162
rect 47124 18964 47176 18970
rect 47124 18906 47176 18912
rect 47228 18902 47256 21134
rect 47306 21040 47362 21049
rect 47306 20975 47362 20984
rect 47216 18896 47268 18902
rect 47216 18838 47268 18844
rect 47044 18686 47256 18714
rect 47032 18624 47084 18630
rect 47032 18566 47084 18572
rect 47044 18426 47072 18566
rect 47032 18420 47084 18426
rect 47032 18362 47084 18368
rect 46848 17740 46900 17746
rect 46848 17682 46900 17688
rect 46756 17536 46808 17542
rect 46756 17478 46808 17484
rect 46768 17202 46796 17478
rect 46756 17196 46808 17202
rect 46756 17138 46808 17144
rect 46768 17066 46796 17138
rect 46756 17060 46808 17066
rect 46756 17002 46808 17008
rect 46860 16522 46888 17682
rect 47032 17536 47084 17542
rect 47032 17478 47084 17484
rect 47044 17270 47072 17478
rect 47032 17264 47084 17270
rect 47032 17206 47084 17212
rect 47124 17264 47176 17270
rect 47124 17206 47176 17212
rect 47030 17096 47086 17105
rect 47030 17031 47086 17040
rect 47044 16538 47072 17031
rect 46848 16516 46900 16522
rect 46848 16458 46900 16464
rect 46952 16510 47072 16538
rect 46756 16108 46808 16114
rect 46756 16050 46808 16056
rect 46768 14414 46796 16050
rect 46860 15910 46888 16458
rect 46848 15904 46900 15910
rect 46848 15846 46900 15852
rect 46848 15156 46900 15162
rect 46848 15098 46900 15104
rect 46756 14408 46808 14414
rect 46756 14350 46808 14356
rect 46768 12753 46796 14350
rect 46860 13938 46888 15098
rect 46848 13932 46900 13938
rect 46848 13874 46900 13880
rect 46952 13394 46980 16510
rect 47032 16448 47084 16454
rect 47032 16390 47084 16396
rect 47044 16250 47072 16390
rect 47032 16244 47084 16250
rect 47032 16186 47084 16192
rect 47032 15020 47084 15026
rect 47032 14962 47084 14968
rect 47044 14618 47072 14962
rect 47032 14612 47084 14618
rect 47032 14554 47084 14560
rect 47044 13938 47072 14554
rect 47032 13932 47084 13938
rect 47032 13874 47084 13880
rect 46940 13388 46992 13394
rect 46940 13330 46992 13336
rect 47032 13184 47084 13190
rect 47032 13126 47084 13132
rect 47044 12986 47072 13126
rect 47032 12980 47084 12986
rect 47032 12922 47084 12928
rect 46940 12844 46992 12850
rect 46940 12786 46992 12792
rect 46754 12744 46810 12753
rect 46754 12679 46810 12688
rect 46848 12708 46900 12714
rect 46848 12650 46900 12656
rect 46756 12640 46808 12646
rect 46756 12582 46808 12588
rect 46768 10713 46796 12582
rect 46860 12238 46888 12650
rect 46848 12232 46900 12238
rect 46848 12174 46900 12180
rect 46860 11626 46888 12174
rect 46952 11762 46980 12786
rect 47032 12096 47084 12102
rect 47032 12038 47084 12044
rect 47044 11898 47072 12038
rect 47032 11892 47084 11898
rect 47032 11834 47084 11840
rect 46940 11756 46992 11762
rect 46940 11698 46992 11704
rect 46848 11620 46900 11626
rect 46848 11562 46900 11568
rect 46860 11218 46888 11562
rect 46952 11354 46980 11698
rect 46940 11348 46992 11354
rect 46940 11290 46992 11296
rect 46848 11212 46900 11218
rect 46848 11154 46900 11160
rect 46860 10810 46888 11154
rect 46848 10804 46900 10810
rect 46848 10746 46900 10752
rect 46754 10704 46810 10713
rect 46754 10639 46810 10648
rect 46940 10464 46992 10470
rect 46940 10406 46992 10412
rect 46952 9654 46980 10406
rect 47032 9920 47084 9926
rect 47032 9862 47084 9868
rect 47044 9722 47072 9862
rect 47032 9716 47084 9722
rect 47032 9658 47084 9664
rect 46664 9648 46716 9654
rect 46664 9590 46716 9596
rect 46940 9648 46992 9654
rect 46940 9590 46992 9596
rect 46676 8498 46704 9590
rect 46756 9512 46808 9518
rect 46756 9454 46808 9460
rect 46768 9178 46796 9454
rect 46756 9172 46808 9178
rect 46756 9114 46808 9120
rect 46756 8560 46808 8566
rect 46756 8502 46808 8508
rect 46664 8492 46716 8498
rect 46664 8434 46716 8440
rect 46768 7342 46796 8502
rect 47136 8090 47164 17206
rect 47228 9110 47256 18686
rect 47216 9104 47268 9110
rect 47216 9046 47268 9052
rect 47124 8084 47176 8090
rect 47124 8026 47176 8032
rect 47032 7744 47084 7750
rect 47032 7686 47084 7692
rect 47044 7546 47072 7686
rect 47032 7540 47084 7546
rect 47032 7482 47084 7488
rect 46756 7336 46808 7342
rect 46756 7278 46808 7284
rect 46756 6792 46808 6798
rect 46756 6734 46808 6740
rect 46768 5846 46796 6734
rect 46940 6724 46992 6730
rect 46940 6666 46992 6672
rect 46846 6488 46902 6497
rect 46846 6423 46902 6432
rect 46860 6322 46888 6423
rect 46848 6316 46900 6322
rect 46848 6258 46900 6264
rect 46756 5840 46808 5846
rect 46952 5817 46980 6666
rect 46756 5782 46808 5788
rect 46938 5808 46994 5817
rect 46938 5743 46994 5752
rect 47136 5234 47164 8026
rect 47228 7954 47256 9046
rect 47216 7948 47268 7954
rect 47216 7890 47268 7896
rect 47320 6882 47348 20975
rect 47412 19242 47440 33322
rect 47492 25152 47544 25158
rect 47492 25094 47544 25100
rect 47504 21049 47532 25094
rect 47490 21040 47546 21049
rect 47490 20975 47546 20984
rect 47492 20936 47544 20942
rect 47492 20878 47544 20884
rect 47504 20505 47532 20878
rect 47596 20777 47624 34478
rect 47780 26926 47808 38762
rect 48056 38593 48084 38898
rect 48042 38584 48098 38593
rect 48042 38519 48098 38528
rect 48044 38276 48096 38282
rect 48044 38218 48096 38224
rect 48056 38049 48084 38218
rect 48042 38040 48098 38049
rect 48042 37975 48098 37984
rect 48044 37868 48096 37874
rect 48044 37810 48096 37816
rect 47860 37732 47912 37738
rect 47860 37674 47912 37680
rect 47768 26920 47820 26926
rect 47768 26862 47820 26868
rect 47872 26330 47900 37674
rect 48056 37466 48084 37810
rect 48044 37460 48096 37466
rect 48044 37402 48096 37408
rect 48056 37369 48084 37402
rect 48042 37360 48098 37369
rect 48042 37295 48098 37304
rect 48044 37120 48096 37126
rect 48044 37062 48096 37068
rect 48056 36786 48084 37062
rect 48044 36780 48096 36786
rect 48044 36722 48096 36728
rect 48056 36689 48084 36722
rect 48042 36680 48098 36689
rect 48042 36615 48098 36624
rect 48044 36100 48096 36106
rect 48044 36042 48096 36048
rect 47952 36032 48004 36038
rect 48056 36009 48084 36042
rect 47952 35974 48004 35980
rect 48042 36000 48098 36009
rect 47964 26926 47992 35974
rect 48042 35935 48098 35944
rect 48044 35692 48096 35698
rect 48044 35634 48096 35640
rect 48056 35465 48084 35634
rect 48042 35456 48098 35465
rect 48042 35391 48098 35400
rect 48044 35012 48096 35018
rect 48044 34954 48096 34960
rect 48056 34785 48084 34954
rect 48042 34776 48098 34785
rect 48042 34711 48098 34720
rect 48044 34604 48096 34610
rect 48044 34546 48096 34552
rect 48056 34202 48084 34546
rect 48044 34196 48096 34202
rect 48044 34138 48096 34144
rect 48056 34105 48084 34138
rect 48042 34096 48098 34105
rect 48042 34031 48098 34040
rect 48044 33856 48096 33862
rect 48044 33798 48096 33804
rect 48056 33522 48084 33798
rect 48044 33516 48096 33522
rect 48044 33458 48096 33464
rect 48056 33425 48084 33458
rect 48042 33416 48098 33425
rect 48042 33351 48098 33360
rect 48044 32836 48096 32842
rect 48044 32778 48096 32784
rect 48056 32745 48084 32778
rect 48042 32736 48098 32745
rect 48042 32671 48098 32680
rect 48044 32428 48096 32434
rect 48044 32370 48096 32376
rect 48056 32201 48084 32370
rect 48042 32192 48098 32201
rect 48042 32127 48098 32136
rect 48044 31816 48096 31822
rect 48044 31758 48096 31764
rect 48056 31521 48084 31758
rect 48042 31512 48098 31521
rect 48042 31447 48098 31456
rect 48044 31340 48096 31346
rect 48044 31282 48096 31288
rect 48056 30938 48084 31282
rect 48044 30932 48096 30938
rect 48044 30874 48096 30880
rect 48056 30841 48084 30874
rect 48042 30832 48098 30841
rect 48042 30767 48098 30776
rect 48044 30592 48096 30598
rect 48044 30534 48096 30540
rect 48056 30258 48084 30534
rect 48044 30252 48096 30258
rect 48044 30194 48096 30200
rect 48056 30161 48084 30194
rect 48042 30152 48098 30161
rect 48042 30087 48098 30096
rect 48042 29608 48098 29617
rect 48042 29543 48044 29552
rect 48096 29543 48098 29552
rect 48044 29514 48096 29520
rect 48044 29164 48096 29170
rect 48044 29106 48096 29112
rect 48056 28937 48084 29106
rect 48042 28928 48098 28937
rect 48042 28863 48098 28872
rect 48044 28484 48096 28490
rect 48044 28426 48096 28432
rect 48056 28257 48084 28426
rect 48042 28248 48098 28257
rect 48042 28183 48098 28192
rect 48044 27328 48096 27334
rect 48044 27270 48096 27276
rect 48056 26994 48084 27270
rect 48044 26988 48096 26994
rect 48044 26930 48096 26936
rect 47952 26920 48004 26926
rect 48056 26897 48084 26930
rect 47952 26862 48004 26868
rect 48042 26888 48098 26897
rect 48042 26823 48098 26832
rect 47952 26580 48004 26586
rect 47952 26522 48004 26528
rect 47964 26489 47992 26522
rect 47950 26480 48006 26489
rect 47950 26415 48006 26424
rect 48042 26344 48098 26353
rect 47872 26302 47992 26330
rect 47676 25764 47728 25770
rect 47676 25706 47728 25712
rect 47688 20856 47716 25706
rect 47860 24676 47912 24682
rect 47860 24618 47912 24624
rect 47768 22500 47820 22506
rect 47768 22442 47820 22448
rect 47780 21049 47808 22442
rect 47766 21040 47822 21049
rect 47766 20975 47822 20984
rect 47688 20828 47808 20856
rect 47582 20768 47638 20777
rect 47582 20703 47638 20712
rect 47582 20632 47638 20641
rect 47780 20584 47808 20828
rect 47582 20567 47638 20576
rect 47490 20496 47546 20505
rect 47490 20431 47546 20440
rect 47596 20346 47624 20567
rect 47504 20318 47624 20346
rect 47688 20556 47808 20584
rect 47400 19236 47452 19242
rect 47400 19178 47452 19184
rect 47400 18964 47452 18970
rect 47400 18906 47452 18912
rect 47412 16674 47440 18906
rect 47504 17270 47532 20318
rect 47584 20256 47636 20262
rect 47584 20198 47636 20204
rect 47596 19854 47624 20198
rect 47584 19848 47636 19854
rect 47584 19790 47636 19796
rect 47584 19168 47636 19174
rect 47584 19110 47636 19116
rect 47596 18766 47624 19110
rect 47584 18760 47636 18766
rect 47584 18702 47636 18708
rect 47584 18080 47636 18086
rect 47584 18022 47636 18028
rect 47492 17264 47544 17270
rect 47492 17206 47544 17212
rect 47596 17134 47624 18022
rect 47584 17128 47636 17134
rect 47584 17070 47636 17076
rect 47412 16646 47532 16674
rect 47400 16584 47452 16590
rect 47400 16526 47452 16532
rect 47412 15570 47440 16526
rect 47504 15570 47532 16646
rect 47584 16584 47636 16590
rect 47584 16526 47636 16532
rect 47596 15978 47624 16526
rect 47584 15972 47636 15978
rect 47584 15914 47636 15920
rect 47400 15564 47452 15570
rect 47400 15506 47452 15512
rect 47492 15564 47544 15570
rect 47492 15506 47544 15512
rect 47412 14958 47440 15506
rect 47400 14952 47452 14958
rect 47400 14894 47452 14900
rect 47412 14482 47440 14894
rect 47584 14816 47636 14822
rect 47584 14758 47636 14764
rect 47400 14476 47452 14482
rect 47400 14418 47452 14424
rect 47412 13870 47440 14418
rect 47596 14414 47624 14758
rect 47584 14408 47636 14414
rect 47584 14350 47636 14356
rect 47400 13864 47452 13870
rect 47400 13806 47452 13812
rect 47584 13728 47636 13734
rect 47584 13670 47636 13676
rect 47596 13326 47624 13670
rect 47584 13320 47636 13326
rect 47584 13262 47636 13268
rect 47584 12640 47636 12646
rect 47584 12582 47636 12588
rect 47596 12238 47624 12582
rect 47584 12232 47636 12238
rect 47584 12174 47636 12180
rect 47584 11552 47636 11558
rect 47584 11494 47636 11500
rect 47596 11150 47624 11494
rect 47584 11144 47636 11150
rect 47584 11086 47636 11092
rect 47584 10464 47636 10470
rect 47584 10406 47636 10412
rect 47596 10062 47624 10406
rect 47400 10056 47452 10062
rect 47400 9998 47452 10004
rect 47584 10056 47636 10062
rect 47584 9998 47636 10004
rect 47412 9178 47440 9998
rect 47400 9172 47452 9178
rect 47400 9114 47452 9120
rect 47412 9042 47440 9114
rect 47400 9036 47452 9042
rect 47400 8978 47452 8984
rect 47492 8356 47544 8362
rect 47492 8298 47544 8304
rect 47400 7880 47452 7886
rect 47400 7822 47452 7828
rect 47228 6866 47348 6882
rect 47412 6866 47440 7822
rect 47216 6860 47348 6866
rect 47268 6854 47348 6860
rect 47216 6802 47268 6808
rect 47214 6352 47270 6361
rect 47214 6287 47270 6296
rect 47228 5846 47256 6287
rect 47320 5846 47348 6854
rect 47400 6860 47452 6866
rect 47400 6802 47452 6808
rect 47412 6186 47440 6802
rect 47504 6322 47532 8298
rect 47688 8022 47716 20556
rect 47768 19916 47820 19922
rect 47768 19858 47820 19864
rect 47780 18834 47808 19858
rect 47768 18828 47820 18834
rect 47768 18770 47820 18776
rect 47780 18290 47808 18770
rect 47768 18284 47820 18290
rect 47768 18226 47820 18232
rect 47780 17746 47808 18226
rect 47768 17740 47820 17746
rect 47768 17682 47820 17688
rect 47780 17202 47808 17682
rect 47768 17196 47820 17202
rect 47768 17138 47820 17144
rect 47780 16250 47808 17138
rect 47768 16244 47820 16250
rect 47768 16186 47820 16192
rect 47766 16144 47822 16153
rect 47766 16079 47822 16088
rect 47780 14414 47808 16079
rect 47768 14408 47820 14414
rect 47768 14350 47820 14356
rect 47780 14074 47808 14350
rect 47768 14068 47820 14074
rect 47768 14010 47820 14016
rect 47872 12434 47900 24618
rect 47964 22094 47992 26302
rect 48042 26279 48044 26288
rect 48096 26279 48098 26288
rect 48044 26250 48096 26256
rect 48044 25900 48096 25906
rect 48044 25842 48096 25848
rect 48056 25673 48084 25842
rect 48042 25664 48098 25673
rect 48042 25599 48098 25608
rect 48044 25220 48096 25226
rect 48044 25162 48096 25168
rect 48056 24993 48084 25162
rect 48042 24984 48098 24993
rect 48042 24919 48098 24928
rect 48044 24812 48096 24818
rect 48044 24754 48096 24760
rect 48056 24313 48084 24754
rect 48042 24304 48098 24313
rect 48042 24239 48098 24248
rect 48044 24132 48096 24138
rect 48044 24074 48096 24080
rect 48056 23769 48084 24074
rect 48042 23760 48098 23769
rect 48042 23695 48098 23704
rect 48042 23080 48098 23089
rect 48042 23015 48044 23024
rect 48096 23015 48098 23024
rect 48044 22986 48096 22992
rect 48044 22636 48096 22642
rect 48044 22578 48096 22584
rect 48056 22409 48084 22578
rect 48042 22400 48098 22409
rect 48042 22335 48098 22344
rect 48044 22094 48096 22098
rect 47964 22092 48096 22094
rect 47964 22066 48044 22092
rect 48044 22034 48096 22040
rect 47952 22024 48004 22030
rect 47952 21966 48004 21972
rect 47964 21570 47992 21966
rect 48044 21956 48096 21962
rect 48044 21898 48096 21904
rect 48056 21729 48084 21898
rect 48042 21720 48098 21729
rect 48042 21655 48098 21664
rect 48148 21570 48176 39782
rect 48228 28076 48280 28082
rect 48228 28018 48280 28024
rect 48240 27606 48268 28018
rect 48320 27872 48372 27878
rect 48320 27814 48372 27820
rect 48228 27600 48280 27606
rect 48226 27568 48228 27577
rect 48280 27568 48282 27577
rect 48226 27503 48282 27512
rect 48228 26920 48280 26926
rect 48228 26862 48280 26868
rect 48240 22166 48268 26862
rect 48228 22160 48280 22166
rect 48228 22102 48280 22108
rect 48228 22024 48280 22030
rect 48228 21966 48280 21972
rect 48240 21690 48268 21966
rect 48228 21684 48280 21690
rect 48228 21626 48280 21632
rect 47964 21554 48084 21570
rect 47964 21548 48096 21554
rect 47964 21542 48044 21548
rect 48148 21542 48268 21570
rect 48044 21490 48096 21496
rect 47952 21480 48004 21486
rect 47952 21422 48004 21428
rect 47964 20754 47992 21422
rect 48056 21049 48084 21490
rect 48136 21412 48188 21418
rect 48136 21354 48188 21360
rect 48042 21040 48098 21049
rect 48042 20975 48098 20984
rect 48148 20942 48176 21354
rect 48136 20936 48188 20942
rect 48136 20878 48188 20884
rect 47964 20726 48084 20754
rect 47952 20596 48004 20602
rect 47952 20538 48004 20544
rect 47964 19854 47992 20538
rect 47952 19848 48004 19854
rect 47952 19790 48004 19796
rect 48056 19530 48084 20726
rect 48148 19825 48176 20878
rect 48240 20602 48268 21542
rect 48228 20596 48280 20602
rect 48228 20538 48280 20544
rect 48228 20460 48280 20466
rect 48228 20402 48280 20408
rect 48134 19816 48190 19825
rect 48134 19751 48190 19760
rect 47964 19502 48084 19530
rect 47964 17814 47992 19502
rect 48044 19372 48096 19378
rect 48044 19314 48096 19320
rect 48056 17921 48084 19314
rect 48136 19236 48188 19242
rect 48136 19178 48188 19184
rect 48148 18442 48176 19178
rect 48240 19145 48268 20402
rect 48226 19136 48282 19145
rect 48226 19071 48282 19080
rect 48148 18414 48268 18442
rect 48136 18284 48188 18290
rect 48136 18226 48188 18232
rect 48042 17912 48098 17921
rect 48042 17847 48098 17856
rect 47952 17808 48004 17814
rect 47952 17750 48004 17756
rect 47964 17678 47992 17750
rect 47952 17672 48004 17678
rect 47952 17614 48004 17620
rect 47952 17536 48004 17542
rect 47952 17478 48004 17484
rect 47964 12918 47992 17478
rect 48148 17241 48176 18226
rect 48240 17542 48268 18414
rect 48228 17536 48280 17542
rect 48228 17478 48280 17484
rect 48134 17232 48190 17241
rect 48134 17167 48190 17176
rect 48228 17196 48280 17202
rect 48228 17138 48280 17144
rect 48044 16584 48096 16590
rect 48044 16526 48096 16532
rect 48056 15502 48084 16526
rect 48136 15700 48188 15706
rect 48136 15642 48188 15648
rect 48044 15496 48096 15502
rect 48044 15438 48096 15444
rect 48056 15026 48084 15438
rect 48148 15026 48176 15642
rect 48240 15201 48268 17138
rect 48226 15192 48282 15201
rect 48226 15127 48282 15136
rect 48044 15020 48096 15026
rect 48044 14962 48096 14968
rect 48136 15020 48188 15026
rect 48136 14962 48188 14968
rect 48056 14414 48084 14962
rect 48044 14408 48096 14414
rect 48044 14350 48096 14356
rect 48044 13932 48096 13938
rect 48044 13874 48096 13880
rect 48056 13530 48084 13874
rect 48044 13524 48096 13530
rect 48044 13466 48096 13472
rect 48044 13320 48096 13326
rect 48148 13297 48176 14962
rect 48228 13524 48280 13530
rect 48228 13466 48280 13472
rect 48044 13262 48096 13268
rect 48134 13288 48190 13297
rect 47952 12912 48004 12918
rect 47952 12854 48004 12860
rect 48056 12850 48084 13262
rect 48134 13223 48190 13232
rect 48044 12844 48096 12850
rect 48044 12786 48096 12792
rect 47780 12406 47900 12434
rect 47676 8016 47728 8022
rect 47676 7958 47728 7964
rect 47584 7880 47636 7886
rect 47584 7822 47636 7828
rect 47492 6316 47544 6322
rect 47492 6258 47544 6264
rect 47400 6180 47452 6186
rect 47400 6122 47452 6128
rect 47412 5914 47440 6122
rect 47400 5908 47452 5914
rect 47400 5850 47452 5856
rect 47216 5840 47268 5846
rect 47216 5782 47268 5788
rect 47308 5840 47360 5846
rect 47308 5782 47360 5788
rect 47412 5710 47440 5850
rect 47400 5704 47452 5710
rect 47400 5646 47452 5652
rect 47124 5228 47176 5234
rect 47124 5170 47176 5176
rect 46664 5024 46716 5030
rect 46664 4966 46716 4972
rect 47032 5024 47084 5030
rect 47032 4966 47084 4972
rect 46572 4616 46624 4622
rect 46572 4558 46624 4564
rect 46388 3936 46440 3942
rect 46388 3878 46440 3884
rect 46480 1352 46532 1358
rect 46480 1294 46532 1300
rect 18 0 74 800
rect 110 0 166 800
rect 202 0 258 800
rect 294 0 350 800
rect 386 0 442 800
rect 478 0 534 800
rect 570 0 626 800
rect 662 0 718 800
rect 754 0 810 800
rect 846 0 902 800
rect 938 0 994 800
rect 1030 0 1086 800
rect 1214 0 1270 800
rect 1306 0 1362 800
rect 1398 0 1454 800
rect 1490 0 1546 800
rect 1582 0 1638 800
rect 1674 0 1730 800
rect 1766 0 1822 800
rect 1858 0 1914 800
rect 1950 0 2006 800
rect 2042 0 2098 800
rect 2134 0 2190 800
rect 2226 0 2282 800
rect 2410 0 2466 800
rect 2502 0 2558 800
rect 2594 0 2650 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2870 0 2926 800
rect 2962 0 3018 800
rect 3054 0 3110 800
rect 3146 0 3202 800
rect 3238 0 3294 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3606 0 3662 800
rect 3698 0 3754 800
rect 3790 0 3846 800
rect 3882 0 3938 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4158 0 4214 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4434 0 4490 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4802 0 4858 800
rect 4894 0 4950 800
rect 4986 0 5042 800
rect 5078 0 5134 800
rect 5170 0 5226 800
rect 5262 0 5318 800
rect 5354 0 5410 800
rect 5446 0 5502 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 7010 0 7066 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46492 377 46520 1294
rect 46676 800 46704 4966
rect 46940 4548 46992 4554
rect 46940 4490 46992 4496
rect 46952 4185 46980 4490
rect 46938 4176 46994 4185
rect 46938 4111 46994 4120
rect 46848 2644 46900 2650
rect 46848 2586 46900 2592
rect 46756 2576 46808 2582
rect 46756 2518 46808 2524
rect 46768 1601 46796 2518
rect 46860 2281 46888 2586
rect 47044 2530 47072 4966
rect 47412 4690 47440 5646
rect 47504 5642 47532 6258
rect 47596 6118 47624 7822
rect 47688 6798 47716 7958
rect 47676 6792 47728 6798
rect 47676 6734 47728 6740
rect 47584 6112 47636 6118
rect 47584 6054 47636 6060
rect 47492 5636 47544 5642
rect 47492 5578 47544 5584
rect 47400 4684 47452 4690
rect 47400 4626 47452 4632
rect 47780 4622 47808 12406
rect 48056 12306 48084 12786
rect 48044 12300 48096 12306
rect 48044 12242 48096 12248
rect 48056 11150 48084 12242
rect 48240 12073 48268 13466
rect 48226 12064 48282 12073
rect 48226 11999 48282 12008
rect 48136 11756 48188 11762
rect 48136 11698 48188 11704
rect 48148 11626 48176 11698
rect 48136 11620 48188 11626
rect 48136 11562 48188 11568
rect 48044 11144 48096 11150
rect 48044 11086 48096 11092
rect 48044 10056 48096 10062
rect 48148 10033 48176 11562
rect 48228 10668 48280 10674
rect 48228 10610 48280 10616
rect 48044 9998 48096 10004
rect 48134 10024 48190 10033
rect 48056 9586 48084 9998
rect 48134 9959 48190 9968
rect 48044 9580 48096 9586
rect 48044 9522 48096 9528
rect 48136 9580 48188 9586
rect 48136 9522 48188 9528
rect 47952 9376 48004 9382
rect 47952 9318 48004 9324
rect 47964 7478 47992 9318
rect 48056 8974 48084 9522
rect 48044 8968 48096 8974
rect 48044 8910 48096 8916
rect 48056 8634 48084 8910
rect 48044 8628 48096 8634
rect 48044 8570 48096 8576
rect 48044 7880 48096 7886
rect 48044 7822 48096 7828
rect 47952 7472 48004 7478
rect 47952 7414 48004 7420
rect 47860 7200 47912 7206
rect 47860 7142 47912 7148
rect 47768 4616 47820 4622
rect 47768 4558 47820 4564
rect 47780 4282 47808 4558
rect 47768 4276 47820 4282
rect 47768 4218 47820 4224
rect 47216 4072 47268 4078
rect 47216 4014 47268 4020
rect 47124 3188 47176 3194
rect 47124 3130 47176 3136
rect 46952 2502 47072 2530
rect 46846 2272 46902 2281
rect 46846 2207 46902 2216
rect 46754 1592 46810 1601
rect 46754 1527 46810 1536
rect 46952 800 46980 2502
rect 47136 2446 47164 3130
rect 47124 2440 47176 2446
rect 47124 2382 47176 2388
rect 47228 800 47256 4014
rect 47492 3732 47544 3738
rect 47492 3674 47544 3680
rect 47306 3360 47362 3369
rect 47306 3295 47362 3304
rect 47320 3194 47348 3295
rect 47308 3188 47360 3194
rect 47308 3130 47360 3136
rect 47504 800 47532 3674
rect 47872 800 47900 7142
rect 48056 6798 48084 7822
rect 48148 7449 48176 9522
rect 48240 8809 48268 10610
rect 48332 9042 48360 27814
rect 48412 22160 48464 22166
rect 48412 22102 48464 22108
rect 48424 15094 48452 22102
rect 48412 15088 48464 15094
rect 48412 15030 48464 15036
rect 48320 9036 48372 9042
rect 48320 8978 48372 8984
rect 48226 8800 48282 8809
rect 48226 8735 48282 8744
rect 48134 7440 48190 7449
rect 48134 7375 48190 7384
rect 48044 6792 48096 6798
rect 48044 6734 48096 6740
rect 48056 6458 48084 6734
rect 48044 6452 48096 6458
rect 48044 6394 48096 6400
rect 48056 5710 48084 6394
rect 48044 5704 48096 5710
rect 48044 5646 48096 5652
rect 48056 4622 48084 5646
rect 48044 4616 48096 4622
rect 48044 4558 48096 4564
rect 48688 4140 48740 4146
rect 48688 4082 48740 4088
rect 48136 4004 48188 4010
rect 48136 3946 48188 3952
rect 48148 800 48176 3946
rect 48412 3188 48464 3194
rect 48412 3130 48464 3136
rect 48424 800 48452 3130
rect 48700 800 48728 4082
rect 49792 3936 49844 3942
rect 49792 3878 49844 3884
rect 49148 3664 49200 3670
rect 49148 3606 49200 3612
rect 48964 3596 49016 3602
rect 48964 3538 49016 3544
rect 48976 800 49004 3538
rect 49056 3120 49108 3126
rect 49056 3062 49108 3068
rect 49068 800 49096 3062
rect 49160 800 49188 3606
rect 49516 3392 49568 3398
rect 49516 3334 49568 3340
rect 49332 2848 49384 2854
rect 49332 2790 49384 2796
rect 49240 2304 49292 2310
rect 49240 2246 49292 2252
rect 49252 800 49280 2246
rect 49344 800 49372 2790
rect 49424 2576 49476 2582
rect 49424 2518 49476 2524
rect 49436 800 49464 2518
rect 49528 800 49556 3334
rect 49608 2916 49660 2922
rect 49608 2858 49660 2864
rect 49620 800 49648 2858
rect 49700 2372 49752 2378
rect 49700 2314 49752 2320
rect 49712 800 49740 2314
rect 49804 800 49832 3878
rect 46478 368 46534 377
rect 46478 303 46534 312
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
<< via2 >>
rect 46478 49680 46534 49736
rect 1490 47252 1546 47288
rect 1490 47232 1492 47252
rect 1492 47232 1544 47252
rect 1544 47232 1546 47252
rect 1490 41656 1546 41712
rect 1490 36080 1546 36136
rect 1490 30540 1492 30560
rect 1492 30540 1544 30560
rect 1544 30540 1546 30560
rect 1490 30504 1546 30540
rect 1490 24928 1546 24984
rect 1490 19352 1546 19408
rect 1490 13796 1546 13832
rect 1490 13776 1492 13796
rect 1492 13776 1544 13796
rect 1544 13776 1546 13796
rect 1490 8200 1546 8256
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4526 45484 4582 45520
rect 4526 45464 4528 45484
rect 4528 45464 4580 45484
rect 4580 45464 4582 45484
rect 4894 45464 4950 45520
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 2042 11056 2098 11112
rect 1766 4392 1822 4448
rect 2318 8336 2374 8392
rect 2042 4664 2098 4720
rect 2410 6976 2466 7032
rect 2318 4140 2374 4176
rect 2318 4120 2320 4140
rect 2320 4120 2372 4140
rect 2372 4120 2374 4140
rect 2318 3984 2374 4040
rect 2042 2896 2098 2952
rect 2226 2624 2282 2680
rect 2778 7248 2834 7304
rect 2778 6704 2834 6760
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 2962 8880 3018 8936
rect 3054 6976 3110 7032
rect 3054 3984 3110 4040
rect 2962 3576 3018 3632
rect 2778 3304 2834 3360
rect 2870 3188 2926 3224
rect 2870 3168 2872 3188
rect 2872 3168 2924 3188
rect 2924 3168 2926 3188
rect 2778 2896 2834 2952
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 7194 45484 7250 45520
rect 7194 45464 7196 45484
rect 7196 45464 7248 45484
rect 7248 45464 7250 45484
rect 7746 42508 7748 42528
rect 7748 42508 7800 42528
rect 7800 42508 7802 42528
rect 7746 42472 7802 42508
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 3238 5480 3294 5536
rect 3238 4392 3294 4448
rect 3146 3032 3202 3088
rect 3238 2896 3294 2952
rect 3054 2352 3110 2408
rect 2870 1944 2926 2000
rect 3238 2216 3294 2272
rect 3790 6976 3846 7032
rect 3790 6160 3846 6216
rect 3514 2624 3570 2680
rect 3514 2488 3570 2544
rect 3698 4256 3754 4312
rect 3698 2916 3754 2952
rect 3698 2896 3700 2916
rect 3700 2896 3752 2916
rect 3752 2896 3754 2916
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4158 9424 4214 9480
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4342 8780 4344 8800
rect 4344 8780 4396 8800
rect 4396 8780 4398 8800
rect 4342 8744 4398 8780
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4526 7828 4528 7848
rect 4528 7828 4580 7848
rect 4580 7828 4582 7848
rect 3974 7384 4030 7440
rect 3790 2352 3846 2408
rect 3698 1808 3754 1864
rect 4526 7792 4582 7828
rect 4434 7248 4490 7304
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4342 6840 4398 6896
rect 4342 6332 4344 6352
rect 4344 6332 4396 6352
rect 4396 6332 4398 6352
rect 4342 6296 4398 6332
rect 4250 6160 4306 6216
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4158 5772 4214 5808
rect 4158 5752 4160 5772
rect 4160 5752 4212 5772
rect 4212 5752 4214 5772
rect 4710 8356 4766 8392
rect 4710 8336 4712 8356
rect 4712 8336 4764 8356
rect 4764 8336 4766 8356
rect 4894 8608 4950 8664
rect 4250 5480 4306 5536
rect 4158 5344 4214 5400
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4526 4664 4582 4720
rect 4434 4548 4490 4584
rect 4434 4528 4436 4548
rect 4436 4528 4488 4548
rect 4488 4528 4490 4548
rect 4342 4392 4398 4448
rect 4342 4256 4398 4312
rect 4434 4120 4490 4176
rect 4986 7248 5042 7304
rect 4802 6840 4858 6896
rect 4710 3984 4766 4040
rect 4066 3848 4122 3904
rect 4618 3848 4674 3904
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4250 3304 4306 3360
rect 4526 3440 4582 3496
rect 4434 3188 4490 3224
rect 4434 3168 4436 3188
rect 4436 3168 4488 3188
rect 4488 3168 4490 3188
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4250 2488 4306 2544
rect 3974 1264 4030 1320
rect 5078 6160 5134 6216
rect 4802 992 4858 1048
rect 5078 3168 5134 3224
rect 5354 6840 5410 6896
rect 10230 43696 10286 43752
rect 5630 7248 5686 7304
rect 5538 6704 5594 6760
rect 5446 6024 5502 6080
rect 5354 5072 5410 5128
rect 5170 2760 5226 2816
rect 5170 1128 5226 1184
rect 5446 3168 5502 3224
rect 5722 3304 5778 3360
rect 5906 4276 5962 4312
rect 5906 4256 5908 4276
rect 5908 4256 5960 4276
rect 5960 4256 5962 4276
rect 5814 3168 5870 3224
rect 5722 3032 5778 3088
rect 6182 5480 6238 5536
rect 6090 4664 6146 4720
rect 5998 3304 6054 3360
rect 5814 2488 5870 2544
rect 5998 2760 6054 2816
rect 5630 856 5686 912
rect 6366 2216 6422 2272
rect 7194 7248 7250 7304
rect 6734 5072 6790 5128
rect 6918 5364 6974 5400
rect 6918 5344 6920 5364
rect 6920 5344 6972 5364
rect 6972 5344 6974 5364
rect 6642 3168 6698 3224
rect 7010 3984 7066 4040
rect 7378 5908 7434 5944
rect 7378 5888 7380 5908
rect 7380 5888 7432 5908
rect 7432 5888 7434 5908
rect 7286 5480 7342 5536
rect 7470 5208 7526 5264
rect 7194 2896 7250 2952
rect 6642 1944 6698 2000
rect 7102 2624 7158 2680
rect 6826 2352 6882 2408
rect 7010 2372 7066 2408
rect 7010 2352 7012 2372
rect 7012 2352 7064 2372
rect 7064 2352 7066 2372
rect 7102 1536 7158 1592
rect 7286 1672 7342 1728
rect 7930 6976 7986 7032
rect 7838 4120 7894 4176
rect 8206 6740 8208 6760
rect 8208 6740 8260 6760
rect 8260 6740 8262 6760
rect 8206 6704 8262 6740
rect 8206 5908 8262 5944
rect 8206 5888 8208 5908
rect 8208 5888 8260 5908
rect 8260 5888 8262 5908
rect 8206 5344 8262 5400
rect 8298 4972 8300 4992
rect 8300 4972 8352 4992
rect 8352 4972 8354 4992
rect 8298 4936 8354 4972
rect 8574 4800 8630 4856
rect 8206 4528 8262 4584
rect 7930 3984 7986 4040
rect 7930 3440 7986 3496
rect 8206 4120 8262 4176
rect 8114 3712 8170 3768
rect 7838 2760 7894 2816
rect 7930 2488 7986 2544
rect 8482 4528 8538 4584
rect 8482 4140 8538 4176
rect 8482 4120 8484 4140
rect 8484 4120 8536 4140
rect 8536 4120 8538 4140
rect 8482 3848 8538 3904
rect 8298 2624 8354 2680
rect 9034 6604 9036 6624
rect 9036 6604 9088 6624
rect 9088 6604 9090 6624
rect 9034 6568 9090 6604
rect 9034 5344 9090 5400
rect 8942 4664 8998 4720
rect 8850 4564 8852 4584
rect 8852 4564 8904 4584
rect 8904 4564 8906 4584
rect 8850 4528 8906 4564
rect 8942 4256 8998 4312
rect 8666 3440 8722 3496
rect 9034 3596 9090 3632
rect 9034 3576 9036 3596
rect 9036 3576 9088 3596
rect 9088 3576 9090 3596
rect 8574 2624 8630 2680
rect 8482 2352 8538 2408
rect 8758 3168 8814 3224
rect 9494 6432 9550 6488
rect 9402 4800 9458 4856
rect 9310 4664 9366 4720
rect 9862 4936 9918 4992
rect 9218 4256 9274 4312
rect 10046 5888 10102 5944
rect 10598 6740 10600 6760
rect 10600 6740 10652 6760
rect 10652 6740 10654 6760
rect 10598 6704 10654 6740
rect 10322 6432 10378 6488
rect 9218 3848 9274 3904
rect 9402 3712 9458 3768
rect 9034 2624 9090 2680
rect 9310 3052 9366 3088
rect 9310 3032 9312 3052
rect 9312 3032 9364 3052
rect 9364 3032 9366 3052
rect 8942 1944 8998 2000
rect 9034 1264 9090 1320
rect 10138 5364 10194 5400
rect 10138 5344 10140 5364
rect 10140 5344 10192 5364
rect 10192 5344 10194 5364
rect 10230 4936 10286 4992
rect 10230 4256 10286 4312
rect 10046 3848 10102 3904
rect 9586 3032 9642 3088
rect 10138 3168 10194 3224
rect 9678 2796 9680 2816
rect 9680 2796 9732 2816
rect 9732 2796 9734 2816
rect 9678 2760 9734 2796
rect 10230 2624 10286 2680
rect 9678 2508 9734 2544
rect 10598 6568 10654 6624
rect 11058 6024 11114 6080
rect 10966 5772 11022 5808
rect 10966 5752 10968 5772
rect 10968 5752 11020 5772
rect 11020 5752 11022 5772
rect 10874 5480 10930 5536
rect 10690 4392 10746 4448
rect 10506 3712 10562 3768
rect 10690 4020 10692 4040
rect 10692 4020 10744 4040
rect 10744 4020 10746 4040
rect 10690 3984 10746 4020
rect 9678 2488 9680 2508
rect 9680 2488 9732 2508
rect 9732 2488 9734 2508
rect 9954 2352 10010 2408
rect 10322 2080 10378 2136
rect 10966 4392 11022 4448
rect 11058 4256 11114 4312
rect 10782 2760 10838 2816
rect 10874 2216 10930 2272
rect 11058 3712 11114 3768
rect 11058 3168 11114 3224
rect 11610 6740 11612 6760
rect 11612 6740 11664 6760
rect 11664 6740 11666 6760
rect 11610 6704 11666 6740
rect 11242 2896 11298 2952
rect 11426 4120 11482 4176
rect 11426 3304 11482 3360
rect 11334 2760 11390 2816
rect 11886 5072 11942 5128
rect 11794 2624 11850 2680
rect 11978 4256 12034 4312
rect 11978 2388 11980 2408
rect 11980 2388 12032 2408
rect 12032 2388 12034 2408
rect 11978 2352 12034 2388
rect 12254 5752 12310 5808
rect 12162 4528 12218 4584
rect 12162 3848 12218 3904
rect 12806 3712 12862 3768
rect 12806 3440 12862 3496
rect 12714 3032 12770 3088
rect 13082 3712 13138 3768
rect 12898 2488 12954 2544
rect 13450 3712 13506 3768
rect 13174 2352 13230 2408
rect 14094 4120 14150 4176
rect 15750 43716 15806 43752
rect 15750 43696 15752 43716
rect 15752 43696 15804 43716
rect 15804 43696 15806 43716
rect 14830 3984 14886 4040
rect 15750 4392 15806 4448
rect 16762 5480 16818 5536
rect 16946 4684 17002 4720
rect 16946 4664 16948 4684
rect 16948 4664 17000 4684
rect 17000 4664 17002 4684
rect 17498 43716 17554 43752
rect 17498 43696 17500 43716
rect 17500 43696 17552 43716
rect 17552 43696 17554 43716
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 17774 2624 17830 2680
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 18602 5888 18658 5944
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 22926 43732 22928 43752
rect 22928 43732 22980 43752
rect 22980 43732 22982 43752
rect 22926 43696 22982 43732
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 23386 43696 23442 43752
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 29090 44396 29146 44432
rect 29090 44376 29092 44396
rect 29092 44376 29144 44396
rect 29144 44376 29146 44396
rect 23754 3612 23756 3632
rect 23756 3612 23808 3632
rect 23808 3612 23810 3632
rect 23754 3576 23810 3612
rect 30930 45484 30986 45520
rect 30930 45464 30932 45484
rect 30932 45464 30984 45484
rect 30984 45464 30986 45484
rect 30746 44260 30802 44296
rect 30746 44240 30748 44260
rect 30748 44240 30800 44260
rect 30800 44240 30802 44260
rect 29458 3440 29514 3496
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 31390 44396 31446 44432
rect 31390 44376 31392 44396
rect 31392 44376 31444 44396
rect 31444 44376 31446 44396
rect 31206 44260 31262 44296
rect 31206 44240 31208 44260
rect 31208 44240 31260 44260
rect 31260 44240 31262 44260
rect 29826 3068 29828 3088
rect 29828 3068 29880 3088
rect 29880 3068 29882 3088
rect 29826 3032 29882 3068
rect 30378 3440 30434 3496
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 39946 46416 40002 46472
rect 40498 46572 40554 46608
rect 40498 46552 40500 46572
rect 40500 46552 40552 46572
rect 40552 46552 40554 46572
rect 41050 46280 41106 46336
rect 41786 46572 41842 46608
rect 41786 46552 41788 46572
rect 41788 46552 41840 46572
rect 41840 46552 41842 46572
rect 45650 49000 45706 49056
rect 45098 45484 45154 45520
rect 45098 45464 45100 45484
rect 45100 45464 45152 45484
rect 45152 45464 45154 45484
rect 46202 48320 46258 48376
rect 46018 46280 46074 46336
rect 46662 46416 46718 46472
rect 46846 47132 46848 47152
rect 46848 47132 46900 47152
rect 46900 47132 46902 47152
rect 46846 47096 46902 47132
rect 46846 45056 46902 45112
rect 46846 44376 46902 44432
rect 47306 47640 47362 47696
rect 47858 46416 47914 46472
rect 48042 46436 48098 46472
rect 48042 46416 48044 46436
rect 48044 46416 48096 46436
rect 48096 46416 48098 46436
rect 48042 45772 48044 45792
rect 48044 45772 48096 45792
rect 48096 45772 48098 45792
rect 48042 45736 48098 45772
rect 48042 43832 48098 43888
rect 48042 43172 48098 43208
rect 48042 43152 48044 43172
rect 48044 43152 48096 43172
rect 48096 43152 48098 43172
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 32218 6024 32274 6080
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 43258 6724 43314 6760
rect 43258 6704 43260 6724
rect 43260 6704 43312 6724
rect 43312 6704 43314 6724
rect 44086 6452 44142 6488
rect 44086 6432 44088 6452
rect 44088 6432 44140 6452
rect 44140 6432 44142 6452
rect 40406 3984 40462 4040
rect 41878 3576 41934 3632
rect 42798 3304 42854 3360
rect 42614 856 42670 912
rect 43626 4800 43682 4856
rect 44822 6740 44824 6760
rect 44824 6740 44876 6760
rect 44876 6740 44878 6760
rect 44822 6704 44878 6740
rect 44178 3984 44234 4040
rect 44914 4256 44970 4312
rect 45558 14592 45614 14648
rect 45926 15816 45982 15872
rect 48042 42508 48044 42528
rect 48044 42508 48096 42528
rect 48096 42508 48098 42528
rect 48042 42472 48098 42508
rect 48042 41792 48098 41848
rect 48042 41248 48098 41304
rect 45834 12688 45890 12744
rect 46018 12416 46074 12472
rect 46110 12144 46166 12200
rect 45558 8064 45614 8120
rect 46294 18400 46350 18456
rect 46294 16532 46296 16552
rect 46296 16532 46348 16552
rect 46348 16532 46350 16552
rect 46294 16496 46350 16532
rect 46294 13912 46350 13968
rect 48042 40568 48098 40624
rect 48042 39888 48098 39944
rect 48042 39208 48098 39264
rect 46294 12552 46350 12608
rect 46294 11328 46350 11384
rect 46478 11600 46534 11656
rect 46294 9288 46350 9344
rect 45926 6840 45982 6896
rect 45650 6740 45652 6760
rect 45652 6740 45704 6760
rect 45704 6740 45706 6760
rect 45650 6704 45706 6740
rect 45558 6196 45560 6216
rect 45560 6196 45612 6216
rect 45612 6196 45614 6216
rect 45558 6160 45614 6196
rect 45374 5480 45430 5536
rect 44914 3732 44970 3768
rect 44914 3712 44916 3732
rect 44916 3712 44968 3732
rect 44968 3712 44970 3732
rect 44822 3440 44878 3496
rect 45098 3168 45154 3224
rect 45650 3712 45706 3768
rect 45650 3168 45706 3224
rect 45558 2896 45614 2952
rect 45834 3576 45890 3632
rect 46478 4664 46534 4720
rect 46754 17992 46810 18048
rect 47214 21256 47270 21312
rect 47306 20984 47362 21040
rect 47030 17040 47086 17096
rect 46754 12688 46810 12744
rect 46754 10648 46810 10704
rect 46846 6432 46902 6488
rect 46938 5752 46994 5808
rect 47490 20984 47546 21040
rect 48042 38528 48098 38584
rect 48042 37984 48098 38040
rect 48042 37304 48098 37360
rect 48042 36624 48098 36680
rect 48042 35944 48098 36000
rect 48042 35400 48098 35456
rect 48042 34720 48098 34776
rect 48042 34040 48098 34096
rect 48042 33360 48098 33416
rect 48042 32680 48098 32736
rect 48042 32136 48098 32192
rect 48042 31456 48098 31512
rect 48042 30776 48098 30832
rect 48042 30096 48098 30152
rect 48042 29572 48098 29608
rect 48042 29552 48044 29572
rect 48044 29552 48096 29572
rect 48096 29552 48098 29572
rect 48042 28872 48098 28928
rect 48042 28192 48098 28248
rect 48042 26832 48098 26888
rect 47950 26424 48006 26480
rect 47766 20984 47822 21040
rect 47582 20712 47638 20768
rect 47582 20576 47638 20632
rect 47490 20440 47546 20496
rect 47214 6296 47270 6352
rect 47766 16088 47822 16144
rect 48042 26308 48098 26344
rect 48042 26288 48044 26308
rect 48044 26288 48096 26308
rect 48096 26288 48098 26308
rect 48042 25608 48098 25664
rect 48042 24928 48098 24984
rect 48042 24248 48098 24304
rect 48042 23704 48098 23760
rect 48042 23044 48098 23080
rect 48042 23024 48044 23044
rect 48044 23024 48096 23044
rect 48096 23024 48098 23044
rect 48042 22344 48098 22400
rect 48042 21664 48098 21720
rect 48226 27548 48228 27568
rect 48228 27548 48280 27568
rect 48280 27548 48282 27568
rect 48226 27512 48282 27548
rect 48042 20984 48098 21040
rect 48134 19760 48190 19816
rect 48226 19080 48282 19136
rect 48042 17856 48098 17912
rect 48134 17176 48190 17232
rect 48226 15136 48282 15192
rect 48134 13232 48190 13288
rect 46938 4120 46994 4176
rect 48226 12008 48282 12064
rect 48134 9968 48190 10024
rect 46846 2216 46902 2272
rect 46754 1536 46810 1592
rect 47306 3304 47362 3360
rect 48226 8744 48282 8800
rect 48134 7384 48190 7440
rect 46478 312 46534 368
<< metal3 >>
rect 46473 49738 46539 49741
rect 49200 49738 50000 49768
rect 46473 49736 50000 49738
rect 46473 49680 46478 49736
rect 46534 49680 50000 49736
rect 46473 49678 50000 49680
rect 46473 49675 46539 49678
rect 49200 49648 50000 49678
rect 45645 49058 45711 49061
rect 49200 49058 50000 49088
rect 45645 49056 50000 49058
rect 45645 49000 45650 49056
rect 45706 49000 50000 49056
rect 45645 48998 50000 49000
rect 45645 48995 45711 48998
rect 49200 48968 50000 48998
rect 46197 48378 46263 48381
rect 49200 48378 50000 48408
rect 46197 48376 50000 48378
rect 46197 48320 46202 48376
rect 46258 48320 50000 48376
rect 46197 48318 50000 48320
rect 46197 48315 46263 48318
rect 49200 48288 50000 48318
rect 47301 47698 47367 47701
rect 49200 47698 50000 47728
rect 47301 47696 50000 47698
rect 47301 47640 47306 47696
rect 47362 47640 50000 47696
rect 47301 47638 50000 47640
rect 47301 47635 47367 47638
rect 49200 47608 50000 47638
rect 4208 47360 4528 47361
rect 0 47290 800 47320
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 1485 47290 1551 47293
rect 0 47288 1551 47290
rect 0 47232 1490 47288
rect 1546 47232 1551 47288
rect 0 47230 1551 47232
rect 0 47200 800 47230
rect 1485 47227 1551 47230
rect 46841 47154 46907 47157
rect 49200 47154 50000 47184
rect 46841 47152 50000 47154
rect 46841 47096 46846 47152
rect 46902 47096 50000 47152
rect 46841 47094 50000 47096
rect 46841 47091 46907 47094
rect 49200 47064 50000 47094
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 40493 46610 40559 46613
rect 41781 46610 41847 46613
rect 40493 46608 41847 46610
rect 40493 46552 40498 46608
rect 40554 46552 41786 46608
rect 41842 46552 41847 46608
rect 40493 46550 41847 46552
rect 40493 46547 40559 46550
rect 41781 46547 41847 46550
rect 39941 46474 40007 46477
rect 46657 46474 46723 46477
rect 47853 46474 47919 46477
rect 39941 46472 47919 46474
rect 39941 46416 39946 46472
rect 40002 46416 46662 46472
rect 46718 46416 47858 46472
rect 47914 46416 47919 46472
rect 39941 46414 47919 46416
rect 39941 46411 40007 46414
rect 46657 46411 46723 46414
rect 47853 46411 47919 46414
rect 48037 46474 48103 46477
rect 49200 46474 50000 46504
rect 48037 46472 50000 46474
rect 48037 46416 48042 46472
rect 48098 46416 50000 46472
rect 48037 46414 50000 46416
rect 48037 46411 48103 46414
rect 49200 46384 50000 46414
rect 41045 46338 41111 46341
rect 46013 46338 46079 46341
rect 41045 46336 46079 46338
rect 41045 46280 41050 46336
rect 41106 46280 46018 46336
rect 46074 46280 46079 46336
rect 41045 46278 46079 46280
rect 41045 46275 41111 46278
rect 46013 46275 46079 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 48037 45794 48103 45797
rect 49200 45794 50000 45824
rect 48037 45792 50000 45794
rect 48037 45736 48042 45792
rect 48098 45736 50000 45792
rect 48037 45734 50000 45736
rect 48037 45731 48103 45734
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 49200 45704 50000 45734
rect 19568 45663 19888 45664
rect 4521 45522 4587 45525
rect 4889 45522 4955 45525
rect 7189 45522 7255 45525
rect 4521 45520 7255 45522
rect 4521 45464 4526 45520
rect 4582 45464 4894 45520
rect 4950 45464 7194 45520
rect 7250 45464 7255 45520
rect 4521 45462 7255 45464
rect 4521 45459 4587 45462
rect 4889 45459 4955 45462
rect 7189 45459 7255 45462
rect 30925 45522 30991 45525
rect 45093 45522 45159 45525
rect 30925 45520 45159 45522
rect 30925 45464 30930 45520
rect 30986 45464 45098 45520
rect 45154 45464 45159 45520
rect 30925 45462 45159 45464
rect 30925 45459 30991 45462
rect 45093 45459 45159 45462
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 46841 45114 46907 45117
rect 49200 45114 50000 45144
rect 46841 45112 50000 45114
rect 46841 45056 46846 45112
rect 46902 45056 50000 45112
rect 46841 45054 50000 45056
rect 46841 45051 46907 45054
rect 49200 45024 50000 45054
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 29085 44434 29151 44437
rect 31385 44434 31451 44437
rect 29085 44432 31451 44434
rect 29085 44376 29090 44432
rect 29146 44376 31390 44432
rect 31446 44376 31451 44432
rect 29085 44374 31451 44376
rect 29085 44371 29151 44374
rect 31385 44371 31451 44374
rect 46841 44434 46907 44437
rect 49200 44434 50000 44464
rect 46841 44432 50000 44434
rect 46841 44376 46846 44432
rect 46902 44376 50000 44432
rect 46841 44374 50000 44376
rect 46841 44371 46907 44374
rect 49200 44344 50000 44374
rect 30741 44298 30807 44301
rect 31201 44298 31267 44301
rect 30741 44296 31267 44298
rect 30741 44240 30746 44296
rect 30802 44240 31206 44296
rect 31262 44240 31267 44296
rect 30741 44238 31267 44240
rect 30741 44235 30807 44238
rect 31201 44235 31267 44238
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 48037 43890 48103 43893
rect 49200 43890 50000 43920
rect 48037 43888 50000 43890
rect 48037 43832 48042 43888
rect 48098 43832 50000 43888
rect 48037 43830 50000 43832
rect 48037 43827 48103 43830
rect 49200 43800 50000 43830
rect 10225 43754 10291 43757
rect 15745 43754 15811 43757
rect 17493 43754 17559 43757
rect 10225 43752 17559 43754
rect 10225 43696 10230 43752
rect 10286 43696 15750 43752
rect 15806 43696 17498 43752
rect 17554 43696 17559 43752
rect 10225 43694 17559 43696
rect 10225 43691 10291 43694
rect 15745 43691 15811 43694
rect 17493 43691 17559 43694
rect 22921 43754 22987 43757
rect 23381 43754 23447 43757
rect 22921 43752 23447 43754
rect 22921 43696 22926 43752
rect 22982 43696 23386 43752
rect 23442 43696 23447 43752
rect 22921 43694 23447 43696
rect 22921 43691 22987 43694
rect 23381 43691 23447 43694
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 48037 43210 48103 43213
rect 49200 43210 50000 43240
rect 48037 43208 50000 43210
rect 48037 43152 48042 43208
rect 48098 43152 50000 43208
rect 48037 43150 50000 43152
rect 48037 43147 48103 43150
rect 49200 43120 50000 43150
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 7741 42530 7807 42533
rect 7966 42530 7972 42532
rect 7741 42528 7972 42530
rect 7741 42472 7746 42528
rect 7802 42472 7972 42528
rect 7741 42470 7972 42472
rect 7741 42467 7807 42470
rect 7966 42468 7972 42470
rect 8036 42468 8042 42532
rect 48037 42530 48103 42533
rect 49200 42530 50000 42560
rect 48037 42528 50000 42530
rect 48037 42472 48042 42528
rect 48098 42472 50000 42528
rect 48037 42470 50000 42472
rect 48037 42467 48103 42470
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 49200 42440 50000 42470
rect 19568 42399 19888 42400
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 48037 41850 48103 41853
rect 49200 41850 50000 41880
rect 48037 41848 50000 41850
rect 48037 41792 48042 41848
rect 48098 41792 50000 41848
rect 48037 41790 50000 41792
rect 48037 41787 48103 41790
rect 49200 41760 50000 41790
rect 0 41714 800 41744
rect 1485 41714 1551 41717
rect 0 41712 1551 41714
rect 0 41656 1490 41712
rect 1546 41656 1551 41712
rect 0 41654 1551 41656
rect 0 41624 800 41654
rect 1485 41651 1551 41654
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 48037 41306 48103 41309
rect 49200 41306 50000 41336
rect 48037 41304 50000 41306
rect 48037 41248 48042 41304
rect 48098 41248 50000 41304
rect 48037 41246 50000 41248
rect 48037 41243 48103 41246
rect 49200 41216 50000 41246
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 48037 40626 48103 40629
rect 49200 40626 50000 40656
rect 48037 40624 50000 40626
rect 48037 40568 48042 40624
rect 48098 40568 50000 40624
rect 48037 40566 50000 40568
rect 48037 40563 48103 40566
rect 49200 40536 50000 40566
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 48037 39946 48103 39949
rect 49200 39946 50000 39976
rect 48037 39944 50000 39946
rect 48037 39888 48042 39944
rect 48098 39888 50000 39944
rect 48037 39886 50000 39888
rect 48037 39883 48103 39886
rect 49200 39856 50000 39886
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 48037 39266 48103 39269
rect 49200 39266 50000 39296
rect 48037 39264 50000 39266
rect 48037 39208 48042 39264
rect 48098 39208 50000 39264
rect 48037 39206 50000 39208
rect 48037 39203 48103 39206
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 49200 39176 50000 39206
rect 19568 39135 19888 39136
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 48037 38586 48103 38589
rect 49200 38586 50000 38616
rect 48037 38584 50000 38586
rect 48037 38528 48042 38584
rect 48098 38528 50000 38584
rect 48037 38526 50000 38528
rect 48037 38523 48103 38526
rect 49200 38496 50000 38526
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 48037 38042 48103 38045
rect 49200 38042 50000 38072
rect 48037 38040 50000 38042
rect 48037 37984 48042 38040
rect 48098 37984 50000 38040
rect 48037 37982 50000 37984
rect 48037 37979 48103 37982
rect 49200 37952 50000 37982
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 48037 37362 48103 37365
rect 49200 37362 50000 37392
rect 48037 37360 50000 37362
rect 48037 37304 48042 37360
rect 48098 37304 50000 37360
rect 48037 37302 50000 37304
rect 48037 37299 48103 37302
rect 49200 37272 50000 37302
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 48037 36682 48103 36685
rect 49200 36682 50000 36712
rect 48037 36680 50000 36682
rect 48037 36624 48042 36680
rect 48098 36624 50000 36680
rect 48037 36622 50000 36624
rect 48037 36619 48103 36622
rect 49200 36592 50000 36622
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36138 800 36168
rect 1485 36138 1551 36141
rect 0 36136 1551 36138
rect 0 36080 1490 36136
rect 1546 36080 1551 36136
rect 0 36078 1551 36080
rect 0 36048 800 36078
rect 1485 36075 1551 36078
rect 48037 36002 48103 36005
rect 49200 36002 50000 36032
rect 48037 36000 50000 36002
rect 48037 35944 48042 36000
rect 48098 35944 50000 36000
rect 48037 35942 50000 35944
rect 48037 35939 48103 35942
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 49200 35912 50000 35942
rect 19568 35871 19888 35872
rect 48037 35458 48103 35461
rect 49200 35458 50000 35488
rect 48037 35456 50000 35458
rect 48037 35400 48042 35456
rect 48098 35400 50000 35456
rect 48037 35398 50000 35400
rect 48037 35395 48103 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 49200 35368 50000 35398
rect 34928 35327 35248 35328
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48037 34778 48103 34781
rect 49200 34778 50000 34808
rect 48037 34776 50000 34778
rect 48037 34720 48042 34776
rect 48098 34720 50000 34776
rect 48037 34718 50000 34720
rect 48037 34715 48103 34718
rect 49200 34688 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 48037 34098 48103 34101
rect 49200 34098 50000 34128
rect 48037 34096 50000 34098
rect 48037 34040 48042 34096
rect 48098 34040 50000 34096
rect 48037 34038 50000 34040
rect 48037 34035 48103 34038
rect 49200 34008 50000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 48037 33418 48103 33421
rect 49200 33418 50000 33448
rect 48037 33416 50000 33418
rect 48037 33360 48042 33416
rect 48098 33360 50000 33416
rect 48037 33358 50000 33360
rect 48037 33355 48103 33358
rect 49200 33328 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 48037 32738 48103 32741
rect 49200 32738 50000 32768
rect 48037 32736 50000 32738
rect 48037 32680 48042 32736
rect 48098 32680 50000 32736
rect 48037 32678 50000 32680
rect 48037 32675 48103 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 49200 32648 50000 32678
rect 19568 32607 19888 32608
rect 48037 32194 48103 32197
rect 49200 32194 50000 32224
rect 48037 32192 50000 32194
rect 48037 32136 48042 32192
rect 48098 32136 50000 32192
rect 48037 32134 50000 32136
rect 48037 32131 48103 32134
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 49200 32104 50000 32134
rect 34928 32063 35248 32064
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 48037 31514 48103 31517
rect 49200 31514 50000 31544
rect 48037 31512 50000 31514
rect 48037 31456 48042 31512
rect 48098 31456 50000 31512
rect 48037 31454 50000 31456
rect 48037 31451 48103 31454
rect 49200 31424 50000 31454
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 48037 30834 48103 30837
rect 49200 30834 50000 30864
rect 48037 30832 50000 30834
rect 48037 30776 48042 30832
rect 48098 30776 50000 30832
rect 48037 30774 50000 30776
rect 48037 30771 48103 30774
rect 49200 30744 50000 30774
rect 0 30562 800 30592
rect 1485 30562 1551 30565
rect 0 30560 1551 30562
rect 0 30504 1490 30560
rect 1546 30504 1551 30560
rect 0 30502 1551 30504
rect 0 30472 800 30502
rect 1485 30499 1551 30502
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 48037 30154 48103 30157
rect 49200 30154 50000 30184
rect 48037 30152 50000 30154
rect 48037 30096 48042 30152
rect 48098 30096 50000 30152
rect 48037 30094 50000 30096
rect 48037 30091 48103 30094
rect 49200 30064 50000 30094
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 48037 29610 48103 29613
rect 49200 29610 50000 29640
rect 48037 29608 50000 29610
rect 48037 29552 48042 29608
rect 48098 29552 50000 29608
rect 48037 29550 50000 29552
rect 48037 29547 48103 29550
rect 49200 29520 50000 29550
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 48037 28930 48103 28933
rect 49200 28930 50000 28960
rect 48037 28928 50000 28930
rect 48037 28872 48042 28928
rect 48098 28872 50000 28928
rect 48037 28870 50000 28872
rect 48037 28867 48103 28870
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 49200 28840 50000 28870
rect 34928 28799 35248 28800
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 48037 28250 48103 28253
rect 49200 28250 50000 28280
rect 48037 28248 50000 28250
rect 48037 28192 48042 28248
rect 48098 28192 50000 28248
rect 48037 28190 50000 28192
rect 48037 28187 48103 28190
rect 49200 28160 50000 28190
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 48221 27570 48287 27573
rect 49200 27570 50000 27600
rect 48221 27568 50000 27570
rect 48221 27512 48226 27568
rect 48282 27512 50000 27568
rect 48221 27510 50000 27512
rect 48221 27507 48287 27510
rect 49200 27480 50000 27510
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 48037 26890 48103 26893
rect 49200 26890 50000 26920
rect 48037 26888 50000 26890
rect 48037 26832 48042 26888
rect 48098 26832 50000 26888
rect 48037 26830 50000 26832
rect 48037 26827 48103 26830
rect 49200 26800 50000 26830
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 47945 26482 48011 26485
rect 48078 26482 48084 26484
rect 47945 26480 48084 26482
rect 47945 26424 47950 26480
rect 48006 26424 48084 26480
rect 47945 26422 48084 26424
rect 47945 26419 48011 26422
rect 48078 26420 48084 26422
rect 48148 26420 48154 26484
rect 48037 26346 48103 26349
rect 49200 26346 50000 26376
rect 48037 26344 50000 26346
rect 48037 26288 48042 26344
rect 48098 26288 50000 26344
rect 48037 26286 50000 26288
rect 48037 26283 48103 26286
rect 49200 26256 50000 26286
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 48037 25666 48103 25669
rect 49200 25666 50000 25696
rect 48037 25664 50000 25666
rect 48037 25608 48042 25664
rect 48098 25608 50000 25664
rect 48037 25606 50000 25608
rect 48037 25603 48103 25606
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 49200 25576 50000 25606
rect 34928 25535 35248 25536
rect 19568 25056 19888 25057
rect 0 24986 800 25016
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 1485 24986 1551 24989
rect 0 24984 1551 24986
rect 0 24928 1490 24984
rect 1546 24928 1551 24984
rect 0 24926 1551 24928
rect 0 24896 800 24926
rect 1485 24923 1551 24926
rect 48037 24986 48103 24989
rect 49200 24986 50000 25016
rect 48037 24984 50000 24986
rect 48037 24928 48042 24984
rect 48098 24928 50000 24984
rect 48037 24926 50000 24928
rect 48037 24923 48103 24926
rect 49200 24896 50000 24926
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 48037 24306 48103 24309
rect 49200 24306 50000 24336
rect 48037 24304 50000 24306
rect 48037 24248 48042 24304
rect 48098 24248 50000 24304
rect 48037 24246 50000 24248
rect 48037 24243 48103 24246
rect 49200 24216 50000 24246
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 48037 23762 48103 23765
rect 49200 23762 50000 23792
rect 48037 23760 50000 23762
rect 48037 23704 48042 23760
rect 48098 23704 50000 23760
rect 48037 23702 50000 23704
rect 48037 23699 48103 23702
rect 49200 23672 50000 23702
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 48037 23082 48103 23085
rect 49200 23082 50000 23112
rect 48037 23080 50000 23082
rect 48037 23024 48042 23080
rect 48098 23024 50000 23080
rect 48037 23022 50000 23024
rect 48037 23019 48103 23022
rect 49200 22992 50000 23022
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 48037 22402 48103 22405
rect 49200 22402 50000 22432
rect 48037 22400 50000 22402
rect 48037 22344 48042 22400
rect 48098 22344 50000 22400
rect 48037 22342 50000 22344
rect 48037 22339 48103 22342
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 49200 22312 50000 22342
rect 34928 22271 35248 22272
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 48037 21722 48103 21725
rect 49200 21722 50000 21752
rect 48037 21720 50000 21722
rect 48037 21664 48042 21720
rect 48098 21664 50000 21720
rect 48037 21662 50000 21664
rect 48037 21659 48103 21662
rect 49200 21632 50000 21662
rect 47209 21316 47275 21317
rect 47158 21314 47164 21316
rect 47118 21254 47164 21314
rect 47228 21312 47275 21316
rect 47270 21256 47275 21312
rect 47158 21252 47164 21254
rect 47228 21252 47275 21256
rect 47209 21251 47275 21252
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 47301 21042 47367 21045
rect 47485 21042 47551 21045
rect 47301 21040 47551 21042
rect 47301 20984 47306 21040
rect 47362 20984 47490 21040
rect 47546 20984 47551 21040
rect 47301 20982 47551 20984
rect 47301 20979 47367 20982
rect 47485 20979 47551 20982
rect 47761 21042 47827 21045
rect 48037 21042 48103 21045
rect 49200 21042 50000 21072
rect 47761 21040 47962 21042
rect 47761 20984 47766 21040
rect 47822 20984 47962 21040
rect 47761 20982 47962 20984
rect 47761 20979 47827 20982
rect 47577 20770 47643 20773
rect 47710 20770 47716 20772
rect 47577 20768 47716 20770
rect 47577 20712 47582 20768
rect 47638 20712 47716 20768
rect 47577 20710 47716 20712
rect 47577 20707 47643 20710
rect 47710 20708 47716 20710
rect 47780 20708 47786 20772
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 47577 20634 47643 20637
rect 47902 20634 47962 20982
rect 48037 21040 50000 21042
rect 48037 20984 48042 21040
rect 48098 20984 50000 21040
rect 48037 20982 50000 20984
rect 48037 20979 48103 20982
rect 49200 20952 50000 20982
rect 47577 20632 47962 20634
rect 47577 20576 47582 20632
rect 47638 20576 47962 20632
rect 47577 20574 47962 20576
rect 47577 20571 47643 20574
rect 47485 20498 47551 20501
rect 49200 20498 50000 20528
rect 47485 20496 50000 20498
rect 47485 20440 47490 20496
rect 47546 20440 50000 20496
rect 47485 20438 50000 20440
rect 47485 20435 47551 20438
rect 49200 20408 50000 20438
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 48129 19818 48195 19821
rect 49200 19818 50000 19848
rect 48129 19816 50000 19818
rect 48129 19760 48134 19816
rect 48190 19760 50000 19816
rect 48129 19758 50000 19760
rect 48129 19755 48195 19758
rect 49200 19728 50000 19758
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19410 800 19440
rect 1485 19410 1551 19413
rect 0 19408 1551 19410
rect 0 19352 1490 19408
rect 1546 19352 1551 19408
rect 0 19350 1551 19352
rect 0 19320 800 19350
rect 1485 19347 1551 19350
rect 48221 19138 48287 19141
rect 49200 19138 50000 19168
rect 48221 19136 50000 19138
rect 48221 19080 48226 19136
rect 48282 19080 50000 19136
rect 48221 19078 50000 19080
rect 48221 19075 48287 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 49200 19048 50000 19078
rect 34928 19007 35248 19008
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 46289 18458 46355 18461
rect 49200 18458 50000 18488
rect 46289 18456 50000 18458
rect 46289 18400 46294 18456
rect 46350 18400 50000 18456
rect 46289 18398 50000 18400
rect 46289 18395 46355 18398
rect 49200 18368 50000 18398
rect 46054 17988 46060 18052
rect 46124 18050 46130 18052
rect 46749 18050 46815 18053
rect 46124 18048 46815 18050
rect 46124 17992 46754 18048
rect 46810 17992 46815 18048
rect 46124 17990 46815 17992
rect 46124 17988 46130 17990
rect 46749 17987 46815 17990
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 48037 17914 48103 17917
rect 49200 17914 50000 17944
rect 48037 17912 50000 17914
rect 48037 17856 48042 17912
rect 48098 17856 50000 17912
rect 48037 17854 50000 17856
rect 48037 17851 48103 17854
rect 49200 17824 50000 17854
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 48129 17234 48195 17237
rect 49200 17234 50000 17264
rect 48129 17232 50000 17234
rect 48129 17176 48134 17232
rect 48190 17176 50000 17232
rect 48129 17174 50000 17176
rect 48129 17171 48195 17174
rect 49200 17144 50000 17174
rect 47025 17098 47091 17101
rect 47158 17098 47164 17100
rect 47025 17096 47164 17098
rect 47025 17040 47030 17096
rect 47086 17040 47164 17096
rect 47025 17038 47164 17040
rect 47025 17035 47091 17038
rect 47158 17036 47164 17038
rect 47228 17036 47234 17100
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 46289 16554 46355 16557
rect 49200 16554 50000 16584
rect 46289 16552 50000 16554
rect 46289 16496 46294 16552
rect 46350 16496 50000 16552
rect 46289 16494 50000 16496
rect 46289 16491 46355 16494
rect 49200 16464 50000 16494
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 47761 16148 47827 16149
rect 47710 16084 47716 16148
rect 47780 16146 47827 16148
rect 47780 16144 47872 16146
rect 47822 16088 47872 16144
rect 47780 16086 47872 16088
rect 47780 16084 47827 16086
rect 47761 16083 47827 16084
rect 45921 15874 45987 15877
rect 49200 15874 50000 15904
rect 45921 15872 50000 15874
rect 45921 15816 45926 15872
rect 45982 15816 50000 15872
rect 45921 15814 50000 15816
rect 45921 15811 45987 15814
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 49200 15784 50000 15814
rect 34928 15743 35248 15744
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 48221 15194 48287 15197
rect 49200 15194 50000 15224
rect 48221 15192 50000 15194
rect 48221 15136 48226 15192
rect 48282 15136 50000 15192
rect 48221 15134 50000 15136
rect 48221 15131 48287 15134
rect 49200 15104 50000 15134
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 45553 14650 45619 14653
rect 49200 14650 50000 14680
rect 45553 14648 50000 14650
rect 45553 14592 45558 14648
rect 45614 14592 50000 14648
rect 45553 14590 50000 14592
rect 45553 14587 45619 14590
rect 49200 14560 50000 14590
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 46289 13970 46355 13973
rect 49200 13970 50000 14000
rect 46289 13968 50000 13970
rect 46289 13912 46294 13968
rect 46350 13912 50000 13968
rect 46289 13910 50000 13912
rect 46289 13907 46355 13910
rect 49200 13880 50000 13910
rect 0 13834 800 13864
rect 1485 13834 1551 13837
rect 0 13832 1551 13834
rect 0 13776 1490 13832
rect 1546 13776 1551 13832
rect 0 13774 1551 13776
rect 0 13744 800 13774
rect 1485 13771 1551 13774
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 48129 13290 48195 13293
rect 49200 13290 50000 13320
rect 48129 13288 50000 13290
rect 48129 13232 48134 13288
rect 48190 13232 50000 13288
rect 48129 13230 50000 13232
rect 48129 13227 48195 13230
rect 49200 13200 50000 13230
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 45829 12746 45895 12749
rect 46749 12746 46815 12749
rect 45829 12744 46815 12746
rect 45829 12688 45834 12744
rect 45890 12688 46754 12744
rect 46810 12688 46815 12744
rect 45829 12686 46815 12688
rect 45829 12683 45895 12686
rect 46749 12683 46815 12686
rect 46289 12610 46355 12613
rect 49200 12610 50000 12640
rect 46289 12608 50000 12610
rect 46289 12552 46294 12608
rect 46350 12552 50000 12608
rect 46289 12550 50000 12552
rect 46289 12547 46355 12550
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 49200 12520 50000 12550
rect 34928 12479 35248 12480
rect 46013 12476 46079 12477
rect 46013 12474 46060 12476
rect 45968 12472 46060 12474
rect 45968 12416 46018 12472
rect 45968 12414 46060 12416
rect 46013 12412 46060 12414
rect 46124 12412 46130 12476
rect 46013 12411 46079 12412
rect 46105 12202 46171 12205
rect 46105 12200 46490 12202
rect 46105 12144 46110 12200
rect 46166 12144 46490 12200
rect 46105 12142 46490 12144
rect 46105 12139 46171 12142
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 46430 11661 46490 12142
rect 48221 12066 48287 12069
rect 49200 12066 50000 12096
rect 48221 12064 50000 12066
rect 48221 12008 48226 12064
rect 48282 12008 50000 12064
rect 48221 12006 50000 12008
rect 48221 12003 48287 12006
rect 49200 11976 50000 12006
rect 46430 11656 46539 11661
rect 46430 11600 46478 11656
rect 46534 11600 46539 11656
rect 46430 11598 46539 11600
rect 46473 11595 46539 11598
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 46289 11386 46355 11389
rect 49200 11386 50000 11416
rect 46289 11384 50000 11386
rect 46289 11328 46294 11384
rect 46350 11328 50000 11384
rect 46289 11326 50000 11328
rect 46289 11323 46355 11326
rect 49200 11296 50000 11326
rect 1158 11052 1164 11116
rect 1228 11114 1234 11116
rect 2037 11114 2103 11117
rect 1228 11112 2103 11114
rect 1228 11056 2042 11112
rect 2098 11056 2103 11112
rect 1228 11054 2103 11056
rect 1228 11052 1234 11054
rect 2037 11051 2103 11054
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 46749 10706 46815 10709
rect 49200 10706 50000 10736
rect 46749 10704 50000 10706
rect 46749 10648 46754 10704
rect 46810 10648 50000 10704
rect 46749 10646 50000 10648
rect 46749 10643 46815 10646
rect 49200 10616 50000 10646
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 48129 10026 48195 10029
rect 49200 10026 50000 10056
rect 48129 10024 50000 10026
rect 48129 9968 48134 10024
rect 48190 9968 50000 10024
rect 48129 9966 50000 9968
rect 48129 9963 48195 9966
rect 49200 9936 50000 9966
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 3734 9420 3740 9484
rect 3804 9482 3810 9484
rect 4153 9482 4219 9485
rect 3804 9480 4219 9482
rect 3804 9424 4158 9480
rect 4214 9424 4219 9480
rect 3804 9422 4219 9424
rect 3804 9420 3810 9422
rect 4153 9419 4219 9422
rect 46289 9346 46355 9349
rect 49200 9346 50000 9376
rect 46289 9344 50000 9346
rect 46289 9288 46294 9344
rect 46350 9288 50000 9344
rect 46289 9286 50000 9288
rect 46289 9283 46355 9286
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 49200 9256 50000 9286
rect 34928 9215 35248 9216
rect 2957 8938 3023 8941
rect 4838 8938 4844 8940
rect 2957 8936 4844 8938
rect 2957 8880 2962 8936
rect 3018 8880 4844 8936
rect 2957 8878 4844 8880
rect 2957 8875 3023 8878
rect 4838 8876 4844 8878
rect 4908 8876 4914 8940
rect 3550 8740 3556 8804
rect 3620 8802 3626 8804
rect 4337 8802 4403 8805
rect 3620 8800 4403 8802
rect 3620 8744 4342 8800
rect 4398 8744 4403 8800
rect 3620 8742 4403 8744
rect 3620 8740 3626 8742
rect 4337 8739 4403 8742
rect 48221 8802 48287 8805
rect 49200 8802 50000 8832
rect 48221 8800 50000 8802
rect 48221 8744 48226 8800
rect 48282 8744 50000 8800
rect 48221 8742 50000 8744
rect 48221 8739 48287 8742
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 49200 8712 50000 8742
rect 19568 8671 19888 8672
rect 3918 8604 3924 8668
rect 3988 8666 3994 8668
rect 4889 8666 4955 8669
rect 3988 8664 4955 8666
rect 3988 8608 4894 8664
rect 4950 8608 4955 8664
rect 3988 8606 4955 8608
rect 3988 8604 3994 8606
rect 4889 8603 4955 8606
rect 2313 8396 2379 8397
rect 4705 8396 4771 8397
rect 2262 8332 2268 8396
rect 2332 8394 2379 8396
rect 4654 8394 4660 8396
rect 2332 8392 2424 8394
rect 2374 8336 2424 8392
rect 2332 8334 2424 8336
rect 4614 8334 4660 8394
rect 4724 8392 4771 8396
rect 4766 8336 4771 8392
rect 2332 8332 2379 8334
rect 4654 8332 4660 8334
rect 4724 8332 4771 8336
rect 2313 8331 2379 8332
rect 4705 8331 4771 8332
rect 0 8258 800 8288
rect 1485 8258 1551 8261
rect 0 8256 1551 8258
rect 0 8200 1490 8256
rect 1546 8200 1551 8256
rect 0 8198 1551 8200
rect 0 8168 800 8198
rect 1485 8195 1551 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 45553 8122 45619 8125
rect 49200 8122 50000 8152
rect 45553 8120 50000 8122
rect 45553 8064 45558 8120
rect 45614 8064 50000 8120
rect 45553 8062 50000 8064
rect 45553 8059 45619 8062
rect 49200 8032 50000 8062
rect 2078 7788 2084 7852
rect 2148 7850 2154 7852
rect 4521 7850 4587 7853
rect 2148 7848 4587 7850
rect 2148 7792 4526 7848
rect 4582 7792 4587 7848
rect 2148 7790 4587 7792
rect 2148 7788 2154 7790
rect 4521 7787 4587 7790
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 3969 7442 4035 7445
rect 48129 7442 48195 7445
rect 49200 7442 50000 7472
rect 3969 7440 4722 7442
rect 3969 7384 3974 7440
rect 4030 7384 4722 7440
rect 3969 7382 4722 7384
rect 3969 7379 4035 7382
rect 2773 7308 2839 7309
rect 2773 7304 2820 7308
rect 2884 7306 2890 7308
rect 2773 7248 2778 7304
rect 2773 7244 2820 7248
rect 2884 7246 2930 7306
rect 2884 7244 2890 7246
rect 3366 7244 3372 7308
rect 3436 7306 3442 7308
rect 4429 7306 4495 7309
rect 3436 7304 4495 7306
rect 3436 7248 4434 7304
rect 4490 7248 4495 7304
rect 3436 7246 4495 7248
rect 3436 7244 3442 7246
rect 2773 7243 2839 7244
rect 4429 7243 4495 7246
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 2405 7036 2471 7037
rect 3049 7036 3115 7037
rect 2405 7032 2452 7036
rect 2516 7034 2522 7036
rect 2998 7034 3004 7036
rect 2405 6976 2410 7032
rect 2405 6972 2452 6976
rect 2516 6974 2562 7034
rect 2958 6974 3004 7034
rect 3068 7032 3115 7036
rect 3110 6976 3115 7032
rect 2516 6972 2522 6974
rect 2998 6972 3004 6974
rect 3068 6972 3115 6976
rect 3182 6972 3188 7036
rect 3252 7034 3258 7036
rect 3785 7034 3851 7037
rect 3252 7032 3851 7034
rect 3252 6976 3790 7032
rect 3846 6976 3851 7032
rect 3252 6974 3851 6976
rect 3252 6972 3258 6974
rect 2405 6971 2471 6972
rect 3049 6971 3115 6972
rect 3785 6971 3851 6974
rect 4337 6898 4403 6901
rect 4662 6898 4722 7382
rect 48129 7440 50000 7442
rect 48129 7384 48134 7440
rect 48190 7384 50000 7440
rect 48129 7382 50000 7384
rect 48129 7379 48195 7382
rect 49200 7352 50000 7382
rect 4981 7306 5047 7309
rect 5206 7306 5212 7308
rect 4981 7304 5212 7306
rect 4981 7248 4986 7304
rect 5042 7248 5212 7304
rect 4981 7246 5212 7248
rect 4981 7243 5047 7246
rect 5206 7244 5212 7246
rect 5276 7244 5282 7308
rect 5390 7244 5396 7308
rect 5460 7306 5466 7308
rect 5625 7306 5691 7309
rect 5460 7304 5691 7306
rect 5460 7248 5630 7304
rect 5686 7248 5691 7304
rect 5460 7246 5691 7248
rect 5460 7244 5466 7246
rect 5625 7243 5691 7246
rect 7189 7306 7255 7309
rect 7598 7306 7604 7308
rect 7189 7304 7604 7306
rect 7189 7248 7194 7304
rect 7250 7248 7604 7304
rect 7189 7246 7604 7248
rect 7189 7243 7255 7246
rect 7598 7244 7604 7246
rect 7668 7244 7674 7308
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 7925 7034 7991 7037
rect 8334 7034 8340 7036
rect 7925 7032 8340 7034
rect 7925 6976 7930 7032
rect 7986 6976 8340 7032
rect 7925 6974 8340 6976
rect 7925 6971 7991 6974
rect 8334 6972 8340 6974
rect 8404 6972 8410 7036
rect 4337 6896 4722 6898
rect 4337 6840 4342 6896
rect 4398 6840 4722 6896
rect 4337 6838 4722 6840
rect 4797 6898 4863 6901
rect 5349 6898 5415 6901
rect 45921 6898 45987 6901
rect 4797 6896 45987 6898
rect 4797 6840 4802 6896
rect 4858 6840 5354 6896
rect 5410 6840 45926 6896
rect 45982 6840 45987 6896
rect 4797 6838 45987 6840
rect 4337 6835 4403 6838
rect 4797 6835 4863 6838
rect 5349 6835 5415 6838
rect 45921 6835 45987 6838
rect 2630 6700 2636 6764
rect 2700 6762 2706 6764
rect 2773 6762 2839 6765
rect 5533 6764 5599 6765
rect 5533 6762 5580 6764
rect 2700 6760 2839 6762
rect 2700 6704 2778 6760
rect 2834 6704 2839 6760
rect 2700 6702 2839 6704
rect 5488 6760 5580 6762
rect 5488 6704 5538 6760
rect 5488 6702 5580 6704
rect 2700 6700 2706 6702
rect 2773 6699 2839 6702
rect 5533 6700 5580 6702
rect 5644 6700 5650 6764
rect 7414 6700 7420 6764
rect 7484 6762 7490 6764
rect 8201 6762 8267 6765
rect 7484 6760 8267 6762
rect 7484 6704 8206 6760
rect 8262 6704 8267 6760
rect 7484 6702 8267 6704
rect 7484 6700 7490 6702
rect 5533 6699 5599 6700
rect 8201 6699 8267 6702
rect 9806 6700 9812 6764
rect 9876 6762 9882 6764
rect 10593 6762 10659 6765
rect 9876 6760 10659 6762
rect 9876 6704 10598 6760
rect 10654 6704 10659 6760
rect 9876 6702 10659 6704
rect 9876 6700 9882 6702
rect 10593 6699 10659 6702
rect 11462 6700 11468 6764
rect 11532 6762 11538 6764
rect 11605 6762 11671 6765
rect 11532 6760 11671 6762
rect 11532 6704 11610 6760
rect 11666 6704 11671 6760
rect 11532 6702 11671 6704
rect 11532 6700 11538 6702
rect 11605 6699 11671 6702
rect 43253 6762 43319 6765
rect 44817 6762 44883 6765
rect 43253 6760 44883 6762
rect 43253 6704 43258 6760
rect 43314 6704 44822 6760
rect 44878 6704 44883 6760
rect 43253 6702 44883 6704
rect 43253 6699 43319 6702
rect 44817 6699 44883 6702
rect 45645 6762 45711 6765
rect 49200 6762 50000 6792
rect 45645 6760 50000 6762
rect 45645 6704 45650 6760
rect 45706 6704 50000 6760
rect 45645 6702 50000 6704
rect 45645 6699 45711 6702
rect 49200 6672 50000 6702
rect 5022 6564 5028 6628
rect 5092 6626 5098 6628
rect 9029 6626 9095 6629
rect 10593 6626 10659 6629
rect 5092 6624 10659 6626
rect 5092 6568 9034 6624
rect 9090 6568 10598 6624
rect 10654 6568 10659 6624
rect 5092 6566 10659 6568
rect 5092 6564 5098 6566
rect 9029 6563 9095 6566
rect 10593 6563 10659 6566
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 5942 6428 5948 6492
rect 6012 6490 6018 6492
rect 9489 6490 9555 6493
rect 6012 6488 9555 6490
rect 6012 6432 9494 6488
rect 9550 6432 9555 6488
rect 6012 6430 9555 6432
rect 6012 6428 6018 6430
rect 9489 6427 9555 6430
rect 10174 6428 10180 6492
rect 10244 6490 10250 6492
rect 10317 6490 10383 6493
rect 10244 6488 10383 6490
rect 10244 6432 10322 6488
rect 10378 6432 10383 6488
rect 10244 6430 10383 6432
rect 10244 6428 10250 6430
rect 10317 6427 10383 6430
rect 44081 6490 44147 6493
rect 46841 6490 46907 6493
rect 48078 6490 48084 6492
rect 44081 6488 48084 6490
rect 44081 6432 44086 6488
rect 44142 6432 46846 6488
rect 46902 6432 48084 6488
rect 44081 6430 48084 6432
rect 44081 6427 44147 6430
rect 46841 6427 46907 6430
rect 48078 6428 48084 6430
rect 48148 6428 48154 6492
rect 4337 6354 4403 6357
rect 11094 6354 11100 6356
rect 4337 6352 11100 6354
rect 4337 6296 4342 6352
rect 4398 6296 11100 6352
rect 4337 6294 11100 6296
rect 4337 6291 4403 6294
rect 11094 6292 11100 6294
rect 11164 6292 11170 6356
rect 47209 6354 47275 6357
rect 12390 6352 47275 6354
rect 12390 6296 47214 6352
rect 47270 6296 47275 6352
rect 12390 6294 47275 6296
rect 3785 6218 3851 6221
rect 4245 6218 4311 6221
rect 5073 6218 5139 6221
rect 12390 6218 12450 6294
rect 47209 6291 47275 6294
rect 3785 6216 3986 6218
rect 3785 6160 3790 6216
rect 3846 6160 3986 6216
rect 3785 6158 3986 6160
rect 3785 6155 3851 6158
rect 3926 5674 3986 6158
rect 4245 6216 12450 6218
rect 4245 6160 4250 6216
rect 4306 6160 5078 6216
rect 5134 6160 12450 6216
rect 4245 6158 12450 6160
rect 45553 6218 45619 6221
rect 49200 6218 50000 6248
rect 45553 6216 50000 6218
rect 45553 6160 45558 6216
rect 45614 6160 50000 6216
rect 45553 6158 50000 6160
rect 4245 6155 4311 6158
rect 5073 6155 5139 6158
rect 45553 6155 45619 6158
rect 49200 6128 50000 6158
rect 5206 6020 5212 6084
rect 5276 6082 5282 6084
rect 5441 6082 5507 6085
rect 5276 6080 5507 6082
rect 5276 6024 5446 6080
rect 5502 6024 5507 6080
rect 5276 6022 5507 6024
rect 5276 6020 5282 6022
rect 5441 6019 5507 6022
rect 6862 6020 6868 6084
rect 6932 6082 6938 6084
rect 11053 6082 11119 6085
rect 32213 6082 32279 6085
rect 6932 6022 8264 6082
rect 6932 6020 6938 6022
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 8204 5949 8264 6022
rect 11053 6080 32279 6082
rect 11053 6024 11058 6080
rect 11114 6024 32218 6080
rect 32274 6024 32279 6080
rect 11053 6022 32279 6024
rect 11053 6019 11119 6022
rect 32213 6019 32279 6022
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 7230 5884 7236 5948
rect 7300 5946 7306 5948
rect 7373 5946 7439 5949
rect 7300 5944 7439 5946
rect 7300 5888 7378 5944
rect 7434 5888 7439 5944
rect 7300 5886 7439 5888
rect 7300 5884 7306 5886
rect 7373 5883 7439 5886
rect 8201 5944 8267 5949
rect 8201 5888 8206 5944
rect 8262 5888 8267 5944
rect 8201 5883 8267 5888
rect 10041 5946 10107 5949
rect 18597 5946 18663 5949
rect 10041 5944 18663 5946
rect 10041 5888 10046 5944
rect 10102 5888 18602 5944
rect 18658 5888 18663 5944
rect 10041 5886 18663 5888
rect 10041 5883 10107 5886
rect 18597 5883 18663 5886
rect 4153 5810 4219 5813
rect 5206 5810 5212 5812
rect 4153 5808 5212 5810
rect 4153 5752 4158 5808
rect 4214 5752 5212 5808
rect 4153 5750 5212 5752
rect 4153 5747 4219 5750
rect 5206 5748 5212 5750
rect 5276 5810 5282 5812
rect 9990 5810 9996 5812
rect 5276 5750 9996 5810
rect 5276 5748 5282 5750
rect 9990 5748 9996 5750
rect 10060 5748 10066 5812
rect 10961 5810 11027 5813
rect 12249 5810 12315 5813
rect 46933 5810 46999 5813
rect 10961 5808 12315 5810
rect 10961 5752 10966 5808
rect 11022 5752 12254 5808
rect 12310 5752 12315 5808
rect 10961 5750 12315 5752
rect 10961 5747 11027 5750
rect 12249 5747 12315 5750
rect 12390 5808 46999 5810
rect 12390 5752 46938 5808
rect 46994 5752 46999 5808
rect 12390 5750 46999 5752
rect 12390 5674 12450 5750
rect 46933 5747 46999 5750
rect 3926 5614 12450 5674
rect 3233 5536 3299 5541
rect 3233 5480 3238 5536
rect 3294 5480 3299 5536
rect 3233 5475 3299 5480
rect 3734 5476 3740 5540
rect 3804 5538 3810 5540
rect 4245 5538 4311 5541
rect 6177 5538 6243 5541
rect 3804 5536 6243 5538
rect 3804 5480 4250 5536
rect 4306 5480 6182 5536
rect 6238 5480 6243 5536
rect 3804 5478 6243 5480
rect 3804 5476 3810 5478
rect 4245 5475 4311 5478
rect 6177 5475 6243 5478
rect 6494 5476 6500 5540
rect 6564 5538 6570 5540
rect 7281 5538 7347 5541
rect 10869 5538 10935 5541
rect 16757 5538 16823 5541
rect 6564 5536 7347 5538
rect 6564 5480 7286 5536
rect 7342 5480 7347 5536
rect 6564 5478 7347 5480
rect 6564 5476 6570 5478
rect 7281 5475 7347 5478
rect 10366 5536 10935 5538
rect 10366 5480 10874 5536
rect 10930 5480 10935 5536
rect 10366 5478 10935 5480
rect 2037 4722 2103 4725
rect 1902 4720 2103 4722
rect 1902 4664 2042 4720
rect 2098 4664 2103 4720
rect 1902 4662 2103 4664
rect 1761 4450 1827 4453
rect 1902 4450 1962 4662
rect 2037 4659 2103 4662
rect 3236 4453 3296 5475
rect 4153 5400 4219 5405
rect 4153 5344 4158 5400
rect 4214 5344 4219 5400
rect 4153 5339 4219 5344
rect 5574 5340 5580 5404
rect 5644 5402 5650 5404
rect 6913 5402 6979 5405
rect 5644 5400 7666 5402
rect 5644 5344 6918 5400
rect 6974 5344 7666 5400
rect 5644 5342 7666 5344
rect 5644 5340 5650 5342
rect 6913 5339 6979 5342
rect 4156 5130 4216 5339
rect 5206 5266 5212 5268
rect 5030 5206 5212 5266
rect 4156 5070 4722 5130
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 4521 4722 4587 4725
rect 4662 4722 4722 5070
rect 4521 4720 4722 4722
rect 4521 4664 4526 4720
rect 4582 4664 4722 4720
rect 4521 4662 4722 4664
rect 4521 4659 4587 4662
rect 3550 4524 3556 4588
rect 3620 4586 3626 4588
rect 4429 4586 4495 4589
rect 3620 4584 4495 4586
rect 3620 4528 4434 4584
rect 4490 4528 4495 4584
rect 3620 4526 4495 4528
rect 3620 4524 3626 4526
rect 4429 4523 4495 4526
rect 1761 4448 1962 4450
rect 1761 4392 1766 4448
rect 1822 4392 1962 4448
rect 1761 4390 1962 4392
rect 3233 4448 3299 4453
rect 3233 4392 3238 4448
rect 3294 4392 3299 4448
rect 1761 4387 1827 4390
rect 3233 4387 3299 4392
rect 3734 4388 3740 4452
rect 3804 4450 3810 4452
rect 4337 4450 4403 4453
rect 3804 4448 4403 4450
rect 3804 4392 4342 4448
rect 4398 4392 4403 4448
rect 3804 4390 4403 4392
rect 3804 4388 3810 4390
rect 4337 4387 4403 4390
rect 3693 4312 3759 4317
rect 3693 4256 3698 4312
rect 3754 4256 3759 4312
rect 3693 4251 3759 4256
rect 4337 4314 4403 4317
rect 5030 4314 5090 5206
rect 5206 5204 5212 5206
rect 5276 5204 5282 5268
rect 7046 5204 7052 5268
rect 7116 5266 7122 5268
rect 7465 5266 7531 5269
rect 7116 5264 7531 5266
rect 7116 5208 7470 5264
rect 7526 5208 7531 5264
rect 7116 5206 7531 5208
rect 7606 5266 7666 5342
rect 7782 5340 7788 5404
rect 7852 5402 7858 5404
rect 8201 5402 8267 5405
rect 7852 5400 8267 5402
rect 7852 5344 8206 5400
rect 8262 5344 8267 5400
rect 7852 5342 8267 5344
rect 7852 5340 7858 5342
rect 8201 5339 8267 5342
rect 8518 5340 8524 5404
rect 8588 5402 8594 5404
rect 9029 5402 9095 5405
rect 8588 5400 9095 5402
rect 8588 5344 9034 5400
rect 9090 5344 9095 5400
rect 8588 5342 9095 5344
rect 8588 5340 8594 5342
rect 9029 5339 9095 5342
rect 10133 5402 10199 5405
rect 10366 5402 10426 5478
rect 10869 5475 10935 5478
rect 12390 5536 16823 5538
rect 12390 5480 16762 5536
rect 16818 5480 16823 5536
rect 12390 5478 16823 5480
rect 10133 5400 10426 5402
rect 10133 5344 10138 5400
rect 10194 5344 10426 5400
rect 10133 5342 10426 5344
rect 10133 5339 10199 5342
rect 12390 5266 12450 5478
rect 16757 5475 16823 5478
rect 45369 5538 45435 5541
rect 49200 5538 50000 5568
rect 45369 5536 50000 5538
rect 45369 5480 45374 5536
rect 45430 5480 50000 5536
rect 45369 5478 50000 5480
rect 45369 5475 45435 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 49200 5448 50000 5478
rect 19568 5407 19888 5408
rect 7606 5206 12450 5266
rect 7116 5204 7122 5206
rect 7465 5203 7531 5206
rect 5206 5068 5212 5132
rect 5276 5130 5282 5132
rect 5349 5130 5415 5133
rect 6729 5132 6795 5133
rect 6678 5130 6684 5132
rect 5276 5128 5415 5130
rect 5276 5072 5354 5128
rect 5410 5072 5415 5128
rect 5276 5070 5415 5072
rect 6638 5070 6684 5130
rect 6748 5128 6795 5132
rect 11881 5130 11947 5133
rect 6790 5072 6795 5128
rect 5276 5068 5282 5070
rect 5349 5067 5415 5070
rect 6678 5068 6684 5070
rect 6748 5068 6795 5072
rect 6729 5067 6795 5068
rect 9630 5128 11947 5130
rect 9630 5072 11886 5128
rect 11942 5072 11947 5128
rect 9630 5070 11947 5072
rect 8293 4994 8359 4997
rect 9630 4994 9690 5070
rect 11881 5067 11947 5070
rect 8293 4992 9690 4994
rect 8293 4936 8298 4992
rect 8354 4936 9690 4992
rect 8293 4934 9690 4936
rect 9857 4994 9923 4997
rect 10225 4994 10291 4997
rect 9857 4992 10291 4994
rect 9857 4936 9862 4992
rect 9918 4936 10230 4992
rect 10286 4936 10291 4992
rect 9857 4934 10291 4936
rect 8293 4931 8359 4934
rect 9857 4931 9923 4934
rect 10225 4931 10291 4934
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 8150 4796 8156 4860
rect 8220 4858 8226 4860
rect 8569 4858 8635 4861
rect 8220 4856 8635 4858
rect 8220 4800 8574 4856
rect 8630 4800 8635 4856
rect 8220 4798 8635 4800
rect 8220 4796 8226 4798
rect 8569 4795 8635 4798
rect 9254 4796 9260 4860
rect 9324 4858 9330 4860
rect 9397 4858 9463 4861
rect 9324 4856 9463 4858
rect 9324 4800 9402 4856
rect 9458 4800 9463 4856
rect 9324 4798 9463 4800
rect 9324 4796 9330 4798
rect 9397 4795 9463 4798
rect 43621 4858 43687 4861
rect 49200 4858 50000 4888
rect 43621 4856 50000 4858
rect 43621 4800 43626 4856
rect 43682 4800 50000 4856
rect 43621 4798 50000 4800
rect 43621 4795 43687 4798
rect 49200 4768 50000 4798
rect 6085 4722 6151 4725
rect 8937 4722 9003 4725
rect 5904 4720 6151 4722
rect 5904 4664 6090 4720
rect 6146 4664 6151 4720
rect 5904 4662 6151 4664
rect 5904 4317 5964 4662
rect 6085 4659 6151 4662
rect 8296 4720 9003 4722
rect 8296 4664 8942 4720
rect 8998 4664 9003 4720
rect 8296 4662 9003 4664
rect 8296 4620 8356 4662
rect 8937 4659 9003 4662
rect 9070 4660 9076 4724
rect 9140 4722 9146 4724
rect 9305 4722 9371 4725
rect 9140 4720 9371 4722
rect 9140 4664 9310 4720
rect 9366 4664 9371 4720
rect 9140 4662 9371 4664
rect 9140 4660 9146 4662
rect 9305 4659 9371 4662
rect 11094 4660 11100 4724
rect 11164 4722 11170 4724
rect 16941 4722 17007 4725
rect 46473 4722 46539 4725
rect 11164 4662 12450 4722
rect 11164 4660 11170 4662
rect 8204 4589 8356 4620
rect 8201 4584 8356 4589
rect 8201 4528 8206 4584
rect 8262 4560 8356 4584
rect 8477 4586 8543 4589
rect 8702 4586 8708 4588
rect 8477 4584 8708 4586
rect 8262 4528 8267 4560
rect 8201 4523 8267 4528
rect 8477 4528 8482 4584
rect 8538 4528 8708 4584
rect 8477 4526 8708 4528
rect 8477 4523 8543 4526
rect 8702 4524 8708 4526
rect 8772 4586 8778 4588
rect 8845 4586 8911 4589
rect 12157 4586 12223 4589
rect 8772 4584 12223 4586
rect 8772 4528 8850 4584
rect 8906 4528 12162 4584
rect 12218 4528 12223 4584
rect 8772 4526 12223 4528
rect 12390 4586 12450 4662
rect 16941 4720 46539 4722
rect 16941 4664 16946 4720
rect 17002 4664 46478 4720
rect 46534 4664 46539 4720
rect 16941 4662 46539 4664
rect 16941 4659 17007 4662
rect 46473 4659 46539 4662
rect 12390 4526 22110 4586
rect 8772 4524 8778 4526
rect 8845 4523 8911 4526
rect 12157 4523 12223 4526
rect 8886 4388 8892 4452
rect 8956 4450 8962 4452
rect 10685 4450 10751 4453
rect 10961 4452 11027 4453
rect 10910 4450 10916 4452
rect 8956 4448 10751 4450
rect 8956 4392 10690 4448
rect 10746 4392 10751 4448
rect 8956 4390 10751 4392
rect 10870 4390 10916 4450
rect 10980 4448 11027 4452
rect 11022 4392 11027 4448
rect 8956 4388 8962 4390
rect 10685 4387 10751 4390
rect 10910 4388 10916 4390
rect 10980 4388 11027 4392
rect 11094 4388 11100 4452
rect 11164 4450 11170 4452
rect 15745 4450 15811 4453
rect 11164 4448 15811 4450
rect 11164 4392 15750 4448
rect 15806 4392 15811 4448
rect 11164 4390 15811 4392
rect 11164 4388 11170 4390
rect 10961 4387 11027 4388
rect 15745 4387 15811 4390
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 4337 4312 5090 4314
rect 4337 4256 4342 4312
rect 4398 4256 5090 4312
rect 4337 4254 5090 4256
rect 4337 4251 4403 4254
rect 5758 4252 5764 4316
rect 5828 4314 5834 4316
rect 5901 4314 5967 4317
rect 5828 4312 5967 4314
rect 5828 4256 5906 4312
rect 5962 4256 5967 4312
rect 5828 4254 5967 4256
rect 5828 4252 5834 4254
rect 5901 4251 5967 4254
rect 8937 4314 9003 4317
rect 9213 4314 9279 4317
rect 8937 4312 9279 4314
rect 8937 4256 8942 4312
rect 8998 4256 9218 4312
rect 9274 4256 9279 4312
rect 8937 4254 9279 4256
rect 8937 4251 9003 4254
rect 9213 4251 9279 4254
rect 9438 4252 9444 4316
rect 9508 4314 9514 4316
rect 10225 4314 10291 4317
rect 9508 4312 10291 4314
rect 9508 4256 10230 4312
rect 10286 4256 10291 4312
rect 9508 4254 10291 4256
rect 9508 4252 9514 4254
rect 10225 4251 10291 4254
rect 11053 4314 11119 4317
rect 11973 4314 12039 4317
rect 11053 4312 12039 4314
rect 11053 4256 11058 4312
rect 11114 4256 11978 4312
rect 12034 4256 12039 4312
rect 11053 4254 12039 4256
rect 11053 4251 11119 4254
rect 11973 4251 12039 4254
rect 2313 4180 2379 4181
rect 2262 4178 2268 4180
rect 2222 4118 2268 4178
rect 2332 4176 2379 4180
rect 2374 4120 2379 4176
rect 2262 4116 2268 4118
rect 2332 4116 2379 4120
rect 2313 4115 2379 4116
rect 2313 4042 2379 4045
rect 3049 4044 3115 4045
rect 2446 4042 2452 4044
rect 2313 4040 2452 4042
rect 2313 3984 2318 4040
rect 2374 3984 2452 4040
rect 2313 3982 2452 3984
rect 2313 3979 2379 3982
rect 2446 3980 2452 3982
rect 2516 3980 2522 4044
rect 2998 3980 3004 4044
rect 3068 4042 3115 4044
rect 3068 4040 3160 4042
rect 3110 3984 3160 4040
rect 3068 3982 3160 3984
rect 3068 3980 3115 3982
rect 3049 3979 3115 3980
rect 2998 3844 3004 3908
rect 3068 3906 3074 3908
rect 3696 3906 3756 4251
rect 4429 4178 4495 4181
rect 5574 4178 5580 4180
rect 4429 4176 5580 4178
rect 4429 4120 4434 4176
rect 4490 4120 5580 4176
rect 4429 4118 5580 4120
rect 4429 4115 4495 4118
rect 5574 4116 5580 4118
rect 5644 4116 5650 4180
rect 6310 4116 6316 4180
rect 6380 4178 6386 4180
rect 7833 4178 7899 4181
rect 6380 4176 7899 4178
rect 6380 4120 7838 4176
rect 7894 4120 7899 4176
rect 6380 4118 7899 4120
rect 6380 4116 6386 4118
rect 7833 4115 7899 4118
rect 8201 4178 8267 4181
rect 8334 4178 8340 4180
rect 8201 4176 8340 4178
rect 8201 4120 8206 4176
rect 8262 4120 8340 4176
rect 8201 4118 8340 4120
rect 8201 4115 8267 4118
rect 8334 4116 8340 4118
rect 8404 4178 8410 4180
rect 8477 4178 8543 4181
rect 8404 4176 8543 4178
rect 8404 4120 8482 4176
rect 8538 4120 8543 4176
rect 8404 4118 8543 4120
rect 8404 4116 8410 4118
rect 8477 4115 8543 4118
rect 11421 4178 11487 4181
rect 14089 4178 14155 4181
rect 11421 4176 14155 4178
rect 11421 4120 11426 4176
rect 11482 4120 14094 4176
rect 14150 4120 14155 4176
rect 11421 4118 14155 4120
rect 22050 4178 22110 4526
rect 44909 4314 44975 4317
rect 44909 4312 47226 4314
rect 44909 4256 44914 4312
rect 44970 4256 47226 4312
rect 44909 4254 47226 4256
rect 44909 4251 44975 4254
rect 46933 4178 46999 4181
rect 22050 4176 46999 4178
rect 22050 4120 46938 4176
rect 46994 4120 46999 4176
rect 22050 4118 46999 4120
rect 47166 4178 47226 4254
rect 49200 4178 50000 4208
rect 47166 4118 50000 4178
rect 11421 4115 11487 4118
rect 14089 4115 14155 4118
rect 46933 4115 46999 4118
rect 49200 4088 50000 4118
rect 4705 4044 4771 4045
rect 4654 3980 4660 4044
rect 4724 4042 4771 4044
rect 7005 4042 7071 4045
rect 7925 4044 7991 4045
rect 7230 4042 7236 4044
rect 4724 4040 4816 4042
rect 4766 3984 4816 4040
rect 4724 3982 4816 3984
rect 7005 4040 7236 4042
rect 7005 3984 7010 4040
rect 7066 3984 7236 4040
rect 7005 3982 7236 3984
rect 4724 3980 4771 3982
rect 4705 3979 4771 3980
rect 7005 3979 7071 3982
rect 7230 3980 7236 3982
rect 7300 3980 7306 4044
rect 7925 4040 7972 4044
rect 8036 4042 8042 4044
rect 9400 4042 9690 4076
rect 10174 4042 10180 4044
rect 7925 3984 7930 4040
rect 7925 3980 7972 3984
rect 8036 3982 8082 4042
rect 8158 4016 10180 4042
rect 8158 3982 9460 4016
rect 9630 3982 10180 4016
rect 8036 3980 8042 3982
rect 7925 3979 7991 3980
rect 3068 3846 3756 3906
rect 3068 3844 3074 3846
rect 3918 3844 3924 3908
rect 3988 3906 3994 3908
rect 4061 3906 4127 3909
rect 3988 3904 4127 3906
rect 3988 3848 4066 3904
rect 4122 3848 4127 3904
rect 3988 3846 4127 3848
rect 3988 3844 3994 3846
rect 4061 3843 4127 3846
rect 4613 3908 4679 3909
rect 4613 3904 4660 3908
rect 4724 3906 4730 3908
rect 4613 3848 4618 3904
rect 4613 3844 4660 3848
rect 4724 3846 4770 3906
rect 4724 3844 4730 3846
rect 6126 3844 6132 3908
rect 6196 3906 6202 3908
rect 8158 3906 8218 3982
rect 10174 3980 10180 3982
rect 10244 3980 10250 4044
rect 10685 4042 10751 4045
rect 14825 4042 14891 4045
rect 10685 4040 14891 4042
rect 10685 3984 10690 4040
rect 10746 3984 14830 4040
rect 14886 3984 14891 4040
rect 10685 3982 14891 3984
rect 6196 3846 8218 3906
rect 8477 3906 8543 3909
rect 9213 3906 9279 3909
rect 10041 3906 10107 3909
rect 8477 3904 9279 3906
rect 8477 3848 8482 3904
rect 8538 3848 9218 3904
rect 9274 3848 9279 3904
rect 8477 3846 9279 3848
rect 6196 3844 6202 3846
rect 4613 3843 4679 3844
rect 8477 3843 8543 3846
rect 9213 3843 9279 3846
rect 9446 3904 10107 3906
rect 9446 3848 10046 3904
rect 10102 3848 10107 3904
rect 9446 3846 10107 3848
rect 10182 3906 10242 3980
rect 10685 3979 10751 3982
rect 14825 3979 14891 3982
rect 40401 4042 40467 4045
rect 44173 4042 44239 4045
rect 40401 4040 44239 4042
rect 40401 3984 40406 4040
rect 40462 3984 44178 4040
rect 44234 3984 44239 4040
rect 40401 3982 44239 3984
rect 40401 3979 40467 3982
rect 44173 3979 44239 3982
rect 10182 3846 11300 3906
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 9446 3773 9506 3846
rect 10041 3843 10107 3846
rect 8109 3770 8175 3773
rect 8518 3770 8524 3772
rect 8109 3768 8524 3770
rect 8109 3712 8114 3768
rect 8170 3712 8524 3768
rect 8109 3710 8524 3712
rect 8109 3707 8175 3710
rect 8518 3708 8524 3710
rect 8588 3708 8594 3772
rect 9397 3768 9506 3773
rect 9397 3712 9402 3768
rect 9458 3712 9506 3768
rect 9397 3710 9506 3712
rect 10501 3770 10567 3773
rect 11053 3770 11119 3773
rect 10501 3768 11119 3770
rect 10501 3712 10506 3768
rect 10562 3712 11058 3768
rect 11114 3712 11119 3768
rect 10501 3710 11119 3712
rect 11240 3770 11300 3846
rect 12014 3844 12020 3908
rect 12084 3906 12090 3908
rect 12157 3906 12223 3909
rect 12084 3904 12223 3906
rect 12084 3848 12162 3904
rect 12218 3848 12223 3904
rect 12084 3846 12223 3848
rect 12084 3844 12090 3846
rect 12157 3843 12223 3846
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 12801 3770 12867 3773
rect 11240 3768 12867 3770
rect 11240 3712 12806 3768
rect 12862 3712 12867 3768
rect 11240 3710 12867 3712
rect 9397 3707 9463 3710
rect 10501 3707 10567 3710
rect 11053 3707 11119 3710
rect 12801 3707 12867 3710
rect 13077 3770 13143 3773
rect 13445 3770 13511 3773
rect 13077 3768 13511 3770
rect 13077 3712 13082 3768
rect 13138 3712 13450 3768
rect 13506 3712 13511 3768
rect 13077 3710 13511 3712
rect 13077 3707 13143 3710
rect 13445 3707 13511 3710
rect 44909 3770 44975 3773
rect 45645 3770 45711 3773
rect 44909 3768 45711 3770
rect 44909 3712 44914 3768
rect 44970 3712 45650 3768
rect 45706 3712 45711 3768
rect 44909 3710 45711 3712
rect 44909 3707 44975 3710
rect 45645 3707 45711 3710
rect 2957 3634 3023 3637
rect 5022 3634 5028 3636
rect 2957 3632 5028 3634
rect 2957 3576 2962 3632
rect 3018 3576 5028 3632
rect 2957 3574 5028 3576
rect 2957 3571 3023 3574
rect 5022 3572 5028 3574
rect 5092 3572 5098 3636
rect 8334 3572 8340 3636
rect 8404 3634 8410 3636
rect 9029 3634 9095 3637
rect 23749 3634 23815 3637
rect 8404 3574 8954 3634
rect 8404 3572 8410 3574
rect 4521 3498 4587 3501
rect 4838 3498 4844 3500
rect 4521 3496 4844 3498
rect 4521 3440 4526 3496
rect 4582 3440 4844 3496
rect 4521 3438 4844 3440
rect 4521 3435 4587 3438
rect 4838 3436 4844 3438
rect 4908 3436 4914 3500
rect 7925 3498 7991 3501
rect 8661 3498 8727 3501
rect 7925 3496 8727 3498
rect 7925 3440 7930 3496
rect 7986 3440 8666 3496
rect 8722 3440 8727 3496
rect 7925 3438 8727 3440
rect 8894 3498 8954 3574
rect 9029 3632 23815 3634
rect 9029 3576 9034 3632
rect 9090 3576 23754 3632
rect 23810 3576 23815 3632
rect 9029 3574 23815 3576
rect 9029 3571 9095 3574
rect 23749 3571 23815 3574
rect 41873 3634 41939 3637
rect 45829 3634 45895 3637
rect 41873 3632 45895 3634
rect 41873 3576 41878 3632
rect 41934 3576 45834 3632
rect 45890 3576 45895 3632
rect 41873 3574 45895 3576
rect 41873 3571 41939 3574
rect 45829 3571 45895 3574
rect 9806 3498 9812 3500
rect 8894 3438 9812 3498
rect 7925 3435 7991 3438
rect 8661 3435 8727 3438
rect 9806 3436 9812 3438
rect 9876 3436 9882 3500
rect 9990 3436 9996 3500
rect 10060 3498 10066 3500
rect 12801 3498 12867 3501
rect 29453 3498 29519 3501
rect 30373 3498 30439 3501
rect 10060 3438 12266 3498
rect 10060 3436 10066 3438
rect 2773 3362 2839 3365
rect 4245 3362 4311 3365
rect 5717 3362 5783 3365
rect 5993 3364 6059 3365
rect 2773 3360 4311 3362
rect 2773 3304 2778 3360
rect 2834 3304 4250 3360
rect 4306 3304 4311 3360
rect 2773 3302 4311 3304
rect 2773 3299 2839 3302
rect 4245 3299 4311 3302
rect 5214 3360 5783 3362
rect 5214 3304 5722 3360
rect 5778 3304 5783 3360
rect 5214 3302 5783 3304
rect 2630 3164 2636 3228
rect 2700 3226 2706 3228
rect 2865 3226 2931 3229
rect 4429 3226 4495 3229
rect 2700 3224 2931 3226
rect 2700 3168 2870 3224
rect 2926 3168 2931 3224
rect 2700 3166 2931 3168
rect 2700 3164 2706 3166
rect 2865 3163 2931 3166
rect 3558 3224 4495 3226
rect 3558 3168 4434 3224
rect 4490 3168 4495 3224
rect 3558 3166 4495 3168
rect 3141 3092 3207 3093
rect 3141 3090 3188 3092
rect 3096 3088 3188 3090
rect 3096 3032 3146 3088
rect 3096 3030 3188 3032
rect 3141 3028 3188 3030
rect 3252 3028 3258 3092
rect 3141 3027 3207 3028
rect 1894 2892 1900 2956
rect 1964 2954 1970 2956
rect 2037 2954 2103 2957
rect 1964 2952 2103 2954
rect 1964 2896 2042 2952
rect 2098 2896 2103 2952
rect 1964 2894 2103 2896
rect 1964 2892 1970 2894
rect 2037 2891 2103 2894
rect 2773 2956 2839 2957
rect 2773 2952 2820 2956
rect 2884 2954 2890 2956
rect 3233 2954 3299 2957
rect 3366 2954 3372 2956
rect 2773 2896 2778 2952
rect 2773 2892 2820 2896
rect 2884 2894 2930 2954
rect 3233 2952 3372 2954
rect 3233 2896 3238 2952
rect 3294 2896 3372 2952
rect 3233 2894 3372 2896
rect 2884 2892 2890 2894
rect 2773 2891 2839 2892
rect 3233 2891 3299 2894
rect 3366 2892 3372 2894
rect 3436 2892 3442 2956
rect 0 2818 800 2848
rect 3558 2818 3618 3166
rect 4429 3163 4495 3166
rect 5073 3226 5139 3229
rect 5214 3226 5274 3302
rect 5717 3299 5783 3302
rect 5942 3300 5948 3364
rect 6012 3362 6059 3364
rect 6012 3360 6104 3362
rect 6054 3304 6104 3360
rect 6012 3302 6104 3304
rect 6012 3300 6059 3302
rect 8518 3300 8524 3364
rect 8588 3362 8594 3364
rect 11421 3362 11487 3365
rect 12014 3362 12020 3364
rect 8588 3360 12020 3362
rect 8588 3304 11426 3360
rect 11482 3304 12020 3360
rect 8588 3302 12020 3304
rect 8588 3300 8594 3302
rect 5993 3299 6059 3300
rect 11421 3299 11487 3302
rect 12014 3300 12020 3302
rect 12084 3300 12090 3364
rect 12206 3362 12266 3438
rect 12801 3496 30439 3498
rect 12801 3440 12806 3496
rect 12862 3440 29458 3496
rect 29514 3440 30378 3496
rect 30434 3440 30439 3496
rect 12801 3438 30439 3440
rect 12801 3435 12867 3438
rect 29453 3435 29519 3438
rect 30373 3435 30439 3438
rect 44817 3498 44883 3501
rect 49200 3498 50000 3528
rect 44817 3496 50000 3498
rect 44817 3440 44822 3496
rect 44878 3440 50000 3496
rect 44817 3438 50000 3440
rect 44817 3435 44883 3438
rect 49200 3408 50000 3438
rect 42793 3362 42859 3365
rect 47301 3362 47367 3365
rect 12206 3302 17234 3362
rect 5441 3228 5507 3229
rect 5390 3226 5396 3228
rect 5073 3224 5274 3226
rect 5073 3168 5078 3224
rect 5134 3168 5274 3224
rect 5073 3166 5274 3168
rect 5350 3166 5396 3226
rect 5460 3224 5507 3228
rect 5502 3168 5507 3224
rect 5073 3163 5139 3166
rect 5390 3164 5396 3166
rect 5460 3164 5507 3168
rect 5441 3163 5507 3164
rect 5809 3226 5875 3229
rect 6637 3228 6703 3229
rect 5942 3226 5948 3228
rect 5809 3224 5948 3226
rect 5809 3168 5814 3224
rect 5870 3168 5948 3224
rect 5809 3166 5948 3168
rect 5809 3163 5875 3166
rect 5942 3164 5948 3166
rect 6012 3164 6018 3228
rect 6637 3226 6684 3228
rect 6592 3224 6684 3226
rect 6592 3168 6642 3224
rect 6592 3166 6684 3168
rect 6637 3164 6684 3166
rect 6748 3164 6754 3228
rect 8753 3226 8819 3229
rect 9070 3226 9076 3228
rect 8753 3224 9076 3226
rect 8753 3168 8758 3224
rect 8814 3168 9076 3224
rect 8753 3166 9076 3168
rect 6637 3163 6703 3164
rect 8753 3163 8819 3166
rect 9070 3164 9076 3166
rect 9140 3164 9146 3228
rect 9990 3164 9996 3228
rect 10060 3226 10066 3228
rect 10133 3226 10199 3229
rect 11053 3228 11119 3229
rect 11053 3226 11100 3228
rect 10060 3224 10199 3226
rect 10060 3168 10138 3224
rect 10194 3168 10199 3224
rect 10060 3166 10199 3168
rect 11008 3224 11100 3226
rect 11008 3168 11058 3224
rect 11008 3166 11100 3168
rect 10060 3164 10066 3166
rect 10133 3163 10199 3166
rect 11053 3164 11100 3166
rect 11164 3164 11170 3228
rect 11053 3163 11119 3164
rect 5717 3092 5783 3093
rect 5717 3088 5764 3092
rect 5828 3090 5834 3092
rect 5717 3032 5722 3088
rect 5717 3028 5764 3032
rect 5828 3030 5874 3090
rect 6318 3030 7482 3090
rect 5828 3028 5834 3030
rect 5717 3027 5783 3028
rect 3693 2954 3759 2957
rect 6126 2954 6132 2956
rect 3693 2952 6132 2954
rect 3693 2896 3698 2952
rect 3754 2896 6132 2952
rect 3693 2894 6132 2896
rect 3693 2891 3759 2894
rect 6126 2892 6132 2894
rect 6196 2892 6202 2956
rect 0 2758 3618 2818
rect 5165 2820 5231 2821
rect 5165 2816 5212 2820
rect 5276 2818 5282 2820
rect 5993 2818 6059 2821
rect 6318 2818 6378 3030
rect 7189 2956 7255 2957
rect 7189 2954 7236 2956
rect 7144 2952 7236 2954
rect 7144 2896 7194 2952
rect 7144 2894 7236 2896
rect 7189 2892 7236 2894
rect 7300 2892 7306 2956
rect 7422 2954 7482 3030
rect 8702 3028 8708 3092
rect 8772 3090 8778 3092
rect 9305 3090 9371 3093
rect 8772 3088 9371 3090
rect 8772 3032 9310 3088
rect 9366 3032 9371 3088
rect 8772 3030 9371 3032
rect 8772 3028 8778 3030
rect 9305 3027 9371 3030
rect 9581 3090 9647 3093
rect 12709 3090 12775 3093
rect 9581 3088 12775 3090
rect 9581 3032 9586 3088
rect 9642 3032 12714 3088
rect 12770 3032 12775 3088
rect 9581 3030 12775 3032
rect 17174 3090 17234 3302
rect 42793 3360 47367 3362
rect 42793 3304 42798 3360
rect 42854 3304 47306 3360
rect 47362 3304 47367 3360
rect 42793 3302 47367 3304
rect 42793 3299 42859 3302
rect 47301 3299 47367 3302
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 45093 3226 45159 3229
rect 45645 3226 45711 3229
rect 45093 3224 45711 3226
rect 45093 3168 45098 3224
rect 45154 3168 45650 3224
rect 45706 3168 45711 3224
rect 45093 3166 45711 3168
rect 45093 3163 45159 3166
rect 45645 3163 45711 3166
rect 29821 3090 29887 3093
rect 17174 3088 29887 3090
rect 17174 3032 29826 3088
rect 29882 3032 29887 3088
rect 17174 3030 29887 3032
rect 9581 3027 9647 3030
rect 12709 3027 12775 3030
rect 29821 3027 29887 3030
rect 10174 2954 10180 2956
rect 7422 2894 10180 2954
rect 10174 2892 10180 2894
rect 10244 2892 10250 2956
rect 11237 2954 11303 2957
rect 10366 2952 11303 2954
rect 10366 2896 11242 2952
rect 11298 2896 11303 2952
rect 10366 2894 11303 2896
rect 7189 2891 7255 2892
rect 5165 2760 5170 2816
rect 0 2728 800 2758
rect 5165 2756 5212 2760
rect 5276 2758 5322 2818
rect 5993 2816 6378 2818
rect 5993 2760 5998 2816
rect 6054 2760 6378 2816
rect 5993 2758 6378 2760
rect 7833 2818 7899 2821
rect 8150 2818 8156 2820
rect 7833 2816 8156 2818
rect 7833 2760 7838 2816
rect 7894 2760 8156 2816
rect 7833 2758 8156 2760
rect 5276 2756 5282 2758
rect 5165 2755 5231 2756
rect 5993 2755 6059 2758
rect 7833 2755 7899 2758
rect 8150 2756 8156 2758
rect 8220 2756 8226 2820
rect 9438 2818 9444 2820
rect 8342 2758 9444 2818
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 8342 2685 8402 2758
rect 9438 2756 9444 2758
rect 9508 2756 9514 2820
rect 9673 2818 9739 2821
rect 10366 2818 10426 2894
rect 11237 2891 11303 2894
rect 45553 2954 45619 2957
rect 49200 2954 50000 2984
rect 45553 2952 50000 2954
rect 45553 2896 45558 2952
rect 45614 2896 50000 2952
rect 45553 2894 50000 2896
rect 45553 2891 45619 2894
rect 49200 2864 50000 2894
rect 9673 2816 10426 2818
rect 9673 2760 9678 2816
rect 9734 2760 10426 2816
rect 9673 2758 10426 2760
rect 10777 2818 10843 2821
rect 11329 2818 11395 2821
rect 10777 2816 11395 2818
rect 10777 2760 10782 2816
rect 10838 2760 11334 2816
rect 11390 2760 11395 2816
rect 10777 2758 11395 2760
rect 9673 2755 9739 2758
rect 10777 2755 10843 2758
rect 11329 2755 11395 2758
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 1894 2620 1900 2684
rect 1964 2682 1970 2684
rect 2221 2682 2287 2685
rect 3509 2682 3575 2685
rect 1964 2680 2287 2682
rect 1964 2624 2226 2680
rect 2282 2624 2287 2680
rect 1964 2622 2287 2624
rect 1964 2620 1970 2622
rect 2221 2619 2287 2622
rect 3374 2680 3575 2682
rect 3374 2624 3514 2680
rect 3570 2624 3575 2680
rect 3374 2622 3575 2624
rect 3049 2412 3115 2413
rect 2998 2410 3004 2412
rect 2958 2350 3004 2410
rect 3068 2408 3115 2412
rect 3110 2352 3115 2408
rect 2998 2348 3004 2350
rect 3068 2348 3115 2352
rect 3049 2347 3115 2348
rect 3233 2274 3299 2277
rect 3374 2274 3434 2622
rect 3509 2619 3575 2622
rect 5574 2620 5580 2684
rect 5644 2682 5650 2684
rect 7097 2682 7163 2685
rect 5644 2680 7163 2682
rect 5644 2624 7102 2680
rect 7158 2624 7163 2680
rect 5644 2622 7163 2624
rect 5644 2620 5650 2622
rect 7097 2619 7163 2622
rect 8293 2680 8402 2685
rect 8293 2624 8298 2680
rect 8354 2624 8402 2680
rect 8293 2622 8402 2624
rect 8569 2682 8635 2685
rect 8886 2682 8892 2684
rect 8569 2680 8892 2682
rect 8569 2624 8574 2680
rect 8630 2624 8892 2680
rect 8569 2622 8892 2624
rect 8293 2619 8359 2622
rect 8569 2619 8635 2622
rect 8886 2620 8892 2622
rect 8956 2620 8962 2684
rect 9029 2682 9095 2685
rect 10225 2682 10291 2685
rect 9029 2680 10291 2682
rect 9029 2624 9034 2680
rect 9090 2624 10230 2680
rect 10286 2624 10291 2680
rect 9029 2622 10291 2624
rect 9029 2619 9095 2622
rect 10225 2619 10291 2622
rect 11789 2682 11855 2685
rect 17769 2682 17835 2685
rect 11789 2680 17835 2682
rect 11789 2624 11794 2680
rect 11850 2624 17774 2680
rect 17830 2624 17835 2680
rect 11789 2622 17835 2624
rect 11789 2619 11855 2622
rect 17769 2619 17835 2622
rect 3509 2546 3575 2549
rect 3734 2546 3740 2548
rect 3509 2544 3740 2546
rect 3509 2488 3514 2544
rect 3570 2488 3740 2544
rect 3509 2486 3740 2488
rect 3509 2483 3575 2486
rect 3734 2484 3740 2486
rect 3804 2484 3810 2548
rect 4245 2546 4311 2549
rect 4654 2546 4660 2548
rect 4245 2544 4660 2546
rect 4245 2488 4250 2544
rect 4306 2488 4660 2544
rect 4245 2486 4660 2488
rect 4245 2483 4311 2486
rect 4654 2484 4660 2486
rect 4724 2484 4730 2548
rect 5809 2546 5875 2549
rect 7230 2546 7236 2548
rect 5809 2544 7236 2546
rect 5809 2488 5814 2544
rect 5870 2488 7236 2544
rect 5809 2486 7236 2488
rect 5809 2483 5875 2486
rect 7230 2484 7236 2486
rect 7300 2484 7306 2548
rect 7925 2546 7991 2549
rect 8518 2546 8524 2548
rect 7925 2544 8524 2546
rect 7925 2488 7930 2544
rect 7986 2488 8524 2544
rect 7925 2486 8524 2488
rect 7925 2483 7991 2486
rect 8518 2484 8524 2486
rect 8588 2484 8594 2548
rect 9673 2546 9739 2549
rect 9990 2546 9996 2548
rect 9673 2544 9996 2546
rect 9673 2488 9678 2544
rect 9734 2488 9996 2544
rect 9673 2486 9996 2488
rect 9673 2483 9739 2486
rect 9990 2484 9996 2486
rect 10060 2546 10066 2548
rect 12893 2546 12959 2549
rect 10060 2544 12959 2546
rect 10060 2488 12898 2544
rect 12954 2488 12959 2544
rect 10060 2486 12959 2488
rect 10060 2484 10066 2486
rect 12893 2483 12959 2486
rect 3785 2410 3851 2413
rect 6821 2412 6887 2413
rect 7005 2412 7071 2413
rect 3918 2410 3924 2412
rect 3785 2408 3924 2410
rect 3785 2352 3790 2408
rect 3846 2352 3924 2408
rect 3785 2350 3924 2352
rect 3785 2347 3851 2350
rect 3918 2348 3924 2350
rect 3988 2348 3994 2412
rect 6821 2410 6868 2412
rect 6776 2408 6868 2410
rect 6776 2352 6826 2408
rect 6776 2350 6868 2352
rect 6821 2348 6868 2350
rect 6932 2348 6938 2412
rect 7005 2408 7052 2412
rect 7116 2410 7122 2412
rect 8477 2410 8543 2413
rect 9254 2410 9260 2412
rect 7005 2352 7010 2408
rect 7005 2348 7052 2352
rect 7116 2350 7162 2410
rect 8477 2408 9260 2410
rect 8477 2352 8482 2408
rect 8538 2352 9260 2408
rect 8477 2350 9260 2352
rect 7116 2348 7122 2350
rect 6821 2347 6887 2348
rect 7005 2347 7071 2348
rect 8477 2347 8543 2350
rect 9254 2348 9260 2350
rect 9324 2348 9330 2412
rect 9949 2410 10015 2413
rect 11462 2410 11468 2412
rect 9949 2408 11468 2410
rect 9949 2352 9954 2408
rect 10010 2352 11468 2408
rect 9949 2350 11468 2352
rect 9949 2347 10015 2350
rect 11462 2348 11468 2350
rect 11532 2348 11538 2412
rect 11973 2410 12039 2413
rect 13169 2410 13235 2413
rect 11973 2408 13235 2410
rect 11973 2352 11978 2408
rect 12034 2352 13174 2408
rect 13230 2352 13235 2408
rect 11973 2350 13235 2352
rect 11973 2347 12039 2350
rect 13169 2347 13235 2350
rect 3233 2272 3434 2274
rect 3233 2216 3238 2272
rect 3294 2216 3434 2272
rect 3233 2214 3434 2216
rect 6361 2274 6427 2277
rect 7414 2274 7420 2276
rect 6361 2272 7420 2274
rect 6361 2216 6366 2272
rect 6422 2216 7420 2272
rect 6361 2214 7420 2216
rect 3233 2211 3299 2214
rect 6361 2211 6427 2214
rect 7414 2212 7420 2214
rect 7484 2212 7490 2276
rect 10174 2212 10180 2276
rect 10244 2274 10250 2276
rect 10869 2274 10935 2277
rect 10244 2272 10935 2274
rect 10244 2216 10874 2272
rect 10930 2216 10935 2272
rect 10244 2214 10935 2216
rect 10244 2212 10250 2214
rect 10869 2211 10935 2214
rect 46841 2274 46907 2277
rect 49200 2274 50000 2304
rect 46841 2272 50000 2274
rect 46841 2216 46846 2272
rect 46902 2216 50000 2272
rect 46841 2214 50000 2216
rect 46841 2211 46907 2214
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 49200 2184 50000 2214
rect 19568 2143 19888 2144
rect 1158 2076 1164 2140
rect 1228 2138 1234 2140
rect 10317 2138 10383 2141
rect 1228 2136 10383 2138
rect 1228 2080 10322 2136
rect 10378 2080 10383 2136
rect 1228 2078 10383 2080
rect 1228 2076 1234 2078
rect 10317 2075 10383 2078
rect 2865 2002 2931 2005
rect 3550 2002 3556 2004
rect 2865 2000 3556 2002
rect 2865 1944 2870 2000
rect 2926 1944 3556 2000
rect 2865 1942 3556 1944
rect 2865 1939 2931 1942
rect 3550 1940 3556 1942
rect 3620 1940 3626 2004
rect 6637 2002 6703 2005
rect 7598 2002 7604 2004
rect 6637 2000 7604 2002
rect 6637 1944 6642 2000
rect 6698 1944 7604 2000
rect 6637 1942 7604 1944
rect 6637 1939 6703 1942
rect 7598 1940 7604 1942
rect 7668 1940 7674 2004
rect 8937 2002 9003 2005
rect 10910 2002 10916 2004
rect 8937 2000 10916 2002
rect 8937 1944 8942 2000
rect 8998 1944 10916 2000
rect 8937 1942 10916 1944
rect 8937 1939 9003 1942
rect 10910 1940 10916 1942
rect 10980 1940 10986 2004
rect 2078 1804 2084 1868
rect 2148 1866 2154 1868
rect 3693 1866 3759 1869
rect 2148 1864 3759 1866
rect 2148 1808 3698 1864
rect 3754 1808 3759 1864
rect 2148 1806 3759 1808
rect 2148 1804 2154 1806
rect 3693 1803 3759 1806
rect 7281 1730 7347 1733
rect 7238 1728 7347 1730
rect 7238 1672 7286 1728
rect 7342 1672 7347 1728
rect 7238 1667 7347 1672
rect 7097 1594 7163 1597
rect 7238 1594 7298 1667
rect 7097 1592 7298 1594
rect 7097 1536 7102 1592
rect 7158 1536 7298 1592
rect 7097 1534 7298 1536
rect 46749 1594 46815 1597
rect 49200 1594 50000 1624
rect 46749 1592 50000 1594
rect 46749 1536 46754 1592
rect 46810 1536 50000 1592
rect 46749 1534 50000 1536
rect 7097 1531 7163 1534
rect 46749 1531 46815 1534
rect 49200 1504 50000 1534
rect 3969 1322 4035 1325
rect 5758 1322 5764 1324
rect 3969 1320 5764 1322
rect 3969 1264 3974 1320
rect 4030 1264 5764 1320
rect 3969 1262 5764 1264
rect 3969 1259 4035 1262
rect 5758 1260 5764 1262
rect 5828 1260 5834 1324
rect 8334 1260 8340 1324
rect 8404 1322 8410 1324
rect 9029 1322 9095 1325
rect 8404 1320 9095 1322
rect 8404 1264 9034 1320
rect 9090 1264 9095 1320
rect 8404 1262 9095 1264
rect 8404 1260 8410 1262
rect 9029 1259 9095 1262
rect 5165 1186 5231 1189
rect 6494 1186 6500 1188
rect 5165 1184 6500 1186
rect 5165 1128 5170 1184
rect 5226 1128 6500 1184
rect 5165 1126 6500 1128
rect 5165 1123 5231 1126
rect 6494 1124 6500 1126
rect 6564 1124 6570 1188
rect 4797 1050 4863 1053
rect 6310 1050 6316 1052
rect 4797 1048 6316 1050
rect 4797 992 4802 1048
rect 4858 992 6316 1048
rect 4797 990 6316 992
rect 4797 987 4863 990
rect 6310 988 6316 990
rect 6380 988 6386 1052
rect 5625 914 5691 917
rect 7782 914 7788 916
rect 5625 912 7788 914
rect 5625 856 5630 912
rect 5686 856 7788 912
rect 5625 854 7788 856
rect 5625 851 5691 854
rect 7782 852 7788 854
rect 7852 852 7858 916
rect 42609 914 42675 917
rect 49200 914 50000 944
rect 42609 912 50000 914
rect 42609 856 42614 912
rect 42670 856 50000 912
rect 42609 854 50000 856
rect 42609 851 42675 854
rect 49200 824 50000 854
rect 46473 370 46539 373
rect 49200 370 50000 400
rect 46473 368 50000 370
rect 46473 312 46478 368
rect 46534 312 50000 368
rect 46473 310 50000 312
rect 46473 307 46539 310
rect 49200 280 50000 310
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 7972 42468 8036 42532
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 48084 26420 48148 26484
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 47164 21312 47228 21316
rect 47164 21256 47214 21312
rect 47214 21256 47228 21312
rect 47164 21252 47228 21256
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 47716 20708 47780 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 46060 17988 46124 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 47164 17036 47228 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 47716 16144 47780 16148
rect 47716 16088 47766 16144
rect 47766 16088 47780 16144
rect 47716 16084 47780 16088
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 46060 12472 46124 12476
rect 46060 12416 46074 12472
rect 46074 12416 46124 12472
rect 46060 12412 46124 12416
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 1164 11052 1228 11116
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 3740 9420 3804 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4844 8876 4908 8940
rect 3556 8740 3620 8804
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 3924 8604 3988 8668
rect 2268 8392 2332 8396
rect 2268 8336 2318 8392
rect 2318 8336 2332 8392
rect 2268 8332 2332 8336
rect 4660 8392 4724 8396
rect 4660 8336 4710 8392
rect 4710 8336 4724 8392
rect 4660 8332 4724 8336
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 2084 7788 2148 7852
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 2820 7304 2884 7308
rect 2820 7248 2834 7304
rect 2834 7248 2884 7304
rect 2820 7244 2884 7248
rect 3372 7244 3436 7308
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 2452 7032 2516 7036
rect 2452 6976 2466 7032
rect 2466 6976 2516 7032
rect 2452 6972 2516 6976
rect 3004 7032 3068 7036
rect 3004 6976 3054 7032
rect 3054 6976 3068 7032
rect 3004 6972 3068 6976
rect 3188 6972 3252 7036
rect 5212 7244 5276 7308
rect 5396 7244 5460 7308
rect 7604 7244 7668 7308
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 8340 6972 8404 7036
rect 2636 6700 2700 6764
rect 5580 6760 5644 6764
rect 5580 6704 5594 6760
rect 5594 6704 5644 6760
rect 5580 6700 5644 6704
rect 7420 6700 7484 6764
rect 9812 6700 9876 6764
rect 11468 6700 11532 6764
rect 5028 6564 5092 6628
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 5948 6428 6012 6492
rect 10180 6428 10244 6492
rect 48084 6428 48148 6492
rect 11100 6292 11164 6356
rect 5212 6020 5276 6084
rect 6868 6020 6932 6084
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 7236 5884 7300 5948
rect 5212 5748 5276 5812
rect 9996 5748 10060 5812
rect 3740 5476 3804 5540
rect 6500 5476 6564 5540
rect 5580 5340 5644 5404
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 3556 4524 3620 4588
rect 3740 4388 3804 4452
rect 5212 5204 5276 5268
rect 7052 5204 7116 5268
rect 7788 5340 7852 5404
rect 8524 5340 8588 5404
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 5212 5068 5276 5132
rect 6684 5128 6748 5132
rect 6684 5072 6734 5128
rect 6734 5072 6748 5128
rect 6684 5068 6748 5072
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 8156 4796 8220 4860
rect 9260 4796 9324 4860
rect 9076 4660 9140 4724
rect 11100 4660 11164 4724
rect 8708 4524 8772 4588
rect 8892 4388 8956 4452
rect 10916 4448 10980 4452
rect 10916 4392 10966 4448
rect 10966 4392 10980 4448
rect 10916 4388 10980 4392
rect 11100 4388 11164 4452
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 5764 4252 5828 4316
rect 9444 4252 9508 4316
rect 2268 4176 2332 4180
rect 2268 4120 2318 4176
rect 2318 4120 2332 4176
rect 2268 4116 2332 4120
rect 2452 3980 2516 4044
rect 3004 4040 3068 4044
rect 3004 3984 3054 4040
rect 3054 3984 3068 4040
rect 3004 3980 3068 3984
rect 3004 3844 3068 3908
rect 5580 4116 5644 4180
rect 6316 4116 6380 4180
rect 8340 4116 8404 4180
rect 4660 4040 4724 4044
rect 4660 3984 4710 4040
rect 4710 3984 4724 4040
rect 4660 3980 4724 3984
rect 7236 3980 7300 4044
rect 7972 4040 8036 4044
rect 7972 3984 7986 4040
rect 7986 3984 8036 4040
rect 7972 3980 8036 3984
rect 3924 3844 3988 3908
rect 4660 3904 4724 3908
rect 4660 3848 4674 3904
rect 4674 3848 4724 3904
rect 4660 3844 4724 3848
rect 6132 3844 6196 3908
rect 10180 3980 10244 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 8524 3708 8588 3772
rect 12020 3844 12084 3908
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 5028 3572 5092 3636
rect 8340 3572 8404 3636
rect 4844 3436 4908 3500
rect 9812 3436 9876 3500
rect 9996 3436 10060 3500
rect 2636 3164 2700 3228
rect 3188 3088 3252 3092
rect 3188 3032 3202 3088
rect 3202 3032 3252 3088
rect 3188 3028 3252 3032
rect 1900 2892 1964 2956
rect 2820 2952 2884 2956
rect 2820 2896 2834 2952
rect 2834 2896 2884 2952
rect 2820 2892 2884 2896
rect 3372 2892 3436 2956
rect 5948 3360 6012 3364
rect 5948 3304 5998 3360
rect 5998 3304 6012 3360
rect 5948 3300 6012 3304
rect 8524 3300 8588 3364
rect 12020 3300 12084 3364
rect 5396 3224 5460 3228
rect 5396 3168 5446 3224
rect 5446 3168 5460 3224
rect 5396 3164 5460 3168
rect 5948 3164 6012 3228
rect 6684 3224 6748 3228
rect 6684 3168 6698 3224
rect 6698 3168 6748 3224
rect 6684 3164 6748 3168
rect 9076 3164 9140 3228
rect 9996 3164 10060 3228
rect 11100 3224 11164 3228
rect 11100 3168 11114 3224
rect 11114 3168 11164 3224
rect 11100 3164 11164 3168
rect 5764 3088 5828 3092
rect 5764 3032 5778 3088
rect 5778 3032 5828 3088
rect 5764 3028 5828 3032
rect 6132 2892 6196 2956
rect 5212 2816 5276 2820
rect 7236 2952 7300 2956
rect 7236 2896 7250 2952
rect 7250 2896 7300 2952
rect 7236 2892 7300 2896
rect 8708 3028 8772 3092
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 10180 2892 10244 2956
rect 5212 2760 5226 2816
rect 5226 2760 5276 2816
rect 5212 2756 5276 2760
rect 8156 2756 8220 2820
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 9444 2756 9508 2820
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 1900 2620 1964 2684
rect 3004 2408 3068 2412
rect 3004 2352 3054 2408
rect 3054 2352 3068 2408
rect 3004 2348 3068 2352
rect 5580 2620 5644 2684
rect 8892 2620 8956 2684
rect 3740 2484 3804 2548
rect 4660 2484 4724 2548
rect 7236 2484 7300 2548
rect 8524 2484 8588 2548
rect 9996 2484 10060 2548
rect 3924 2348 3988 2412
rect 6868 2408 6932 2412
rect 6868 2352 6882 2408
rect 6882 2352 6932 2408
rect 6868 2348 6932 2352
rect 7052 2408 7116 2412
rect 7052 2352 7066 2408
rect 7066 2352 7116 2408
rect 7052 2348 7116 2352
rect 9260 2348 9324 2412
rect 11468 2348 11532 2412
rect 7420 2212 7484 2276
rect 10180 2212 10244 2276
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 1164 2076 1228 2140
rect 3556 1940 3620 2004
rect 7604 1940 7668 2004
rect 10916 1940 10980 2004
rect 2084 1804 2148 1868
rect 5764 1260 5828 1324
rect 8340 1260 8404 1324
rect 6500 1124 6564 1188
rect 6316 988 6380 1052
rect 7788 852 7852 916
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 7971 42532 8037 42533
rect 7971 42468 7972 42532
rect 8036 42468 8037 42532
rect 7971 42467 8037 42468
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 1163 11116 1229 11117
rect 1163 11052 1164 11116
rect 1228 11052 1229 11116
rect 1163 11051 1229 11052
rect 1166 2141 1226 11051
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 3739 9484 3805 9485
rect 3739 9420 3740 9484
rect 3804 9420 3805 9484
rect 3739 9419 3805 9420
rect 3555 8804 3621 8805
rect 3555 8740 3556 8804
rect 3620 8740 3621 8804
rect 3555 8739 3621 8740
rect 2267 8396 2333 8397
rect 2267 8332 2268 8396
rect 2332 8332 2333 8396
rect 2267 8331 2333 8332
rect 2083 7852 2149 7853
rect 2083 7788 2084 7852
rect 2148 7788 2149 7852
rect 2083 7787 2149 7788
rect 1899 2956 1965 2957
rect 1899 2892 1900 2956
rect 1964 2892 1965 2956
rect 1899 2891 1965 2892
rect 1902 2685 1962 2891
rect 1899 2684 1965 2685
rect 1899 2620 1900 2684
rect 1964 2620 1965 2684
rect 1899 2619 1965 2620
rect 1163 2140 1229 2141
rect 1163 2076 1164 2140
rect 1228 2076 1229 2140
rect 1163 2075 1229 2076
rect 2086 1869 2146 7787
rect 2270 4181 2330 8331
rect 2819 7308 2885 7309
rect 2819 7244 2820 7308
rect 2884 7244 2885 7308
rect 2819 7243 2885 7244
rect 3371 7308 3437 7309
rect 3371 7244 3372 7308
rect 3436 7244 3437 7308
rect 3371 7243 3437 7244
rect 2451 7036 2517 7037
rect 2451 6972 2452 7036
rect 2516 6972 2517 7036
rect 2451 6971 2517 6972
rect 2267 4180 2333 4181
rect 2267 4116 2268 4180
rect 2332 4116 2333 4180
rect 2267 4115 2333 4116
rect 2454 4045 2514 6971
rect 2635 6764 2701 6765
rect 2635 6700 2636 6764
rect 2700 6700 2701 6764
rect 2635 6699 2701 6700
rect 2451 4044 2517 4045
rect 2451 3980 2452 4044
rect 2516 3980 2517 4044
rect 2451 3979 2517 3980
rect 2638 3229 2698 6699
rect 2635 3228 2701 3229
rect 2635 3164 2636 3228
rect 2700 3164 2701 3228
rect 2635 3163 2701 3164
rect 2822 2957 2882 7243
rect 3003 7036 3069 7037
rect 3003 6972 3004 7036
rect 3068 6972 3069 7036
rect 3003 6971 3069 6972
rect 3187 7036 3253 7037
rect 3187 6972 3188 7036
rect 3252 6972 3253 7036
rect 3187 6971 3253 6972
rect 3006 4045 3066 6971
rect 3003 4044 3069 4045
rect 3003 3980 3004 4044
rect 3068 3980 3069 4044
rect 3003 3979 3069 3980
rect 3003 3908 3069 3909
rect 3003 3844 3004 3908
rect 3068 3844 3069 3908
rect 3003 3843 3069 3844
rect 2819 2956 2885 2957
rect 2819 2892 2820 2956
rect 2884 2892 2885 2956
rect 2819 2891 2885 2892
rect 3006 2413 3066 3843
rect 3190 3093 3250 6971
rect 3187 3092 3253 3093
rect 3187 3028 3188 3092
rect 3252 3028 3253 3092
rect 3187 3027 3253 3028
rect 3374 2957 3434 7243
rect 3558 4589 3618 8739
rect 3742 5541 3802 9419
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 3923 8668 3989 8669
rect 3923 8604 3924 8668
rect 3988 8604 3989 8668
rect 3923 8603 3989 8604
rect 3739 5540 3805 5541
rect 3739 5476 3740 5540
rect 3804 5476 3805 5540
rect 3739 5475 3805 5476
rect 3555 4588 3621 4589
rect 3555 4524 3556 4588
rect 3620 4524 3621 4588
rect 3555 4523 3621 4524
rect 3371 2956 3437 2957
rect 3371 2892 3372 2956
rect 3436 2892 3437 2956
rect 3371 2891 3437 2892
rect 3003 2412 3069 2413
rect 3003 2348 3004 2412
rect 3068 2348 3069 2412
rect 3003 2347 3069 2348
rect 3558 2005 3618 4523
rect 3739 4452 3805 4453
rect 3739 4388 3740 4452
rect 3804 4450 3805 4452
rect 3926 4450 3986 8603
rect 3804 4390 3986 4450
rect 4208 8192 4528 9216
rect 4843 8940 4909 8941
rect 4843 8876 4844 8940
rect 4908 8876 4909 8940
rect 4843 8875 4909 8876
rect 4659 8396 4725 8397
rect 4659 8332 4660 8396
rect 4724 8332 4725 8396
rect 4659 8331 4725 8332
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 3804 4388 3805 4390
rect 3739 4387 3805 4388
rect 3742 2549 3802 4387
rect 3923 3908 3989 3909
rect 3923 3844 3924 3908
rect 3988 3844 3989 3908
rect 3923 3843 3989 3844
rect 3739 2548 3805 2549
rect 3739 2484 3740 2548
rect 3804 2484 3805 2548
rect 3739 2483 3805 2484
rect 3926 2413 3986 3843
rect 4208 3840 4528 4864
rect 4662 4045 4722 8331
rect 4659 4044 4725 4045
rect 4659 3980 4660 4044
rect 4724 3980 4725 4044
rect 4659 3979 4725 3980
rect 4659 3908 4725 3909
rect 4659 3844 4660 3908
rect 4724 3844 4725 3908
rect 4659 3843 4725 3844
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 3923 2412 3989 2413
rect 3923 2348 3924 2412
rect 3988 2348 3989 2412
rect 3923 2347 3989 2348
rect 4208 2128 4528 2688
rect 4662 2549 4722 3843
rect 4846 3501 4906 8875
rect 5211 7308 5277 7309
rect 5211 7244 5212 7308
rect 5276 7244 5277 7308
rect 5211 7243 5277 7244
rect 5395 7308 5461 7309
rect 5395 7244 5396 7308
rect 5460 7244 5461 7308
rect 5395 7243 5461 7244
rect 7603 7308 7669 7309
rect 7603 7244 7604 7308
rect 7668 7244 7669 7308
rect 7603 7243 7669 7244
rect 5027 6628 5093 6629
rect 5027 6564 5028 6628
rect 5092 6564 5093 6628
rect 5027 6563 5093 6564
rect 5030 3637 5090 6563
rect 5214 6085 5274 7243
rect 5211 6084 5277 6085
rect 5211 6020 5212 6084
rect 5276 6020 5277 6084
rect 5211 6019 5277 6020
rect 5211 5812 5277 5813
rect 5211 5748 5212 5812
rect 5276 5748 5277 5812
rect 5211 5747 5277 5748
rect 5214 5269 5274 5747
rect 5211 5268 5277 5269
rect 5211 5204 5212 5268
rect 5276 5204 5277 5268
rect 5211 5203 5277 5204
rect 5211 5132 5277 5133
rect 5211 5068 5212 5132
rect 5276 5068 5277 5132
rect 5211 5067 5277 5068
rect 5027 3636 5093 3637
rect 5027 3572 5028 3636
rect 5092 3572 5093 3636
rect 5027 3571 5093 3572
rect 4843 3500 4909 3501
rect 4843 3436 4844 3500
rect 4908 3436 4909 3500
rect 4843 3435 4909 3436
rect 5214 2821 5274 5067
rect 5398 3229 5458 7243
rect 5579 6764 5645 6765
rect 5579 6700 5580 6764
rect 5644 6700 5645 6764
rect 5579 6699 5645 6700
rect 7419 6764 7485 6765
rect 7419 6700 7420 6764
rect 7484 6700 7485 6764
rect 7419 6699 7485 6700
rect 5582 5405 5642 6699
rect 5947 6492 6013 6493
rect 5947 6428 5948 6492
rect 6012 6428 6013 6492
rect 5947 6427 6013 6428
rect 5579 5404 5645 5405
rect 5579 5340 5580 5404
rect 5644 5340 5645 5404
rect 5579 5339 5645 5340
rect 5763 4316 5829 4317
rect 5763 4252 5764 4316
rect 5828 4252 5829 4316
rect 5763 4251 5829 4252
rect 5579 4180 5645 4181
rect 5579 4116 5580 4180
rect 5644 4116 5645 4180
rect 5579 4115 5645 4116
rect 5395 3228 5461 3229
rect 5395 3164 5396 3228
rect 5460 3164 5461 3228
rect 5395 3163 5461 3164
rect 5211 2820 5277 2821
rect 5211 2756 5212 2820
rect 5276 2756 5277 2820
rect 5211 2755 5277 2756
rect 5582 2685 5642 4115
rect 5766 3093 5826 4251
rect 5950 3365 6010 6427
rect 6867 6084 6933 6085
rect 6867 6020 6868 6084
rect 6932 6020 6933 6084
rect 6867 6019 6933 6020
rect 6499 5540 6565 5541
rect 6499 5476 6500 5540
rect 6564 5476 6565 5540
rect 6499 5475 6565 5476
rect 6315 4180 6381 4181
rect 6315 4116 6316 4180
rect 6380 4116 6381 4180
rect 6315 4115 6381 4116
rect 6131 3908 6197 3909
rect 6131 3844 6132 3908
rect 6196 3844 6197 3908
rect 6131 3843 6197 3844
rect 5947 3364 6013 3365
rect 5947 3300 5948 3364
rect 6012 3300 6013 3364
rect 5947 3299 6013 3300
rect 5947 3228 6013 3229
rect 5947 3164 5948 3228
rect 6012 3164 6013 3228
rect 5947 3163 6013 3164
rect 5763 3092 5829 3093
rect 5763 3028 5764 3092
rect 5828 3028 5829 3092
rect 5763 3027 5829 3028
rect 5950 2790 6010 3163
rect 6134 2957 6194 3843
rect 6131 2956 6197 2957
rect 6131 2892 6132 2956
rect 6196 2892 6197 2956
rect 6131 2891 6197 2892
rect 5766 2730 6010 2790
rect 5579 2684 5645 2685
rect 5579 2620 5580 2684
rect 5644 2620 5645 2684
rect 5579 2619 5645 2620
rect 4659 2548 4725 2549
rect 4659 2484 4660 2548
rect 4724 2484 4725 2548
rect 4659 2483 4725 2484
rect 3555 2004 3621 2005
rect 3555 1940 3556 2004
rect 3620 1940 3621 2004
rect 3555 1939 3621 1940
rect 2083 1868 2149 1869
rect 2083 1804 2084 1868
rect 2148 1804 2149 1868
rect 2083 1803 2149 1804
rect 5766 1325 5826 2730
rect 5763 1324 5829 1325
rect 5763 1260 5764 1324
rect 5828 1260 5829 1324
rect 5763 1259 5829 1260
rect 6318 1053 6378 4115
rect 6502 1189 6562 5475
rect 6683 5132 6749 5133
rect 6683 5068 6684 5132
rect 6748 5068 6749 5132
rect 6683 5067 6749 5068
rect 6686 3229 6746 5067
rect 6683 3228 6749 3229
rect 6683 3164 6684 3228
rect 6748 3164 6749 3228
rect 6683 3163 6749 3164
rect 6870 2413 6930 6019
rect 7235 5948 7301 5949
rect 7235 5884 7236 5948
rect 7300 5884 7301 5948
rect 7235 5883 7301 5884
rect 7051 5268 7117 5269
rect 7051 5204 7052 5268
rect 7116 5204 7117 5268
rect 7051 5203 7117 5204
rect 7054 2413 7114 5203
rect 7238 4045 7298 5883
rect 7235 4044 7301 4045
rect 7235 3980 7236 4044
rect 7300 3980 7301 4044
rect 7235 3979 7301 3980
rect 7235 2956 7301 2957
rect 7235 2892 7236 2956
rect 7300 2892 7301 2956
rect 7235 2891 7301 2892
rect 7238 2549 7298 2891
rect 7235 2548 7301 2549
rect 7235 2484 7236 2548
rect 7300 2484 7301 2548
rect 7235 2483 7301 2484
rect 6867 2412 6933 2413
rect 6867 2348 6868 2412
rect 6932 2348 6933 2412
rect 6867 2347 6933 2348
rect 7051 2412 7117 2413
rect 7051 2348 7052 2412
rect 7116 2348 7117 2412
rect 7051 2347 7117 2348
rect 7422 2277 7482 6699
rect 7419 2276 7485 2277
rect 7419 2212 7420 2276
rect 7484 2212 7485 2276
rect 7419 2211 7485 2212
rect 7606 2005 7666 7243
rect 7787 5404 7853 5405
rect 7787 5340 7788 5404
rect 7852 5340 7853 5404
rect 7787 5339 7853 5340
rect 7603 2004 7669 2005
rect 7603 1940 7604 2004
rect 7668 1940 7669 2004
rect 7603 1939 7669 1940
rect 6499 1188 6565 1189
rect 6499 1124 6500 1188
rect 6564 1124 6565 1188
rect 6499 1123 6565 1124
rect 6315 1052 6381 1053
rect 6315 988 6316 1052
rect 6380 988 6381 1052
rect 6315 987 6381 988
rect 7790 917 7850 5339
rect 7974 4045 8034 42467
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 8339 7036 8405 7037
rect 8339 6972 8340 7036
rect 8404 6972 8405 7036
rect 8339 6971 8405 6972
rect 8155 4860 8221 4861
rect 8155 4796 8156 4860
rect 8220 4796 8221 4860
rect 8155 4795 8221 4796
rect 7971 4044 8037 4045
rect 7971 3980 7972 4044
rect 8036 3980 8037 4044
rect 7971 3979 8037 3980
rect 8158 2821 8218 4795
rect 8342 4181 8402 6971
rect 9811 6764 9877 6765
rect 9811 6700 9812 6764
rect 9876 6700 9877 6764
rect 9811 6699 9877 6700
rect 11467 6764 11533 6765
rect 11467 6700 11468 6764
rect 11532 6700 11533 6764
rect 11467 6699 11533 6700
rect 8523 5404 8589 5405
rect 8523 5340 8524 5404
rect 8588 5340 8589 5404
rect 8523 5339 8589 5340
rect 8339 4180 8405 4181
rect 8339 4116 8340 4180
rect 8404 4116 8405 4180
rect 8339 4115 8405 4116
rect 8526 3773 8586 5339
rect 9259 4860 9325 4861
rect 9259 4796 9260 4860
rect 9324 4796 9325 4860
rect 9259 4795 9325 4796
rect 9075 4724 9141 4725
rect 9075 4660 9076 4724
rect 9140 4660 9141 4724
rect 9075 4659 9141 4660
rect 8707 4588 8773 4589
rect 8707 4524 8708 4588
rect 8772 4524 8773 4588
rect 8707 4523 8773 4524
rect 8523 3772 8589 3773
rect 8523 3708 8524 3772
rect 8588 3708 8589 3772
rect 8523 3707 8589 3708
rect 8339 3636 8405 3637
rect 8339 3572 8340 3636
rect 8404 3572 8405 3636
rect 8339 3571 8405 3572
rect 8155 2820 8221 2821
rect 8155 2756 8156 2820
rect 8220 2756 8221 2820
rect 8155 2755 8221 2756
rect 8342 1325 8402 3571
rect 8523 3364 8589 3365
rect 8523 3300 8524 3364
rect 8588 3300 8589 3364
rect 8523 3299 8589 3300
rect 8526 2549 8586 3299
rect 8710 3093 8770 4523
rect 8891 4452 8957 4453
rect 8891 4388 8892 4452
rect 8956 4388 8957 4452
rect 8891 4387 8957 4388
rect 8707 3092 8773 3093
rect 8707 3028 8708 3092
rect 8772 3028 8773 3092
rect 8707 3027 8773 3028
rect 8894 2685 8954 4387
rect 9078 3229 9138 4659
rect 9075 3228 9141 3229
rect 9075 3164 9076 3228
rect 9140 3164 9141 3228
rect 9075 3163 9141 3164
rect 8891 2684 8957 2685
rect 8891 2620 8892 2684
rect 8956 2620 8957 2684
rect 8891 2619 8957 2620
rect 8523 2548 8589 2549
rect 8523 2484 8524 2548
rect 8588 2484 8589 2548
rect 8523 2483 8589 2484
rect 9262 2413 9322 4795
rect 9443 4316 9509 4317
rect 9443 4252 9444 4316
rect 9508 4252 9509 4316
rect 9443 4251 9509 4252
rect 9446 2821 9506 4251
rect 9814 3501 9874 6699
rect 10179 6492 10245 6493
rect 10179 6428 10180 6492
rect 10244 6428 10245 6492
rect 10179 6427 10245 6428
rect 9995 5812 10061 5813
rect 9995 5748 9996 5812
rect 10060 5748 10061 5812
rect 9995 5747 10061 5748
rect 9998 3501 10058 5747
rect 10182 4045 10242 6427
rect 11099 6356 11165 6357
rect 11099 6292 11100 6356
rect 11164 6292 11165 6356
rect 11099 6291 11165 6292
rect 11102 4725 11162 6291
rect 11099 4724 11165 4725
rect 11099 4660 11100 4724
rect 11164 4660 11165 4724
rect 11099 4659 11165 4660
rect 10915 4452 10981 4453
rect 10915 4388 10916 4452
rect 10980 4388 10981 4452
rect 10915 4387 10981 4388
rect 11099 4452 11165 4453
rect 11099 4388 11100 4452
rect 11164 4388 11165 4452
rect 11099 4387 11165 4388
rect 10179 4044 10245 4045
rect 10179 3980 10180 4044
rect 10244 3980 10245 4044
rect 10179 3979 10245 3980
rect 9811 3500 9877 3501
rect 9811 3436 9812 3500
rect 9876 3436 9877 3500
rect 9811 3435 9877 3436
rect 9995 3500 10061 3501
rect 9995 3436 9996 3500
rect 10060 3436 10061 3500
rect 9995 3435 10061 3436
rect 9995 3228 10061 3229
rect 9995 3164 9996 3228
rect 10060 3164 10061 3228
rect 9995 3163 10061 3164
rect 9443 2820 9509 2821
rect 9443 2756 9444 2820
rect 9508 2756 9509 2820
rect 9443 2755 9509 2756
rect 9998 2549 10058 3163
rect 10179 2956 10245 2957
rect 10179 2892 10180 2956
rect 10244 2892 10245 2956
rect 10179 2891 10245 2892
rect 9995 2548 10061 2549
rect 9995 2484 9996 2548
rect 10060 2484 10061 2548
rect 9995 2483 10061 2484
rect 9259 2412 9325 2413
rect 9259 2348 9260 2412
rect 9324 2348 9325 2412
rect 9259 2347 9325 2348
rect 10182 2277 10242 2891
rect 10179 2276 10245 2277
rect 10179 2212 10180 2276
rect 10244 2212 10245 2276
rect 10179 2211 10245 2212
rect 10918 2005 10978 4387
rect 11102 3229 11162 4387
rect 11099 3228 11165 3229
rect 11099 3164 11100 3228
rect 11164 3164 11165 3228
rect 11099 3163 11165 3164
rect 11470 2413 11530 6699
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 12019 3908 12085 3909
rect 12019 3844 12020 3908
rect 12084 3844 12085 3908
rect 12019 3843 12085 3844
rect 12022 3365 12082 3843
rect 12019 3364 12085 3365
rect 12019 3300 12020 3364
rect 12084 3300 12085 3364
rect 12019 3299 12085 3300
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 11467 2412 11533 2413
rect 11467 2348 11468 2412
rect 11532 2348 11533 2412
rect 11467 2347 11533 2348
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 48083 26484 48149 26485
rect 48083 26420 48084 26484
rect 48148 26420 48149 26484
rect 48083 26419 48149 26420
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 47163 21316 47229 21317
rect 47163 21252 47164 21316
rect 47228 21252 47229 21316
rect 47163 21251 47229 21252
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 46059 18052 46125 18053
rect 46059 17988 46060 18052
rect 46124 17988 46125 18052
rect 46059 17987 46125 17988
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 46062 12477 46122 17987
rect 47166 17101 47226 21251
rect 47715 20772 47781 20773
rect 47715 20708 47716 20772
rect 47780 20708 47781 20772
rect 47715 20707 47781 20708
rect 47163 17100 47229 17101
rect 47163 17036 47164 17100
rect 47228 17036 47229 17100
rect 47163 17035 47229 17036
rect 47718 16149 47778 20707
rect 47715 16148 47781 16149
rect 47715 16084 47716 16148
rect 47780 16084 47781 16148
rect 47715 16083 47781 16084
rect 46059 12476 46125 12477
rect 46059 12412 46060 12476
rect 46124 12412 46125 12476
rect 46059 12411 46125 12412
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 48086 6493 48146 26419
rect 48083 6492 48149 6493
rect 48083 6428 48084 6492
rect 48148 6428 48149 6492
rect 48083 6427 48149 6428
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 10915 2004 10981 2005
rect 10915 1940 10916 2004
rect 10980 1940 10981 2004
rect 10915 1939 10981 1940
rect 8339 1324 8405 1325
rect 8339 1260 8340 1324
rect 8404 1260 8405 1324
rect 8339 1259 8405 1260
rect 7787 916 7853 917
rect 7787 852 7788 916
rect 7852 852 7853 916
rect 7787 851 7853 852
use sky130_fd_sc_hd__decap_4  FILLER_0_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 2668 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_12
timestamp 1636043612
transform 1 0 2208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1636043612
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 2576 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _113_
timestamp 1636043612
transform -1 0 3312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input136 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_6  input69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 1380 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _112_
timestamp 1636043612
transform -1 0 4232 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 3128 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1636043612
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input104 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 4140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1636043612
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1636043612
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_42
timestamp 1636043612
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39
timestamp 1636043612
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input105
timestamp 1636043612
transform 1 0 5060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _116_
timestamp 1636043612
transform -1 0 5888 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1636043612
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1636043612
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input106
timestamp 1636043612
transform 1 0 6716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _117_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 6532 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1636043612
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1636043612
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1636043612
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1636043612
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input108
timestamp 1636043612
transform 1 0 7636 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1636043612
transform 1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1636043612
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__CLK $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform -1 0 7912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__or4_1  _105_
timestamp 1636043612
transform -1 0 8832 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1636043612
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77
timestamp 1636043612
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1636043612
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_84
timestamp 1636043612
transform 1 0 8832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1636043612
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1636043612
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input110
timestamp 1636043612
transform 1 0 9292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _106_
timestamp 1636043612
transform -1 0 10304 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1636043612
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95
timestamp 1636043612
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__D
timestamp 1636043612
transform -1 0 9384 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1636043612
transform -1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input127
timestamp 1636043612
transform -1 0 11040 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_100
timestamp 1636043612
transform 1 0 10304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1636043612
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1636043612
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input118 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input116
timestamp 1636043612
transform -1 0 12052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1636043612
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1636043612
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1636043612
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp 1636043612
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input124
timestamp 1636043612
transform 1 0 12420 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input121
timestamp 1636043612
transform 1 0 12420 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1636043612
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129
timestamp 1636043612
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform -1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_135
timestamp 1636043612
transform 1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1636043612
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _377_
timestamp 1636043612
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1636043612
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1636043612
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 1636043612
transform -1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_143
timestamp 1636043612
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145
timestamp 1636043612
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output270
timestamp 1636043612
transform -1 0 14996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1636043612
transform -1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_151
timestamp 1636043612
transform 1 0 14996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform -1 0 15824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _246_
timestamp 1636043612
transform -1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp 1636043612
transform 1 0 15640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1636043612
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _255_
timestamp 1636043612
transform -1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _251_
timestamp 1636043612
transform -1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1636043612
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1636043612
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1636043612
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1636043612
transform -1 0 16192 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1636043612
transform 1 0 16928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_172
timestamp 1636043612
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _262_
timestamp 1636043612
transform -1 0 18216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _259_
timestamp 1636043612
transform -1 0 17572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _256_
timestamp 1636043612
transform -1 0 17572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_179
timestamp 1636043612
transform 1 0 17572 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1636043612
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _381_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1636043612
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_187
timestamp 1636043612
transform 1 0 18308 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1636043612
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_186
timestamp 1636043612
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A
timestamp 1636043612
transform -1 0 18768 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _264_
timestamp 1636043612
transform -1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1636043612
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _268_
timestamp 1636043612
transform -1 0 20148 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _266_
timestamp 1636043612
transform -1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_199
timestamp 1636043612
transform 1 0 19412 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_200
timestamp 1636043612
transform 1 0 19504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _383_
timestamp 1636043612
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _271_
timestamp 1636043612
transform -1 0 20792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_211
timestamp 1636043612
transform 1 0 20516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_214
timestamp 1636043612
transform 1 0 20792 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_207
timestamp 1636043612
transform 1 0 20148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _270_
timestamp 1636043612
transform -1 0 21160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1636043612
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _274_
timestamp 1636043612
transform -1 0 22080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1636043612
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1636043612
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1636043612
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1636043612
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _384_
timestamp 1636043612
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _277_
timestamp 1636043612
transform -1 0 22724 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_233
timestamp 1636043612
transform 1 0 22540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_235
timestamp 1636043612
transform 1 0 22724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1636043612
transform 1 0 22080 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _279_
timestamp 1636043612
transform -1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _276_
timestamp 1636043612
transform -1 0 23184 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_240
timestamp 1636043612
transform 1 0 23184 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_239
timestamp 1636043612
transform 1 0 23092 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _386_
timestamp 1636043612
transform 1 0 24012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_248
timestamp 1636043612
transform 1 0 23920 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243
timestamp 1636043612
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _282_
timestamp 1636043612
transform -1 0 25024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _280_
timestamp 1636043612
transform -1 0 24656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1636043612
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_253
timestamp 1636043612
transform 1 0 24380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_256
timestamp 1636043612
transform 1 0 24656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1636043612
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _283_
timestamp 1636043612
transform -1 0 25300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_260
timestamp 1636043612
transform 1 0 25024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _286_
timestamp 1636043612
transform -1 0 25944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _285_
timestamp 1636043612
transform -1 0 25668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_267
timestamp 1636043612
transform 1 0 25668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_270
timestamp 1636043612
transform 1 0 25944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_263
timestamp 1636043612
transform 1 0 25300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _288_
timestamp 1636043612
transform -1 0 26312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp 1636043612
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1636043612
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _292_
timestamp 1636043612
transform -1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _289_
timestamp 1636043612
transform -1 0 27232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1636043612
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1636043612
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _294_
timestamp 1636043612
transform -1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _293_
timestamp 1636043612
transform -1 0 27876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_291
timestamp 1636043612
transform 1 0 27876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_284
timestamp 1636043612
transform 1 0 27232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1636043612
transform 1 0 27876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_284
timestamp 1636043612
transform 1 0 27232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _440_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 28520 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _296_
timestamp 1636043612
transform -1 0 28520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_297
timestamp 1636043612
transform 1 0 28428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_298
timestamp 1636043612
transform 1 0 28520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A
timestamp 1636043612
transform 1 0 28888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1636043612
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1636043612
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_317
timestamp 1636043612
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_324
timestamp 1636043612
transform 1 0 30912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_307
timestamp 1636043612
transform 1 0 29348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1636043612
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _303_
timestamp 1636043612
transform -1 0 30912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _390_
timestamp 1636043612
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_8  _441_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 29716 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _306_
timestamp 1636043612
transform -1 0 31556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1636043612
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_331
timestamp 1636043612
transform 1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _309_
timestamp 1636043612
transform -1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _308_
timestamp 1636043612
transform -1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1636043612
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1636043612
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_340
timestamp 1636043612
transform 1 0 32384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_340
timestamp 1636043612
transform 1 0 32384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1636043612
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _312_
timestamp 1636043612
transform -1 0 33028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _311_
timestamp 1636043612
transform -1 0 33028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_347
timestamp 1636043612
transform 1 0 33028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_347
timestamp 1636043612
transform 1 0 33028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _316_
timestamp 1636043612
transform 1 0 33580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _315_
timestamp 1636043612
transform -1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _313_
timestamp 1636043612
transform -1 0 33672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_354
timestamp 1636043612
transform 1 0 33672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1636043612
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _318_
timestamp 1636043612
transform -1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _317_
timestamp 1636043612
transform -1 0 34960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1636043612
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1636043612
transform 1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_368
timestamp 1636043612
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1636043612
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _395_
timestamp 1636043612
transform 1 0 35880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _322_
timestamp 1636043612
transform -1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _320_
timestamp 1636043612
transform -1 0 35604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_374
timestamp 1636043612
transform 1 0 35512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1636043612
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A
timestamp 1636043612
transform -1 0 35512 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_382
timestamp 1636043612
transform 1 0 36248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_382
timestamp 1636043612
transform 1 0 36248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _326_
timestamp 1636043612
transform -1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _325_
timestamp 1636043612
transform -1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1636043612
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1636043612
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1636043612
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1636043612
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _329_
timestamp 1636043612
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _328_
timestamp 1636043612
transform -1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_396
timestamp 1636043612
transform 1 0 37536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1636043612
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _333_
timestamp 1636043612
transform 1 0 38640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _330_
timestamp 1636043612
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_410
timestamp 1636043612
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1636043612
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_407
timestamp 1636043612
transform 1 0 38548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1636043612
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _332_
timestamp 1636043612
transform -1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_411
timestamp 1636043612
transform 1 0 38916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _336_
timestamp 1636043612
transform -1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _335_
timestamp 1636043612
transform -1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1636043612
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1636043612
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1636043612
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _337_
timestamp 1636043612
transform -1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1636043612
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_424
timestamp 1636043612
transform 1 0 40112 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _340_
timestamp 1636043612
transform 1 0 40756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _339_
timestamp 1636043612
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1636043612
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_434
timestamp 1636043612
transform 1 0 41032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_430
timestamp 1636043612
transform 1 0 40664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _342_
timestamp 1636043612
transform -1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_438
timestamp 1636043612
transform 1 0 41400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_441
timestamp 1636043612
transform 1 0 41676 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A1
timestamp 1636043612
transform -1 0 41952 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _345_
timestamp 1636043612
transform -1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _343_
timestamp 1636043612
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1636043612
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1636043612
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1636043612
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1636043612
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _346_
timestamp 1636043612
transform -1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1636043612
transform 1 0 42688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_452
timestamp 1636043612
transform 1 0 42688 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _349_
timestamp 1636043612
transform 1 0 43240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _351_
timestamp 1636043612
transform 1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _348_
timestamp 1636043612
transform -1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_466
timestamp 1636043612
transform 1 0 43976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp 1636043612
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1636043612
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _350_
timestamp 1636043612
transform -1 0 44620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1636043612
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1636043612
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_468
timestamp 1636043612
transform 1 0 44160 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _353_
timestamp 1636043612
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _352_
timestamp 1636043612
transform -1 0 45264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_480
timestamp 1636043612
transform 1 0 45264 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_480
timestamp 1636043612
transform 1 0 45264 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_492
timestamp 1636043612
transform 1 0 46368 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1636043612
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_488
timestamp 1636043612
transform 1 0 46000 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_492
timestamp 1636043612
transform 1 0 46368 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1636043612
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _237_
timestamp 1636043612
transform 1 0 46092 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1636043612
transform 1 0 46736 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1636043612
transform 1 0 46736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1636043612
transform 1 0 46000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1636043612
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1636043612
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_505
timestamp 1636043612
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_505
timestamp 1636043612
transform 1 0 47564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1636043612
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1636043612
transform 1 0 47840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1636043612
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1636043612
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1636043612
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1636043612
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1636043612
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1636043612
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1636043612
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input103
timestamp 1636043612
transform -1 0 2300 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input125
timestamp 1636043612
transform 1 0 2668 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1636043612
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1636043612
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_35
timestamp 1636043612
transform 1 0 4324 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1636043612
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _114_
timestamp 1636043612
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input107
timestamp 1636043612
transform 1 0 5060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_49
timestamp 1636043612
transform 1 0 5612 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_55
timestamp 1636043612
transform 1 0 6164 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_62
timestamp 1636043612
transform 1 0 6808 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _115_
timestamp 1636043612
transform -1 0 6808 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1636043612
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1636043612
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1636043612
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 7360 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input113
timestamp 1636043612
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_101
timestamp 1636043612
transform 1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_91
timestamp 1636043612
transform 1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input115
timestamp 1636043612
transform 1 0 9844 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input119
timestamp 1636043612
transform 1 0 10764 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_111
timestamp 1636043612
transform 1 0 11316 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_121
timestamp 1636043612
transform 1 0 12236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1636043612
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input123
timestamp 1636043612
transform 1 0 11684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 1636043612
transform -1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1636043612
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_145
timestamp 1636043612
transform 1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_152
timestamp 1636043612
transform 1 0 15088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1636043612
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _239_
timestamp 1636043612
transform -1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _245_
timestamp 1636043612
transform -1 0 15088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output271
timestamp 1636043612
transform -1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1636043612
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1636043612
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1636043612
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _248_
timestamp 1636043612
transform -1 0 15732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _253_
timestamp 1636043612
transform -1 0 16376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _257_
timestamp 1636043612
transform -1 0 17020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1636043612
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1636043612
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1636043612
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1636043612
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _260_
timestamp 1636043612
transform -1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _263_
timestamp 1636043612
transform -1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_200
timestamp 1636043612
transform 1 0 19504 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1636043612
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_214
timestamp 1636043612
transform 1 0 20792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _267_
timestamp 1636043612
transform -1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _269_
timestamp 1636043612
transform -1 0 20148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _272_
timestamp 1636043612
transform -1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _273_
timestamp 1636043612
transform -1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_221
timestamp 1636043612
transform 1 0 21436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_228
timestamp 1636043612
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_235
timestamp 1636043612
transform 1 0 22724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _275_
timestamp 1636043612
transform -1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _278_
timestamp 1636043612
transform -1 0 22724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _281_
timestamp 1636043612
transform 1 0 23092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1636043612
transform 1 0 23736 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_242
timestamp 1636043612
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1636043612
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_256
timestamp 1636043612
transform 1 0 24656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1636043612
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _284_
timestamp 1636043612
transform -1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _287_
timestamp 1636043612
transform -1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_263
timestamp 1636043612
transform 1 0 25300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_267
timestamp 1636043612
transform 1 0 25668 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_271
timestamp 1636043612
transform 1 0 26036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_278
timestamp 1636043612
transform 1 0 26680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_282
timestamp 1636043612
transform 1 0 27048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _290_
timestamp 1636043612
transform 1 0 25760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _291_
timestamp 1636043612
transform -1 0 26680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _295_
timestamp 1636043612
transform 1 0 27140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_286
timestamp 1636043612
transform 1 0 27416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_293
timestamp 1636043612
transform 1 0 28060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp 1636043612
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _297_
timestamp 1636043612
transform 1 0 27784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _298_
timestamp 1636043612
transform -1 0 28704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_312
timestamp 1636043612
transform 1 0 29808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_319
timestamp 1636043612
transform 1 0 30452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_326
timestamp 1636043612
transform 1 0 31096 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1636043612
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _301_
timestamp 1636043612
transform -1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _302_
timestamp 1636043612
transform -1 0 30452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _305_
timestamp 1636043612
transform -1 0 31096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_333
timestamp 1636043612
transform 1 0 31740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_340
timestamp 1636043612
transform 1 0 32384 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_346
timestamp 1636043612
transform 1 0 32936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _307_
timestamp 1636043612
transform -1 0 31740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _310_
timestamp 1636043612
transform -1 0 32384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _314_
timestamp 1636043612
transform -1 0 33304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_350 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 33304 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1636043612
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_368
timestamp 1636043612
transform 1 0 34960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1636043612
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _319_
timestamp 1636043612
transform -1 0 34960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_375
timestamp 1636043612
transform 1 0 35604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_382
timestamp 1636043612
transform 1 0 36248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_389
timestamp 1636043612
transform 1 0 36892 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _321_
timestamp 1636043612
transform -1 0 35604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _323_
timestamp 1636043612
transform -1 0 36248 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _324_
timestamp 1636043612
transform -1 0 36892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _327_
timestamp 1636043612
transform -1 0 37536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_396
timestamp 1636043612
transform 1 0 37536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_400
timestamp 1636043612
transform 1 0 37904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_404
timestamp 1636043612
transform 1 0 38272 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_410
timestamp 1636043612
transform 1 0 38824 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_414
timestamp 1636043612
transform 1 0 39192 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _331_
timestamp 1636043612
transform 1 0 37996 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _334_
timestamp 1636043612
transform 1 0 38916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_421
timestamp 1636043612
transform 1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_427
timestamp 1636043612
transform 1 0 40388 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_433
timestamp 1636043612
transform 1 0 40940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1636043612
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _338_
timestamp 1636043612
transform 1 0 40112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _341_
timestamp 1636043612
transform 1 0 41032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_437
timestamp 1636043612
transform 1 0 41308 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_443
timestamp 1636043612
transform 1 0 41860 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_447
timestamp 1636043612
transform 1 0 42228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_456
timestamp 1636043612
transform 1 0 43056 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _344_
timestamp 1636043612
transform 1 0 41952 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _347_
timestamp 1636043612
transform 1 0 42780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_465
timestamp 1636043612
transform 1 0 43884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1636043612
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1636043612
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform -1 0 45724 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _354_
timestamp 1636043612
transform 1 0 44252 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _355_
timestamp 1636043612
transform 1 0 43608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_485
timestamp 1636043612
transform 1 0 45724 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_493
timestamp 1636043612
transform 1 0 46460 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_497
timestamp 1636043612
transform 1 0 46828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _236_
timestamp 1636043612
transform 1 0 47196 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _238_
timestamp 1636043612
transform 1 0 46552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_504
timestamp 1636043612
transform 1 0 47472 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1636043612
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1636043612
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1636043612
transform 1 0 47840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_14
timestamp 1636043612
transform 1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1636043612
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1636043612
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1636043612
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _111_
timestamp 1636043612
transform 1 0 2760 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input128
timestamp 1636043612
transform 1 0 1840 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__C
timestamp 1636043612
transform 1 0 3680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1636043612
transform 1 0 3312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1636043612
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _442_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 4232 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1636043612
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1636043612
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1636043612
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input109
timestamp 1636043612
transform 1 0 6716 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_67
timestamp 1636043612
transform 1 0 7268 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_84
timestamp 1636043612
transform 1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_4  _180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform -1 0 8832 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1636043612
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_97
timestamp 1636043612
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _184_
timestamp 1636043612
transform 1 0 9200 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input120
timestamp 1636043612
transform 1 0 10396 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1636043612
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1636043612
transform 1 0 11868 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1636043612
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1636043612
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 1636043612
transform -1 0 11868 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1636043612
transform -1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1636043612
transform -1 0 13340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_133
timestamp 1636043612
transform 1 0 13340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_140
timestamp 1636043612
transform 1 0 13984 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp 1636043612
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _240_
timestamp 1636043612
transform -1 0 13984 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _244_
timestamp 1636043612
transform -1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _247_
timestamp 1636043612
transform -1 0 15272 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_154
timestamp 1636043612
transform 1 0 15272 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1636043612
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1636043612
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1636043612
transform 1 0 16928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1636043612
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _252_
timestamp 1636043612
transform -1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _258_
timestamp 1636043612
transform -1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_179
timestamp 1636043612
transform 1 0 17572 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_185
timestamp 1636043612
transform 1 0 18124 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_189
timestamp 1636043612
transform 1 0 18492 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _261_
timestamp 1636043612
transform -1 0 17572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _265_
timestamp 1636043612
transform 1 0 18216 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1636043612
transform 1 0 19964 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_201
timestamp 1636043612
transform 1 0 19596 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_207
timestamp 1636043612
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1636043612
transform 1 0 21988 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1636043612
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1636043612
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1636043612
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_229
timestamp 1636043612
transform 1 0 22172 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1636043612
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_241
timestamp 1636043612
transform 1 0 23276 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_253
timestamp 1636043612
transform 1 0 24380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_265
timestamp 1636043612
transform 1 0 25484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp 1636043612
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_281
timestamp 1636043612
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1636043612
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__A1
timestamp 1636043612
transform -1 0 28060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_289
timestamp 1636043612
transform 1 0 27692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_293
timestamp 1636043612
transform 1 0 28060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_300
timestamp 1636043612
transform 1 0 28704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _299_
timestamp 1636043612
transform 1 0 28428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _300_
timestamp 1636043612
transform -1 0 29348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_307
timestamp 1636043612
transform 1 0 29348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_316
timestamp 1636043612
transform 1 0 30176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_323
timestamp 1636043612
transform 1 0 30820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _304_
timestamp 1636043612
transform 1 0 29900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 30544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1636043612
transform 1 0 31188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1636043612
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1636043612
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1636043612
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1636043612
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1636043612
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1636043612
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1636043612
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1636043612
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1636043612
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1636043612
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1636043612
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1636043612
transform -1 0 41308 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output140_A
timestamp 1636043612
transform -1 0 40756 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output147_A
timestamp 1636043612
transform -1 0 40204 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_417
timestamp 1636043612
transform 1 0 39468 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_425
timestamp 1636043612
transform 1 0 40204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_431
timestamp 1636043612
transform 1 0 40756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_437
timestamp 1636043612
transform 1 0 41308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_444
timestamp 1636043612
transform 1 0 41952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1636043612
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_454
timestamp 1636043612
transform 1 0 42872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1636043612
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _362_
timestamp 1636043612
transform 1 0 43240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _365_
timestamp 1636043612
transform 1 0 42596 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1636043612
transform -1 0 41952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_461
timestamp 1636043612
transform 1 0 43516 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_468
timestamp 1636043612
transform 1 0 44160 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 44528 0 -1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__conb_1  _361_
timestamp 1636043612
transform 1 0 43884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_486
timestamp 1636043612
transform 1 0 45816 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_493
timestamp 1636043612
transform 1 0 46460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1636043612
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _356_
timestamp 1636043612
transform -1 0 46460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _357_
timestamp 1636043612
transform -1 0 47104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_505
timestamp 1636043612
transform 1 0 47564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1636043612
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1636043612
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1636043612
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1636043612
transform 1 0 47840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1636043612
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7
timestamp 1636043612
transform 1 0 1748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1636043612
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input114
timestamp 1636043612
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input129
timestamp 1636043612
transform -1 0 2852 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1636043612
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1636043612
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1636043612
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1636043612
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input131
timestamp 1636043612
transform 1 0 4140 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input133
timestamp 1636043612
transform 1 0 5060 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_49
timestamp 1636043612
transform 1 0 5612 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_55
timestamp 1636043612
transform 1 0 6164 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_62
timestamp 1636043612
transform 1 0 6808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input111
timestamp 1636043612
transform 1 0 6256 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_72
timestamp 1636043612
transform 1 0 7728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1636043612
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1636043612
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _232_
timestamp 1636043612
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input112
timestamp 1636043612
transform 1 0 7176 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1636043612
transform -1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_101
timestamp 1636043612
transform 1 0 10396 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_91
timestamp 1636043612
transform 1 0 9476 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input122
timestamp 1636043612
transform 1 0 9844 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input126
timestamp 1636043612
transform 1 0 10764 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_111
timestamp 1636043612
transform 1 0 11316 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_119
timestamp 1636043612
transform 1 0 12052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_126
timestamp 1636043612
transform 1 0 12696 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _241_
timestamp 1636043612
transform -1 0 12696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _242_
timestamp 1636043612
transform -1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1636043612
transform -1 0 12052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1636043612
transform -1 0 14904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1636043612
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1636043612
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1636043612
transform 1 0 14352 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_150
timestamp 1636043612
transform 1 0 14904 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1636043612
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _249_
timestamp 1636043612
transform -1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output262_A
timestamp 1636043612
transform 1 0 16284 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output267_A
timestamp 1636043612
transform 1 0 16836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_161
timestamp 1636043612
transform 1 0 15916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_167
timestamp 1636043612
transform 1 0 16468 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_173
timestamp 1636043612
transform 1 0 17020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _254_
timestamp 1636043612
transform -1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_185
timestamp 1636043612
transform 1 0 18124 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1636043612
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1636043612
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1636043612
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1636043612
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1636043612
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1636043612
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1636043612
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1636043612
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1636043612
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1636043612
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1636043612
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1636043612
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1636043612
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1636043612
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1636043612
transform 1 0 28796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__A1
timestamp 1636043612
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1636043612
transform -1 0 30912 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_311
timestamp 1636043612
transform 1 0 29716 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_318
timestamp 1636043612
transform 1 0 30360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_324
timestamp 1636043612
transform 1 0 30912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1636043612
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1636043612
transform -1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1636043612
transform -1 0 31464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_330
timestamp 1636043612
transform 1 0 31464 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_342
timestamp 1636043612
transform 1 0 32568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_354
timestamp 1636043612
transform 1 0 33672 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1636043612
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1636043612
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1636043612
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1636043612
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1636043612
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1636043612
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1636043612
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output144_A
timestamp 1636043612
transform -1 0 41032 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output149_A
timestamp 1636043612
transform -1 0 40480 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1636043612
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_421
timestamp 1636043612
transform 1 0 39836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_425
timestamp 1636043612
transform 1 0 40204 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_428
timestamp 1636043612
transform 1 0 40480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_434
timestamp 1636043612
transform 1 0 41032 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1636043612
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A1
timestamp 1636043612
transform -1 0 42136 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A1
timestamp 1636043612
transform -1 0 41584 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_440
timestamp 1636043612
transform 1 0 41584 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_446
timestamp 1636043612
transform 1 0 42136 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_453
timestamp 1636043612
transform 1 0 42780 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _364_
timestamp 1636043612
transform 1 0 43148 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1636043612
transform -1 0 42780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_460
timestamp 1636043612
transform 1 0 43424 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_472
timestamp 1636043612
transform 1 0 44528 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1636043612
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_4  _188_
timestamp 1636043612
transform 1 0 44988 0 1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _191_
timestamp 1636043612
transform -1 0 44528 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_491
timestamp 1636043612
transform 1 0 46276 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_497
timestamp 1636043612
transform 1 0 46828 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_4  _195_
timestamp 1636043612
transform 1 0 46920 0 1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1636043612
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1636043612
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1636043612
transform -1 0 2300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1636043612
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1636043612
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1636043612
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input130
timestamp 1636043612
transform 1 0 2668 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1636043612
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1636043612
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_33
timestamp 1636043612
transform 1 0 4140 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_43
timestamp 1636043612
transform 1 0 5060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input132
timestamp 1636043612
transform 1 0 3588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input134
timestamp 1636043612
transform 1 0 4508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1636043612
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1636043612
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1636043612
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1636043612
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or3_1  _118_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 6716 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1636043612
transform -1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_66
timestamp 1636043612
transform 1 0 7176 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_78
timestamp 1636043612
transform 1 0 8280 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _230_
timestamp 1636043612
transform 1 0 8832 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  input117
timestamp 1636043612
transform 1 0 7728 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__C
timestamp 1636043612
transform 1 0 10856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_102
timestamp 1636043612
transform 1 0 10488 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1636043612
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_89
timestamp 1636043612
transform 1 0 9292 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_95
timestamp 1636043612
transform 1 0 9844 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  _231_
timestamp 1636043612
transform 1 0 9936 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_117
timestamp 1636043612
transform 1 0 11868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_124
timestamp 1636043612
transform 1 0 12512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_131
timestamp 1636043612
transform 1 0 13156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1636043612
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _243_
timestamp 1636043612
transform -1 0 12512 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1636043612
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output268
timestamp 1636043612
transform -1 0 11868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1636043612
transform -1 0 13708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1636043612
transform -1 0 14260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input127_A
timestamp 1636043612
transform -1 0 14812 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_137
timestamp 1636043612
transform 1 0 13708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_143
timestamp 1636043612
transform 1 0 14260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1636043612
transform 1 0 14812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output254_A
timestamp 1636043612
transform 1 0 15180 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output266_A
timestamp 1636043612
transform 1 0 15732 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_155
timestamp 1636043612
transform 1 0 15364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1636043612
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1636043612
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1636043612
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1636043612
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1636043612
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1636043612
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1636043612
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1636043612
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1636043612
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1636043612
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1636043612
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1636043612
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1636043612
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1636043612
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1636043612
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1636043612
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1636043612
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1636043612
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1636043612
transform -1 0 29256 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_293
timestamp 1636043612
transform 1 0 28060 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_301
timestamp 1636043612
transform 1 0 28796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1636043612
transform -1 0 30084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_306
timestamp 1636043612
transform 1 0 29256 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_312
timestamp 1636043612
transform 1 0 29808 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_315
timestamp 1636043612
transform 1 0 30084 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_327
timestamp 1636043612
transform 1 0 31188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1636043612
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1636043612
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1636043612
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1636043612
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1636043612
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1636043612
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1636043612
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1636043612
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1636043612
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1636043612
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1636043612
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output146_A
timestamp 1636043612
transform -1 0 41400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1636043612
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_429
timestamp 1636043612
transform 1 0 40572 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_435
timestamp 1636043612
transform 1 0 41124 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A1
timestamp 1636043612
transform -1 0 42872 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1636043612
transform -1 0 41952 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_438
timestamp 1636043612
transform 1 0 41400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_444
timestamp 1636043612
transform 1 0 41952 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_449
timestamp 1636043612
transform 1 0 42412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_454
timestamp 1636043612
transform 1 0 42872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1636043612
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1636043612
transform -1 0 43516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_461
timestamp 1636043612
transform 1 0 43516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_468
timestamp 1636043612
transform 1 0 44160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _190_
timestamp 1636043612
transform 1 0 44528 0 -1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1636043612
transform -1 0 44160 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_486
timestamp 1636043612
transform 1 0 45816 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_493
timestamp 1636043612
transform 1 0 46460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1636043612
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _358_
timestamp 1636043612
transform -1 0 46460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _359_
timestamp 1636043612
transform -1 0 47104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_508
timestamp 1636043612
transform 1 0 47840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1636043612
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1636043612
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _360_
timestamp 1636043612
transform -1 0 47840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1636043612
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1636043612
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1636043612
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1636043612
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1636043612
transform -1 0 2024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1636043612
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1636043612
transform -1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_14
timestamp 1636043612
transform 1 0 2392 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_10
timestamp 1636043612
transform 1 0 2024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1636043612
transform -1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output272
timestamp 1636043612
transform -1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_19
timestamp 1636043612
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1636043612
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output274
timestamp 1636043612
transform -1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1636043612
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1636043612
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1636043612
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1636043612
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output275
timestamp 1636043612
transform -1 0 4324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform -1 0 4416 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_7_35
timestamp 1636043612
transform 1 0 4324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1636043612
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output277
timestamp 1636043612
transform -1 0 5060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1636043612
transform -1 0 5152 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_36
timestamp 1636043612
transform 1 0 4416 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_43
timestamp 1636043612
transform 1 0 5060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1636043612
transform -1 0 5888 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_44
timestamp 1636043612
transform 1 0 5152 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1636043612
transform -1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1636043612
transform -1 0 6624 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1636043612
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1636043612
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_52
timestamp 1636043612
transform 1 0 5888 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_61
timestamp 1636043612
transform 1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_60
timestamp 1636043612
transform 1 0 6624 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1636043612
transform -1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1636043612
transform -1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _179_
timestamp 1636043612
transform 1 0 7268 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp 1636043612
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_72
timestamp 1636043612
transform 1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_66
timestamp 1636043612
transform 1 0 7176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1636043612
transform -1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_77
timestamp 1636043612
transform 1 0 8188 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1636043612
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1636043612
transform -1 0 9292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1636043612
transform -1 0 9292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1636043612
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1636043612
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _233_
timestamp 1636043612
transform 1 0 9660 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_96
timestamp 1636043612
transform 1 0 9936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_89
timestamp 1636043612
transform 1 0 9292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_89
timestamp 1636043612
transform 1 0 9292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1636043612
transform 1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_103
timestamp 1636043612
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_99
timestamp 1636043612
transform 1 0 10212 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_105
timestamp 1636043612
transform 1 0 10764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 10856 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1636043612
transform -1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1636043612
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1636043612
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1636043612
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_111
timestamp 1636043612
transform 1 0 11316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _100_
timestamp 1636043612
transform 1 0 11960 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp 1636043612
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_118
timestamp 1636043612
transform 1 0 11960 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__B
timestamp 1636043612
transform 1 0 12328 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_124
timestamp 1636043612
transform 1 0 12512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_124
timestamp 1636043612
transform 1 0 12512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input121_A
timestamp 1636043612
transform -1 0 13064 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1636043612
transform -1 0 13064 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_130
timestamp 1636043612
transform 1 0 13064 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_130
timestamp 1636043612
transform 1 0 13064 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1636043612
transform -1 0 13616 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input124_A
timestamp 1636043612
transform -1 0 13616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1636043612
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1636043612
transform 1 0 13616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1636043612
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output264_A
timestamp 1636043612
transform 1 0 13984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_142
timestamp 1636043612
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_143
timestamp 1636043612
transform 1 0 14260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input126_A
timestamp 1636043612
transform -1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_148
timestamp 1636043612
transform 1 0 14720 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1636043612
transform 1 0 14812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output268_A
timestamp 1636043612
transform 1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output253_A
timestamp 1636043612
transform 1 0 14628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output271_A
timestamp 1636043612
transform 1 0 15088 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output261_A
timestamp 1636043612
transform 1 0 15180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output270_A
timestamp 1636043612
transform 1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_155
timestamp 1636043612
transform 1 0 15364 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_161
timestamp 1636043612
transform 1 0 15916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_173
timestamp 1636043612
transform 1 0 17020 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_154
timestamp 1636043612
transform 1 0 15272 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1636043612
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1636043612
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1636043612
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_185
timestamp 1636043612
transform 1 0 18124 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1636043612
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1636043612
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1636043612
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1636043612
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1636043612
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1636043612
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1636043612
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1636043612
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1636043612
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1636043612
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1636043612
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1636043612
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1636043612
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1636043612
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1636043612
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1636043612
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1636043612
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1636043612
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1636043612
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1636043612
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1636043612
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1636043612
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1636043612
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1636043612
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1636043612
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1636043612
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1636043612
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1636043612
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1636043612
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1636043612
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1636043612
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1636043612
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1636043612
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1636043612
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1636043612
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1636043612
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1636043612
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1636043612
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1636043612
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1636043612
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1636043612
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1636043612
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1636043612
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1636043612
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1636043612
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1636043612
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1636043612
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1636043612
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1636043612
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1636043612
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1636043612
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1636043612
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1636043612
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1636043612
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1636043612
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1636043612
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1636043612
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1636043612
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1636043612
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_433
timestamp 1636043612
transform 1 0 40940 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1636043612
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1636043612
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1636043612
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_441
timestamp 1636043612
transform 1 0 41676 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_440
timestamp 1636043612
transform 1 0 41584 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_437
timestamp 1636043612
transform 1 0 41308 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1636043612
transform -1 0 41584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_444
timestamp 1636043612
transform 1 0 41952 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_446
timestamp 1636043612
transform 1 0 42136 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1636043612
transform -1 0 41952 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1636043612
transform -1 0 42136 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1636043612
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_449
timestamp 1636043612
transform 1 0 42412 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1636043612
transform -1 0 42780 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1636043612
transform -1 0 42688 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_453
timestamp 1636043612
transform 1 0 42780 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_452
timestamp 1636043612
transform 1 0 42688 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A1
timestamp 1636043612
transform -1 0 43240 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_458
timestamp 1636043612
transform 1 0 43240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A1
timestamp 1636043612
transform -1 0 43332 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1636043612
transform -1 0 43976 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1636043612
transform -1 0 43884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_459
timestamp 1636043612
transform 1 0 43332 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_466
timestamp 1636043612
transform 1 0 43976 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_465
timestamp 1636043612
transform 1 0 43884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1636043612
transform -1 0 44620 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1636043612
transform -1 0 44528 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_473
timestamp 1636043612
transform 1 0 44620 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_472
timestamp 1636043612
transform 1 0 44528 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1636043612
transform -1 0 45356 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1636043612
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_477
timestamp 1636043612
transform 1 0 44988 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _194_
timestamp 1636043612
transform 1 0 46184 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _183_
timestamp 1636043612
transform -1 0 45724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_485
timestamp 1636043612
transform 1 0 45724 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_481
timestamp 1636043612
transform 1 0 45356 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_489
timestamp 1636043612
transform 1 0 46092 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_485
timestamp 1636043612
transform 1 0 45724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_500
timestamp 1636043612
transform 1 0 47104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_494
timestamp 1636043612
transform 1 0 46552 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _198_
timestamp 1636043612
transform 1 0 45816 0 -1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _196_
timestamp 1636043612
transform 1 0 46920 0 1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1636043612
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_509
timestamp 1636043612
transform 1 0 47932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_515
timestamp 1636043612
transform 1 0 48484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1636043612
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1636043612
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1636043612
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _193_
timestamp 1636043612
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_13
timestamp 1636043612
transform 1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1636043612
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_6
timestamp 1636043612
transform 1 0 1656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1636043612
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _109_
timestamp 1636043612
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _368_
timestamp 1636043612
transform -1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1636043612
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_33
timestamp 1636043612
transform 1 0 4140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1636043612
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1636043612
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output276
timestamp 1636043612
transform -1 0 4140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1636043612
transform -1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_50
timestamp 1636043612
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_57
timestamp 1636043612
transform 1 0 6348 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_64
timestamp 1636043612
transform 1 0 6992 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1636043612
transform 1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1636043612
transform 1 0 6072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1636043612
transform 1 0 6716 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_71
timestamp 1636043612
transform 1 0 7636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_78
timestamp 1636043612
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1636043612
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _110_
timestamp 1636043612
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1636043612
transform 1 0 7360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1636043612
transform 1 0 8004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_102
timestamp 1636043612
transform 1 0 10488 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1636043612
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1636043612
transform 1 0 9200 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_95
timestamp 1636043612
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1636043612
transform 1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1636043612
transform 1 0 10212 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1636043612
transform 1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input123_A
timestamp 1636043612
transform -1 0 12328 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1636043612
transform -1 0 12880 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_116
timestamp 1636043612
transform 1 0 11776 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_122
timestamp 1636043612
transform 1 0 12328 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1636043612
transform 1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1636043612
transform 1 0 11500 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output263_A
timestamp 1636043612
transform 1 0 13248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_134
timestamp 1636043612
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1636043612
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1636043612
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1636043612
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1636043612
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1636043612
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1636043612
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1636043612
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1636043612
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1636043612
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1636043612
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1636043612
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1636043612
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1636043612
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1636043612
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1636043612
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1636043612
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1636043612
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1636043612
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1636043612
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1636043612
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1636043612
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1636043612
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1636043612
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1636043612
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1636043612
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1636043612
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1636043612
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1636043612
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1636043612
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1636043612
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1636043612
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1636043612
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1636043612
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1636043612
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1636043612
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1636043612
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1636043612
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1636043612
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1636043612
transform -1 0 43332 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1636043612
transform -1 0 42780 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_445
timestamp 1636043612
transform 1 0 42044 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_453
timestamp 1636043612
transform 1 0 42780 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A1
timestamp 1636043612
transform -1 0 43884 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_459
timestamp 1636043612
transform 1 0 43332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_465
timestamp 1636043612
transform 1 0 43884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_472
timestamp 1636043612
transform 1 0 44528 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_480
timestamp 1636043612
transform 1 0 45264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1636043612
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1636043612
transform -1 0 45264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1636043612
transform -1 0 44528 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_487
timestamp 1636043612
transform 1 0 45908 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_494
timestamp 1636043612
transform 1 0 46552 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _197_
timestamp 1636043612
transform 1 0 46920 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__conb_1  _366_
timestamp 1636043612
transform 1 0 46276 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1636043612
transform -1 0 45908 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1636043612
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1636043612
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_13
timestamp 1636043612
transform 1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_20
timestamp 1636043612
transform 1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_6
timestamp 1636043612
transform 1 0 1656 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1636043612
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1636043612
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1636043612
transform -1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1636043612
transform 1 0 2668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1636043612
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_38
timestamp 1636043612
transform 1 0 4600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1636043612
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1636043612
transform 1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1636043612
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1636043612
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1636043612
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_60
timestamp 1636043612
transform 1 0 6624 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1636043612
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1636043612
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1636043612
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1636043612
transform 1 0 6992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_67
timestamp 1636043612
transform 1 0 7268 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_76
timestamp 1636043612
transform 1 0 8096 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_83
timestamp 1636043612
transform 1 0 8740 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1636043612
transform -1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1636043612
transform 1 0 8464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1636043612
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1636043612
transform -1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_102
timestamp 1636043612
transform 1 0 10488 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1636043612
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_90
timestamp 1636043612
transform 1 0 9384 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_98
timestamp 1636043612
transform 1 0 10120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1636043612
transform -1 0 10488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1636043612
transform -1 0 11684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1636043612
transform -1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output265_A
timestamp 1636043612
transform 1 0 12604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_115
timestamp 1636043612
transform 1 0 11684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_121
timestamp 1636043612
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1636043612
transform 1 0 12788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1636043612
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1636043612
transform 1 0 13892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_151
timestamp 1636043612
transform 1 0 14996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1636043612
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1636043612
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1636043612
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1636043612
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1636043612
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1636043612
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1636043612
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1636043612
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1636043612
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1636043612
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1636043612
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1636043612
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1636043612
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1636043612
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1636043612
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1636043612
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1636043612
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1636043612
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1636043612
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1636043612
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1636043612
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1636043612
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1636043612
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1636043612
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1636043612
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1636043612
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1636043612
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1636043612
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1636043612
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1636043612
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1636043612
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1636043612
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1636043612
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1636043612
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1636043612
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1636043612
transform 1 0 43240 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1636043612
transform -1 0 42872 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1636043612
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1636043612
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_449
timestamp 1636043612
transform 1 0 42412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_454
timestamp 1636043612
transform 1 0 42872 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1636043612
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_460
timestamp 1636043612
transform 1 0 43424 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_467
timestamp 1636043612
transform 1 0 44068 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_474
timestamp 1636043612
transform 1 0 44712 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1636043612
transform 1 0 44436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1636043612
transform 1 0 43792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _186_
timestamp 1636043612
transform 1 0 45080 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_482
timestamp 1636043612
transform 1 0 45448 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_500
timestamp 1636043612
transform 1 0 47104 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _203_
timestamp 1636043612
transform 1 0 45816 0 -1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_9_508
timestamp 1636043612
transform 1 0 47840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1636043612
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1636043612
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _363_
timestamp 1636043612
transform 1 0 47564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1636043612
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_6
timestamp 1636043612
transform 1 0 1656 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1636043612
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1636043612
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1636043612
transform -1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1636043612
transform -1 0 3128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1636043612
transform -1 0 5244 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_22
timestamp 1636043612
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1636043612
transform 1 0 4048 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_39
timestamp 1636043612
transform 1 0 4692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1636043612
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1636043612
transform 1 0 4416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1636043612
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1636043612
transform -1 0 5796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1636043612
transform -1 0 6716 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_45
timestamp 1636043612
transform 1 0 5244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1636043612
transform 1 0 5796 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_61
timestamp 1636043612
transform 1 0 6716 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1636043612
transform -1 0 7636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1636043612
transform -1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1636043612
transform -1 0 8188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_71
timestamp 1636043612
transform 1 0 7636 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1636043612
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1636043612
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_87
timestamp 1636043612
transform 1 0 9108 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1636043612
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input122_A
timestamp 1636043612
transform -1 0 9844 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1636043612
transform -1 0 10396 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1636043612
transform -1 0 10948 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_101
timestamp 1636043612
transform 1 0 10396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_107
timestamp 1636043612
transform 1 0 10948 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_95
timestamp 1636043612
transform 1 0 9844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1636043612
transform -1 0 11500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_113
timestamp 1636043612
transform 1 0 11500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_125
timestamp 1636043612
transform 1 0 12604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1636043612
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1636043612
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1636043612
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1636043612
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1636043612
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1636043612
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1636043612
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1636043612
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1636043612
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1636043612
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1636043612
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1636043612
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1636043612
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1636043612
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1636043612
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1636043612
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1636043612
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1636043612
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1636043612
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1636043612
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1636043612
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1636043612
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1636043612
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1636043612
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1636043612
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1636043612
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1636043612
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1636043612
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1636043612
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1636043612
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1636043612
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1636043612
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1636043612
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1636043612
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1636043612
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1636043612
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1636043612
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1636043612
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1636043612
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1636043612
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_457
timestamp 1636043612
transform 1 0 43148 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1636043612
transform -1 0 44436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A1
timestamp 1636043612
transform -1 0 45264 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1636043612
transform -1 0 43884 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_465
timestamp 1636043612
transform 1 0 43884 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_471
timestamp 1636043612
transform 1 0 44436 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1636043612
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_477
timestamp 1636043612
transform 1 0 44988 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_480
timestamp 1636043612
transform 1 0 45264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1636043612
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A1
timestamp 1636043612
transform 1 0 46368 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_488
timestamp 1636043612
transform 1 0 46000 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_494
timestamp 1636043612
transform 1 0 46552 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _182_
timestamp 1636043612
transform 1 0 45632 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _199_
timestamp 1636043612
transform 1 0 46920 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1636043612
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1636043612
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1636043612
transform 1 0 2760 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_14
timestamp 1636043612
transform 1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_20
timestamp 1636043612
transform 1 0 2944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_7
timestamp 1636043612
transform 1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1636043612
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _370_
timestamp 1636043612
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1636043612
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1636043612
transform -1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1636043612
transform -1 0 4784 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_24
timestamp 1636043612
transform 1 0 3312 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_28
timestamp 1636043612
transform 1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_34
timestamp 1636043612
transform 1 0 4232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_40
timestamp 1636043612
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1636043612
transform -1 0 3680 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1636043612
transform -1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1636043612
transform -1 0 6716 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1636043612
transform -1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1636043612
transform -1 0 7268 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_46
timestamp 1636043612
transform 1 0 5336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1636043612
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1636043612
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_61
timestamp 1636043612
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1636043612
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1636043612
transform -1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1636043612
transform -1 0 8372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1636043612
transform -1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_67
timestamp 1636043612
transform 1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_73
timestamp 1636043612
transform 1 0 7820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1636043612
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1636043612
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1636043612
transform -1 0 9476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1636043612
transform -1 0 10028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1636043612
transform -1 0 10580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1636043612
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1636043612
transform 1 0 9476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_97
timestamp 1636043612
transform 1 0 10028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1636043612
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1636043612
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1636043612
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1636043612
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1636043612
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1636043612
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1636043612
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1636043612
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1636043612
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1636043612
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1636043612
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1636043612
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1636043612
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1636043612
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1636043612
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1636043612
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1636043612
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1636043612
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1636043612
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1636043612
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1636043612
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1636043612
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1636043612
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1636043612
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1636043612
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1636043612
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1636043612
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1636043612
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1636043612
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1636043612
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1636043612
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1636043612
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1636043612
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1636043612
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1636043612
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1636043612
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1636043612
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1636043612
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1636043612
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1636043612
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1636043612
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1636043612
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1636043612
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1636043612
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1636043612
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A1
timestamp 1636043612
transform -1 0 44804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1636043612
transform -1 0 44252 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_461
timestamp 1636043612
transform 1 0 43516 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_469
timestamp 1636043612
transform 1 0 44252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_475
timestamp 1636043612
transform 1 0 44804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1636043612
transform -1 0 45448 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_482
timestamp 1636043612
transform 1 0 45448 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_500
timestamp 1636043612
transform 1 0 47104 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _204_
timestamp 1636043612
transform 1 0 45816 0 -1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_11_509
timestamp 1636043612
transform 1 0 47932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_515
timestamp 1636043612
transform 1 0 48484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1636043612
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1636043612
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _200_
timestamp 1636043612
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1636043612
transform 1 0 2392 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input125_A
timestamp 1636043612
transform -1 0 3128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_16
timestamp 1636043612
transform 1 0 2576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_6
timestamp 1636043612
transform 1 0 1656 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1636043612
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1636043612
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input129_A
timestamp 1636043612
transform -1 0 3956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input131_A
timestamp 1636043612
transform -1 0 4508 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input133_A
timestamp 1636043612
transform -1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1636043612
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_31
timestamp 1636043612
transform 1 0 3956 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_37
timestamp 1636043612
transform 1 0 4508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_43
timestamp 1636043612
transform 1 0 5060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1636043612
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1636043612
transform -1 0 5612 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1636043612
transform -1 0 6164 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1636043612
transform -1 0 6716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1636043612
transform -1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_49
timestamp 1636043612
transform 1 0 5612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_55
timestamp 1636043612
transform 1 0 6164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_61
timestamp 1636043612
transform 1 0 6716 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1636043612
transform -1 0 7820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1636043612
transform -1 0 8372 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output250_A
timestamp 1636043612
transform -1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_67
timestamp 1636043612
transform 1 0 7268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_73
timestamp 1636043612
transform 1 0 7820 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1636043612
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1636043612
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1636043612
transform 1 0 9108 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1636043612
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output257_A
timestamp 1636043612
transform 1 0 9476 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output260_A
timestamp 1636043612
transform 1 0 10028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1636043612
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_99
timestamp 1636043612
transform 1 0 10212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_111
timestamp 1636043612
transform 1 0 11316 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1636043612
transform 1 0 12420 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 1636043612
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1636043612
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1636043612
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1636043612
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1636043612
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1636043612
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1636043612
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1636043612
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1636043612
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1636043612
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1636043612
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1636043612
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1636043612
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1636043612
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1636043612
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1636043612
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1636043612
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1636043612
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1636043612
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1636043612
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1636043612
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1636043612
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1636043612
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1636043612
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1636043612
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1636043612
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1636043612
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1636043612
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1636043612
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1636043612
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1636043612
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1636043612
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1636043612
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1636043612
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1636043612
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1636043612
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1636043612
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1636043612
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1636043612
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1636043612
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1636043612
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1636043612
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A1
timestamp 1636043612
transform -1 0 45264 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1636043612
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1636043612
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_477
timestamp 1636043612
transform 1 0 44988 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_480
timestamp 1636043612
transform 1 0 45264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1636043612
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A1
timestamp 1636043612
transform -1 0 45816 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_486
timestamp 1636043612
transform 1 0 45816 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_494
timestamp 1636043612
transform 1 0 46552 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _201_
timestamp 1636043612
transform 1 0 46184 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _202_
timestamp 1636043612
transform 1 0 46920 0 1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1636043612
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1636043612
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1636043612
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1636043612
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input135_A
timestamp 1636043612
transform -1 0 1564 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1636043612
transform -1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_5
timestamp 1636043612
transform 1 0 1564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_5
timestamp 1636043612
transform 1 0 1564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input136_A
timestamp 1636043612
transform -1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1636043612
transform -1 0 2116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp 1636043612
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_11
timestamp 1636043612
transform 1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_17
timestamp 1636043612
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_17
timestamp 1636043612
transform 1 0 2668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1636043612
transform -1 0 2668 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input128_A
timestamp 1636043612
transform -1 0 2668 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1636043612
transform -1 0 3220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input130_A
timestamp 1636043612
transform -1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1636043612
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1636043612
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1636043612
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_23
timestamp 1636043612
transform 1 0 3220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input132_A
timestamp 1636043612
transform -1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_31
timestamp 1636043612
transform 1 0 3956 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_29
timestamp 1636043612
transform 1 0 3772 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1636043612
transform -1 0 4508 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1636043612
transform -1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input134_A
timestamp 1636043612
transform -1 0 4508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_37
timestamp 1636043612
transform 1 0 4508 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_37
timestamp 1636043612
transform 1 0 4508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1636043612
transform -1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_43
timestamp 1636043612
transform 1 0 5060 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_43
timestamp 1636043612
transform 1 0 5060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_53
timestamp 1636043612
transform 1 0 5980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_50
timestamp 1636043612
transform 1 0 5704 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_46
timestamp 1636043612
transform 1 0 5336 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_49
timestamp 1636043612
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output249_A
timestamp 1636043612
transform -1 0 5980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output248_A
timestamp 1636043612
transform -1 0 5336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1636043612
transform -1 0 5612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1636043612
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_65
timestamp 1636043612
transform 1 0 7084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_59
timestamp 1636043612
transform 1 0 6532 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1636043612
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output252_A
timestamp 1636043612
transform 1 0 6900 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output251_A
timestamp 1636043612
transform -1 0 6532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1636043612
transform -1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_59
timestamp 1636043612
transform 1 0 6532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_71
timestamp 1636043612
transform 1 0 7636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output256_A
timestamp 1636043612
transform 1 0 8004 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output255_A
timestamp 1636043612
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1636043612
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1636043612
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_77
timestamp 1636043612
transform 1 0 8188 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output259_A
timestamp 1636043612
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1636043612
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_71
timestamp 1636043612
transform 1 0 7636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_83
timestamp 1636043612
transform 1 0 8740 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1636043612
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_95
timestamp 1636043612
transform 1 0 9844 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1636043612
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1636043612
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1636043612
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1636043612
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1636043612
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1636043612
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1636043612
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1636043612
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1636043612
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1636043612
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1636043612
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1636043612
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1636043612
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1636043612
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1636043612
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1636043612
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1636043612
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1636043612
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1636043612
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1636043612
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1636043612
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1636043612
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1636043612
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1636043612
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1636043612
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1636043612
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1636043612
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1636043612
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1636043612
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1636043612
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1636043612
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1636043612
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1636043612
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1636043612
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1636043612
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1636043612
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1636043612
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1636043612
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1636043612
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1636043612
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1636043612
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1636043612
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1636043612
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1636043612
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1636043612
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1636043612
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1636043612
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1636043612
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1636043612
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1636043612
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1636043612
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1636043612
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1636043612
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1636043612
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1636043612
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1636043612
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1636043612
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1636043612
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1636043612
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1636043612
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1636043612
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1636043612
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1636043612
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1636043612
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1636043612
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1636043612
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1636043612
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1636043612
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1636043612
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1636043612
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1636043612
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1636043612
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1636043612
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1636043612
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1636043612
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1636043612
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1636043612
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1636043612
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1636043612
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1636043612
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1636043612
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1636043612
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1636043612
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1636043612
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1636043612
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1636043612
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1636043612
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1636043612
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1636043612
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1636043612
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1636043612
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1636043612
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_477
timestamp 1636043612
transform 1 0 44988 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1636043612
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_476
timestamp 1636043612
transform 1 0 44896 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_473
timestamp 1636043612
transform 1 0 44620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1636043612
transform -1 0 45356 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A1
timestamp 1636043612
transform -1 0 44896 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A1
timestamp 1636043612
transform -1 0 45448 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1636043612
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A1
timestamp 1636043612
transform -1 0 45908 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_482
timestamp 1636043612
transform 1 0 45448 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_500
timestamp 1636043612
transform 1 0 47104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_481
timestamp 1636043612
transform 1 0 45356 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_487
timestamp 1636043612
transform 1 0 45908 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_494
timestamp 1636043612
transform 1 0 46552 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _205_
timestamp 1636043612
transform 1 0 46920 0 1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _206_
timestamp 1636043612
transform 1 0 45816 0 -1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1636043612
transform -1 0 46552 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_505
timestamp 1636043612
transform 1 0 47564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_512
timestamp 1636043612
transform 1 0 48208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1636043612
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1636043612
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1636043612
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1636043612
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1636043612
transform 1 0 47932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1636043612
transform -1 0 1564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1636043612
transform -1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1636043612
transform -1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_11
timestamp 1636043612
transform 1 0 2116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_17
timestamp 1636043612
transform 1 0 2668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_21
timestamp 1636043612
transform 1 0 3036 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_5
timestamp 1636043612
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1636043612
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1636043612
transform -1 0 3312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1636043612
transform -1 0 3864 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output272_A
timestamp 1636043612
transform -1 0 4416 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output275_A
timestamp 1636043612
transform -1 0 4968 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1636043612
transform 1 0 3312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_30
timestamp 1636043612
transform 1 0 3864 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_36
timestamp 1636043612
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_42
timestamp 1636043612
transform 1 0 4968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output277_A
timestamp 1636043612
transform -1 0 5520 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1636043612
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1636043612
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1636043612
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1636043612
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1636043612
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1636043612
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1636043612
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1636043612
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1636043612
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1636043612
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1636043612
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1636043612
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1636043612
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1636043612
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1636043612
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1636043612
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1636043612
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1636043612
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1636043612
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1636043612
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1636043612
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1636043612
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1636043612
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1636043612
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1636043612
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1636043612
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1636043612
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1636043612
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1636043612
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1636043612
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1636043612
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1636043612
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1636043612
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1636043612
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1636043612
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1636043612
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1636043612
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1636043612
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1636043612
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1636043612
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1636043612
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1636043612
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1636043612
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1636043612
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1636043612
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1636043612
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1636043612
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1636043612
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1636043612
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1636043612
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1636043612
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1636043612
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1636043612
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_473
timestamp 1636043612
transform 1 0 44620 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1636043612
transform -1 0 46184 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1636043612
transform -1 0 45632 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_481
timestamp 1636043612
transform 1 0 45356 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_484
timestamp 1636043612
transform 1 0 45632 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_490
timestamp 1636043612
transform 1 0 46184 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_498
timestamp 1636043612
transform 1 0 46920 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _208_
timestamp 1636043612
transform 1 0 46552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1636043612
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_512
timestamp 1636043612
transform 1 0 48208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1636043612
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1636043612
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1636043612
transform 1 0 47932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output247_A
timestamp 1636043612
transform -1 0 1932 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output258_A
timestamp 1636043612
transform -1 0 2668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output273_A
timestamp 1636043612
transform -1 0 3220 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_17
timestamp 1636043612
transform 1 0 2668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1636043612
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_9
timestamp 1636043612
transform 1 0 1932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1636043612
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output274_A
timestamp 1636043612
transform -1 0 3956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output276_A
timestamp 1636043612
transform -1 0 4508 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output278_A
timestamp 1636043612
transform -1 0 5060 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1636043612
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1636043612
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_31
timestamp 1636043612
transform 1 0 3956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_37
timestamp 1636043612
transform 1 0 4508 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_43
timestamp 1636043612
transform 1 0 5060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1636043612
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_55
timestamp 1636043612
transform 1 0 6164 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_67
timestamp 1636043612
transform 1 0 7268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1636043612
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1636043612
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1636043612
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1636043612
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1636043612
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1636043612
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1636043612
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1636043612
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1636043612
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1636043612
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1636043612
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1636043612
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1636043612
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1636043612
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1636043612
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1636043612
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1636043612
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1636043612
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1636043612
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1636043612
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1636043612
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1636043612
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1636043612
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1636043612
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1636043612
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1636043612
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1636043612
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1636043612
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1636043612
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1636043612
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1636043612
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1636043612
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1636043612
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1636043612
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1636043612
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1636043612
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1636043612
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1636043612
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1636043612
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1636043612
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1636043612
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1636043612
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1636043612
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1636043612
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1636043612
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1636043612
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1636043612
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1636043612
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1636043612
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1636043612
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1636043612
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_477
timestamp 1636043612
transform 1 0 44988 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1636043612
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A1
timestamp 1636043612
transform -1 0 45816 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_483
timestamp 1636043612
transform 1 0 45540 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_486
timestamp 1636043612
transform 1 0 45816 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_494
timestamp 1636043612
transform 1 0 46552 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _207_
timestamp 1636043612
transform 1 0 46184 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _209_
timestamp 1636043612
transform 1 0 46920 0 1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1636043612
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1636043612
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output269_A
timestamp 1636043612
transform -1 0 2208 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_12
timestamp 1636043612
transform 1 0 2208 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1636043612
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1636043612
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1636043612
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_24
timestamp 1636043612
transform 1 0 3312 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_36
timestamp 1636043612
transform 1 0 4416 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_48
timestamp 1636043612
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1636043612
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1636043612
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1636043612
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1636043612
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1636043612
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1636043612
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1636043612
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1636043612
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1636043612
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1636043612
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1636043612
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1636043612
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1636043612
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1636043612
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1636043612
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1636043612
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1636043612
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1636043612
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1636043612
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1636043612
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1636043612
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1636043612
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1636043612
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1636043612
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1636043612
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1636043612
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1636043612
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1636043612
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1636043612
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1636043612
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1636043612
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1636043612
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1636043612
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1636043612
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1636043612
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1636043612
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1636043612
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1636043612
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1636043612
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1636043612
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1636043612
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1636043612
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1636043612
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1636043612
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1636043612
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1636043612
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1636043612
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1636043612
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1636043612
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1636043612
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1636043612
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A1
timestamp 1636043612
transform -1 0 45448 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1636043612
transform -1 0 44896 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1636043612
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_473
timestamp 1636043612
transform 1 0 44620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_476
timestamp 1636043612
transform 1 0 44896 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_482
timestamp 1636043612
transform 1 0 45448 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_500
timestamp 1636043612
transform 1 0 47104 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _211_
timestamp 1636043612
transform 1 0 45816 0 -1 11968
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1636043612
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_512
timestamp 1636043612
transform 1 0 48208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1636043612
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1636043612
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1636043612
transform 1 0 47932 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1636043612
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1636043612
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1636043612
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1636043612
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1636043612
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1636043612
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1636043612
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1636043612
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1636043612
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1636043612
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1636043612
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1636043612
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1636043612
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1636043612
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1636043612
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1636043612
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1636043612
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1636043612
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1636043612
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1636043612
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1636043612
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1636043612
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1636043612
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1636043612
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1636043612
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1636043612
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1636043612
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1636043612
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1636043612
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1636043612
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1636043612
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1636043612
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1636043612
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1636043612
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1636043612
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1636043612
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1636043612
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1636043612
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1636043612
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1636043612
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1636043612
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1636043612
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1636043612
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1636043612
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1636043612
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1636043612
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1636043612
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1636043612
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1636043612
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1636043612
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1636043612
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1636043612
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1636043612
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1636043612
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1636043612
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1636043612
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1636043612
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1636043612
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1636043612
transform -1 0 45356 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1636043612
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1636043612
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_477
timestamp 1636043612
transform 1 0 44988 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1636043612
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A1
timestamp 1636043612
transform -1 0 45908 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_481
timestamp 1636043612
transform 1 0 45356 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_487
timestamp 1636043612
transform 1 0 45908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_494
timestamp 1636043612
transform 1 0 46552 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _210_
timestamp 1636043612
transform 1 0 46920 0 1 11968
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1636043612
transform -1 0 46552 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_512
timestamp 1636043612
transform 1 0 48208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1636043612
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1636043612
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1636043612
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1636043612
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1636043612
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1636043612
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1636043612
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1636043612
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1636043612
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1636043612
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1636043612
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1636043612
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1636043612
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1636043612
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1636043612
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1636043612
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1636043612
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1636043612
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1636043612
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1636043612
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1636043612
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1636043612
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1636043612
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1636043612
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1636043612
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1636043612
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1636043612
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1636043612
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1636043612
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1636043612
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1636043612
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1636043612
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1636043612
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1636043612
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1636043612
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1636043612
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1636043612
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1636043612
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1636043612
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1636043612
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1636043612
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1636043612
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1636043612
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1636043612
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1636043612
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1636043612
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1636043612
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1636043612
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1636043612
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1636043612
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1636043612
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1636043612
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1636043612
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1636043612
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1636043612
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1636043612
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1636043612
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1636043612
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1636043612
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1636043612
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1636043612
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1636043612
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1636043612
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1636043612
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1636043612
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1636043612
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1636043612
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1636043612
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1636043612
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1636043612
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1636043612
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1636043612
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1636043612
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1636043612
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1636043612
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1636043612
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1636043612
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1636043612
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1636043612
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1636043612
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1636043612
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1636043612
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1636043612
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1636043612
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1636043612
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1636043612
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1636043612
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1636043612
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1636043612
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1636043612
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1636043612
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1636043612
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1636043612
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1636043612
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1636043612
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1636043612
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1636043612
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1636043612
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1636043612
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1636043612
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1636043612
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1636043612
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1636043612
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1636043612
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1636043612
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1636043612
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1636043612
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1636043612
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1636043612
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1636043612
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1636043612
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1636043612
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1636043612
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1636043612
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1636043612
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1636043612
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1636043612
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_469
timestamp 1636043612
transform 1 0 44252 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1636043612
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_477
timestamp 1636043612
transform 1 0 44988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_472
timestamp 1636043612
transform 1 0 44528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_476
timestamp 1636043612
transform 1 0 44896 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_473
timestamp 1636043612
transform 1 0 44620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1636043612
transform -1 0 44896 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1636043612
transform -1 0 44528 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1636043612
transform -1 0 45356 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A1
timestamp 1636043612
transform -1 0 45448 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1636043612
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A1
timestamp 1636043612
transform -1 0 45908 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_482
timestamp 1636043612
transform 1 0 45448 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_500
timestamp 1636043612
transform 1 0 47104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_481
timestamp 1636043612
transform 1 0 45356 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_487
timestamp 1636043612
transform 1 0 45908 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_494
timestamp 1636043612
transform 1 0 46552 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _212_
timestamp 1636043612
transform 1 0 46920 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _213_
timestamp 1636043612
transform 1 0 45816 0 -1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1636043612
transform -1 0 46552 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_505
timestamp 1636043612
transform 1 0 47564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_512
timestamp 1636043612
transform 1 0 48208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_512
timestamp 1636043612
transform 1 0 48208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1636043612
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1636043612
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1636043612
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1636043612
transform 1 0 47932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1636043612
transform 1 0 2760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_14
timestamp 1636043612
transform 1 0 2392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_20
timestamp 1636043612
transform 1 0 2944 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_7
timestamp 1636043612
transform 1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1636043612
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _371_
timestamp 1636043612
transform 1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1636043612
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_32
timestamp 1636043612
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_44
timestamp 1636043612
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1636043612
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1636043612
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1636043612
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1636043612
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1636043612
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1636043612
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1636043612
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1636043612
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1636043612
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1636043612
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1636043612
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1636043612
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1636043612
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1636043612
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1636043612
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1636043612
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1636043612
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1636043612
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1636043612
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1636043612
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1636043612
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1636043612
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1636043612
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1636043612
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1636043612
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1636043612
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1636043612
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1636043612
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1636043612
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1636043612
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1636043612
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1636043612
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1636043612
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1636043612
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1636043612
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1636043612
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1636043612
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1636043612
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1636043612
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1636043612
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1636043612
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1636043612
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1636043612
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1636043612
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1636043612
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1636043612
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1636043612
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1636043612
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1636043612
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1636043612
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1636043612
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A1
timestamp 1636043612
transform -1 0 45448 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A1
timestamp 1636043612
transform -1 0 44896 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1636043612
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_473
timestamp 1636043612
transform 1 0 44620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_476
timestamp 1636043612
transform 1 0 44896 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_482
timestamp 1636043612
transform 1 0 45448 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_500
timestamp 1636043612
transform 1 0 47104 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _218_
timestamp 1636043612
transform 1 0 45816 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_21_505
timestamp 1636043612
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_512
timestamp 1636043612
transform 1 0 48208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1636043612
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1636043612
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1636043612
transform 1 0 47932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1636043612
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1636043612
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1636043612
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1636043612
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1636043612
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1636043612
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1636043612
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1636043612
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1636043612
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1636043612
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1636043612
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1636043612
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1636043612
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1636043612
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1636043612
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1636043612
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1636043612
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1636043612
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1636043612
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1636043612
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1636043612
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1636043612
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1636043612
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1636043612
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1636043612
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1636043612
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1636043612
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1636043612
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1636043612
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1636043612
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1636043612
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1636043612
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1636043612
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1636043612
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1636043612
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1636043612
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1636043612
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1636043612
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1636043612
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1636043612
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1636043612
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1636043612
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1636043612
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1636043612
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1636043612
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1636043612
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1636043612
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1636043612
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1636043612
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1636043612
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1636043612
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1636043612
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1636043612
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1636043612
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1636043612
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1636043612
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1636043612
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1636043612
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1636043612
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1636043612
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_477
timestamp 1636043612
transform 1 0 44988 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1636043612
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_481
timestamp 1636043612
transform 1 0 45356 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_486
timestamp 1636043612
transform 1 0 45816 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_494
timestamp 1636043612
transform 1 0 46552 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _214_
timestamp 1636043612
transform 1 0 46184 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _215_
timestamp 1636043612
transform 1 0 45448 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _216_
timestamp 1636043612
transform 1 0 46920 0 1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_22_512
timestamp 1636043612
transform 1 0 48208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1636043612
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1636043612
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1636043612
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1636043612
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1636043612
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1636043612
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1636043612
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1636043612
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1636043612
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1636043612
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1636043612
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1636043612
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1636043612
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1636043612
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1636043612
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1636043612
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1636043612
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1636043612
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1636043612
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1636043612
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1636043612
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1636043612
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1636043612
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1636043612
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1636043612
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1636043612
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1636043612
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1636043612
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1636043612
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1636043612
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1636043612
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1636043612
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1636043612
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1636043612
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1636043612
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1636043612
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1636043612
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1636043612
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1636043612
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1636043612
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1636043612
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1636043612
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1636043612
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1636043612
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1636043612
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1636043612
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1636043612
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1636043612
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1636043612
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1636043612
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1636043612
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1636043612
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1636043612
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1636043612
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1636043612
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1636043612
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1636043612
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1636043612
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1636043612
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A1
timestamp 1636043612
transform -1 0 44804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1636043612
transform -1 0 44252 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_461
timestamp 1636043612
transform 1 0 43516 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_469
timestamp 1636043612
transform 1 0 44252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_475
timestamp 1636043612
transform 1 0 44804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1636043612
transform -1 0 45448 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_482
timestamp 1636043612
transform 1 0 45448 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_500
timestamp 1636043612
transform 1 0 47104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _219_
timestamp 1636043612
transform 1 0 45816 0 -1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_23_505
timestamp 1636043612
transform 1 0 47564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_512
timestamp 1636043612
transform 1 0 48208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1636043612
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1636043612
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1636043612
transform 1 0 47932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1636043612
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1636043612
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1636043612
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1636043612
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1636043612
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1636043612
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1636043612
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1636043612
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1636043612
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1636043612
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1636043612
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1636043612
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1636043612
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1636043612
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1636043612
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1636043612
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1636043612
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1636043612
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1636043612
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1636043612
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1636043612
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1636043612
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1636043612
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1636043612
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1636043612
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1636043612
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1636043612
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1636043612
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1636043612
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1636043612
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1636043612
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1636043612
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1636043612
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1636043612
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1636043612
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1636043612
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1636043612
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1636043612
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1636043612
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1636043612
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1636043612
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1636043612
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1636043612
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1636043612
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1636043612
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1636043612
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1636043612
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1636043612
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1636043612
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1636043612
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1636043612
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1636043612
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1636043612
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1636043612
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1636043612
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1636043612
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1636043612
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1636043612
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1636043612
transform -1 0 45356 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1636043612
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1636043612
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_477
timestamp 1636043612
transform 1 0 44988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1636043612
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A1
timestamp 1636043612
transform -1 0 45908 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_481
timestamp 1636043612
transform 1 0 45356 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_487
timestamp 1636043612
transform 1 0 45908 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_494
timestamp 1636043612
transform 1 0 46552 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _217_
timestamp 1636043612
transform 1 0 46920 0 1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1636043612
transform -1 0 46552 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_512
timestamp 1636043612
transform 1 0 48208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1636043612
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1636043612
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1636043612
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1636043612
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1636043612
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1636043612
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1636043612
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1636043612
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1636043612
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1636043612
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1636043612
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1636043612
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1636043612
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1636043612
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1636043612
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1636043612
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1636043612
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1636043612
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1636043612
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1636043612
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1636043612
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1636043612
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1636043612
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1636043612
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1636043612
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1636043612
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1636043612
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1636043612
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1636043612
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1636043612
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1636043612
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1636043612
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1636043612
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1636043612
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1636043612
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1636043612
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1636043612
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1636043612
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1636043612
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1636043612
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1636043612
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1636043612
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1636043612
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1636043612
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1636043612
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1636043612
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1636043612
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1636043612
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1636043612
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1636043612
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1636043612
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1636043612
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1636043612
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1636043612
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1636043612
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1636043612
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1636043612
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1636043612
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1636043612
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1636043612
transform -1 0 44988 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1636043612
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_473
timestamp 1636043612
transform 1 0 44620 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_477
timestamp 1636043612
transform 1 0 44988 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1636043612
transform -1 0 45540 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_483
timestamp 1636043612
transform 1 0 45540 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_490
timestamp 1636043612
transform 1 0 46184 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_498
timestamp 1636043612
transform 1 0 46920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _222_
timestamp 1636043612
transform 1 0 46552 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1636043612
transform -1 0 46184 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_509
timestamp 1636043612
transform 1 0 47932 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_515
timestamp 1636043612
transform 1 0 48484 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1636043612
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1636043612
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _221_
timestamp 1636043612
transform 1 0 47564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1636043612
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1636043612
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1636043612
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1636043612
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1636043612
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1636043612
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1636043612
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1636043612
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1636043612
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1636043612
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1636043612
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1636043612
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1636043612
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1636043612
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1636043612
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1636043612
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1636043612
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1636043612
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1636043612
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1636043612
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1636043612
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1636043612
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1636043612
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1636043612
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1636043612
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1636043612
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1636043612
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1636043612
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1636043612
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1636043612
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1636043612
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1636043612
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1636043612
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1636043612
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1636043612
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1636043612
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1636043612
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1636043612
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1636043612
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1636043612
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1636043612
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1636043612
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1636043612
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1636043612
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1636043612
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1636043612
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1636043612
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1636043612
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1636043612
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1636043612
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1636043612
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1636043612
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1636043612
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1636043612
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1636043612
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1636043612
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1636043612
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1636043612
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1636043612
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1636043612
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1636043612
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1636043612
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1636043612
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1636043612
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1636043612
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1636043612
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1636043612
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1636043612
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1636043612
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1636043612
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1636043612
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1636043612
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1636043612
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1636043612
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1636043612
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1636043612
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1636043612
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1636043612
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1636043612
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1636043612
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1636043612
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1636043612
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1636043612
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1636043612
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1636043612
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1636043612
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1636043612
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1636043612
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1636043612
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1636043612
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1636043612
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1636043612
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1636043612
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1636043612
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1636043612
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1636043612
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1636043612
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1636043612
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1636043612
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1636043612
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1636043612
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1636043612
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1636043612
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1636043612
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1636043612
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1636043612
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1636043612
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1636043612
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1636043612
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1636043612
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1636043612
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1636043612
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1636043612
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1636043612
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1636043612
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1636043612
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A1
timestamp 1636043612
transform -1 0 45448 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1636043612
transform -1 0 45356 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1636043612
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1636043612
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_477
timestamp 1636043612
transform 1 0 44988 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1636043612
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_473
timestamp 1636043612
transform 1 0 44620 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_479
timestamp 1636043612
transform 1 0 45172 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1636043612
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A1
timestamp 1636043612
transform -1 0 45908 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_481
timestamp 1636043612
transform 1 0 45356 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_487
timestamp 1636043612
transform 1 0 45908 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_494
timestamp 1636043612
transform 1 0 46552 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_482
timestamp 1636043612
transform 1 0 45448 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1636043612
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _220_
timestamp 1636043612
transform 1 0 46920 0 1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _224_
timestamp 1636043612
transform 1 0 45816 0 -1 17408
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1636043612
transform -1 0 46552 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1636043612
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_505
timestamp 1636043612
transform 1 0 47564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_512
timestamp 1636043612
transform 1 0 48208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1636043612
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1636043612
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1636043612
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1636043612
transform 1 0 47932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1636043612
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1636043612
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1636043612
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1636043612
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1636043612
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1636043612
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1636043612
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1636043612
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1636043612
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1636043612
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1636043612
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1636043612
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1636043612
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1636043612
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1636043612
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1636043612
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1636043612
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1636043612
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1636043612
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1636043612
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1636043612
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1636043612
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1636043612
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1636043612
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1636043612
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1636043612
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1636043612
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1636043612
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1636043612
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1636043612
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1636043612
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1636043612
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1636043612
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1636043612
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1636043612
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1636043612
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1636043612
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1636043612
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1636043612
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1636043612
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1636043612
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1636043612
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1636043612
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1636043612
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1636043612
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1636043612
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1636043612
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1636043612
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1636043612
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1636043612
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1636043612
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1636043612
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1636043612
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1636043612
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1636043612
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1636043612
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1636043612
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1636043612
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1636043612
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1636043612
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_477
timestamp 1636043612
transform 1 0 44988 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1636043612
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A1
timestamp 1636043612
transform -1 0 46552 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1636043612
transform -1 0 46000 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_485
timestamp 1636043612
transform 1 0 45724 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_488
timestamp 1636043612
transform 1 0 46000 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_494
timestamp 1636043612
transform 1 0 46552 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _223_
timestamp 1636043612
transform 1 0 46920 0 1 17408
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1636043612
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1636043612
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1636043612
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1636043612
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1636043612
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1636043612
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1636043612
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1636043612
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1636043612
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1636043612
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1636043612
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1636043612
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1636043612
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1636043612
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1636043612
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1636043612
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1636043612
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1636043612
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1636043612
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1636043612
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1636043612
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1636043612
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1636043612
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1636043612
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1636043612
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1636043612
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1636043612
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1636043612
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1636043612
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1636043612
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1636043612
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1636043612
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1636043612
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1636043612
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1636043612
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1636043612
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1636043612
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1636043612
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1636043612
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1636043612
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1636043612
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1636043612
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1636043612
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1636043612
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1636043612
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1636043612
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1636043612
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1636043612
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1636043612
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1636043612
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1636043612
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1636043612
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1636043612
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1636043612
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1636043612
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1636043612
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1636043612
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1636043612
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1636043612
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1636043612
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A1
timestamp 1636043612
transform -1 0 45448 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1636043612
transform -1 0 44896 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1636043612
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_473
timestamp 1636043612
transform 1 0 44620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_476
timestamp 1636043612
transform 1 0 44896 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_482
timestamp 1636043612
transform 1 0 45448 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1636043612
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _226_
timestamp 1636043612
transform 1 0 45816 0 -1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_29_505
timestamp 1636043612
transform 1 0 47564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_512
timestamp 1636043612
transform 1 0 48208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1636043612
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1636043612
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1636043612
transform 1 0 47932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1636043612
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1636043612
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1636043612
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1636043612
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1636043612
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1636043612
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1636043612
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1636043612
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1636043612
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1636043612
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1636043612
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1636043612
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1636043612
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1636043612
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1636043612
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1636043612
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1636043612
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1636043612
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1636043612
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1636043612
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1636043612
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1636043612
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1636043612
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1636043612
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1636043612
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1636043612
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1636043612
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1636043612
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1636043612
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1636043612
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1636043612
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1636043612
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1636043612
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1636043612
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1636043612
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1636043612
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1636043612
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1636043612
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1636043612
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1636043612
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1636043612
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1636043612
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1636043612
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1636043612
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1636043612
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1636043612
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1636043612
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1636043612
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1636043612
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1636043612
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1636043612
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1636043612
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1636043612
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1636043612
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1636043612
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1636043612
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1636043612
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1636043612
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1636043612
transform -1 0 45356 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1636043612
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1636043612
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_477
timestamp 1636043612
transform 1 0 44988 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1636043612
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A1
timestamp 1636043612
transform -1 0 45908 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_481
timestamp 1636043612
transform 1 0 45356 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_487
timestamp 1636043612
transform 1 0 45908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_494
timestamp 1636043612
transform 1 0 46552 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _225_
timestamp 1636043612
transform 1 0 46920 0 1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1636043612
transform -1 0 46552 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1636043612
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1636043612
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1636043612
transform 1 0 2576 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_12
timestamp 1636043612
transform 1 0 2208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_18
timestamp 1636043612
transform 1 0 2760 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1636043612
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1636043612
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _373_
timestamp 1636043612
transform 1 0 1932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_30
timestamp 1636043612
transform 1 0 3864 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_42
timestamp 1636043612
transform 1 0 4968 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1636043612
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1636043612
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1636043612
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1636043612
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1636043612
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1636043612
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1636043612
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1636043612
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1636043612
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1636043612
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1636043612
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1636043612
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1636043612
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1636043612
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1636043612
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1636043612
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1636043612
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1636043612
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1636043612
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1636043612
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1636043612
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1636043612
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1636043612
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1636043612
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1636043612
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1636043612
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1636043612
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1636043612
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1636043612
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1636043612
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1636043612
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1636043612
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1636043612
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1636043612
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1636043612
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1636043612
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1636043612
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1636043612
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1636043612
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1636043612
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1636043612
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1636043612
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1636043612
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1636043612
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1636043612
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1636043612
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1636043612
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1636043612
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1636043612
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1636043612
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1636043612
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1636043612
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A1
timestamp 1636043612
transform -1 0 45448 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1636043612
transform -1 0 44896 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1636043612
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_473
timestamp 1636043612
transform 1 0 44620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_476
timestamp 1636043612
transform 1 0 44896 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_482
timestamp 1636043612
transform 1 0 45448 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_500
timestamp 1636043612
transform 1 0 47104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _228_
timestamp 1636043612
transform 1 0 45816 0 -1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_31_505
timestamp 1636043612
transform 1 0 47564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_512
timestamp 1636043612
transform 1 0 48208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1636043612
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1636043612
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1636043612
transform 1 0 47932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp 1636043612
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_7
timestamp 1636043612
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1636043612
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1636043612
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1636043612
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1636043612
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1636043612
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1636043612
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1636043612
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1636043612
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1636043612
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1636043612
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1636043612
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1636043612
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1636043612
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1636043612
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1636043612
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1636043612
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1636043612
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1636043612
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1636043612
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1636043612
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1636043612
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1636043612
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1636043612
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1636043612
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1636043612
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1636043612
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1636043612
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1636043612
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1636043612
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1636043612
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1636043612
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1636043612
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1636043612
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1636043612
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1636043612
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1636043612
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1636043612
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1636043612
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1636043612
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1636043612
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1636043612
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1636043612
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1636043612
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1636043612
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1636043612
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1636043612
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1636043612
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1636043612
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1636043612
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1636043612
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1636043612
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1636043612
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1636043612
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1636043612
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1636043612
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1636043612
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1636043612
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1636043612
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1636043612
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_477
timestamp 1636043612
transform 1 0 44988 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1636043612
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_4  _229_
timestamp 1636043612
transform 1 0 45264 0 1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_32_494
timestamp 1636043612
transform 1 0 46552 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_4  _227_
timestamp 1636043612
transform 1 0 46920 0 1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1636043612
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1636043612
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1636043612
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1636043612
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1636043612
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1636043612
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1636043612
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1636043612
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1636043612
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1636043612
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1636043612
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1636043612
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1636043612
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1636043612
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1636043612
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1636043612
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1636043612
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1636043612
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1636043612
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1636043612
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1636043612
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1636043612
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1636043612
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1636043612
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1636043612
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1636043612
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1636043612
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1636043612
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1636043612
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1636043612
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1636043612
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1636043612
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1636043612
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1636043612
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1636043612
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1636043612
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1636043612
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1636043612
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1636043612
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1636043612
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1636043612
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1636043612
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1636043612
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1636043612
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1636043612
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1636043612
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1636043612
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1636043612
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1636043612
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1636043612
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1636043612
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1636043612
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1636043612
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1636043612
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1636043612
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1636043612
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1636043612
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1636043612
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1636043612
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1636043612
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1636043612
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1636043612
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1636043612
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1636043612
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1636043612
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1636043612
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1636043612
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1636043612
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1636043612
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1636043612
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1636043612
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1636043612
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1636043612
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1636043612
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1636043612
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1636043612
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1636043612
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1636043612
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1636043612
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1636043612
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1636043612
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1636043612
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1636043612
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1636043612
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1636043612
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1636043612
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1636043612
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1636043612
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1636043612
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1636043612
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1636043612
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1636043612
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1636043612
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1636043612
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1636043612
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1636043612
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1636043612
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1636043612
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1636043612
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1636043612
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1636043612
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1636043612
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1636043612
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1636043612
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1636043612
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1636043612
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1636043612
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1636043612
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1636043612
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1636043612
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1636043612
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1636043612
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1636043612
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1636043612
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1636043612
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1636043612
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1636043612
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1636043612
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1636043612
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1636043612
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1636043612
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1636043612
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1636043612
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1636043612
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_485
timestamp 1636043612
transform 1 0 45724 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_492
timestamp 1636043612
transform 1 0 46368 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_489
timestamp 1636043612
transform 1 0 46092 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_494
timestamp 1636043612
transform 1 0 46552 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_491
timestamp 1636043612
transform 1 0 46276 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1636043612
transform -1 0 46368 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A1
timestamp 1636043612
transform 1 0 46368 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_498
timestamp 1636043612
transform 1 0 46920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1636043612
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1636043612
transform -1 0 46920 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A1
timestamp 1636043612
transform -1 0 47104 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1636043612
transform 1 0 47288 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_505
timestamp 1636043612
transform 1 0 47564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_512
timestamp 1636043612
transform 1 0 48208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_505
timestamp 1636043612
transform 1 0 47564 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1636043612
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1636043612
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1636043612
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1636043612
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1636043612
transform 1 0 47932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1636043612
transform 1 0 47932 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1636043612
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1636043612
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1636043612
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1636043612
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1636043612
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1636043612
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1636043612
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1636043612
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1636043612
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1636043612
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1636043612
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1636043612
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1636043612
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1636043612
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1636043612
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1636043612
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1636043612
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1636043612
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1636043612
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1636043612
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1636043612
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1636043612
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1636043612
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1636043612
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1636043612
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1636043612
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1636043612
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1636043612
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1636043612
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1636043612
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1636043612
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1636043612
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1636043612
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1636043612
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1636043612
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1636043612
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1636043612
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1636043612
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1636043612
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1636043612
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1636043612
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1636043612
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1636043612
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1636043612
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1636043612
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1636043612
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1636043612
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1636043612
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1636043612
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1636043612
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1636043612
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1636043612
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1636043612
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1636043612
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1636043612
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1636043612
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1636043612
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1636043612
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1636043612
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1636043612
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1636043612
transform -1 0 47104 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1636043612
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_497
timestamp 1636043612
transform 1 0 46828 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_500
timestamp 1636043612
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_505
timestamp 1636043612
transform 1 0 47564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_512
timestamp 1636043612
transform 1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1636043612
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1636043612
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1636043612
transform -1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1636043612
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1636043612
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1636043612
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1636043612
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1636043612
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1636043612
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1636043612
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1636043612
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1636043612
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1636043612
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1636043612
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1636043612
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1636043612
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1636043612
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1636043612
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1636043612
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1636043612
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1636043612
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1636043612
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1636043612
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1636043612
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1636043612
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1636043612
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1636043612
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1636043612
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1636043612
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1636043612
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1636043612
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1636043612
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1636043612
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1636043612
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1636043612
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1636043612
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1636043612
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1636043612
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1636043612
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1636043612
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1636043612
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1636043612
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1636043612
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1636043612
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1636043612
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1636043612
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1636043612
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1636043612
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1636043612
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1636043612
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1636043612
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1636043612
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1636043612
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1636043612
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1636043612
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1636043612
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1636043612
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1636043612
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1636043612
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1636043612
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1636043612
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1636043612
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1636043612
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1636043612
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1636043612
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1636043612
transform -1 0 47472 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1636043612
transform -1 0 46920 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_489
timestamp 1636043612
transform 1 0 46092 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_495
timestamp 1636043612
transform 1 0 46644 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_498
timestamp 1636043612
transform 1 0 46920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_504
timestamp 1636043612
transform 1 0 47472 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1636043612
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1636043612
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1636043612
transform -1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1636043612
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1636043612
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1636043612
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1636043612
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1636043612
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1636043612
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1636043612
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1636043612
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1636043612
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1636043612
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1636043612
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1636043612
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1636043612
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1636043612
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1636043612
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1636043612
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1636043612
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1636043612
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1636043612
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1636043612
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1636043612
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1636043612
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1636043612
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1636043612
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1636043612
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1636043612
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1636043612
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1636043612
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1636043612
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1636043612
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1636043612
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1636043612
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1636043612
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1636043612
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1636043612
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1636043612
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1636043612
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1636043612
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1636043612
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1636043612
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1636043612
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1636043612
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1636043612
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1636043612
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1636043612
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1636043612
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1636043612
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1636043612
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1636043612
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1636043612
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1636043612
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1636043612
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1636043612
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1636043612
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1636043612
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1636043612
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1636043612
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1636043612
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1636043612
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1636043612
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1636043612
transform -1 0 47104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1636043612
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_497
timestamp 1636043612
transform 1 0 46828 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1636043612
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_505
timestamp 1636043612
transform 1 0 47564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_512
timestamp 1636043612
transform 1 0 48208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1636043612
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1636043612
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1636043612
transform -1 0 48208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1636043612
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1636043612
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1636043612
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1636043612
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1636043612
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1636043612
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1636043612
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1636043612
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1636043612
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1636043612
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1636043612
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1636043612
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1636043612
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1636043612
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1636043612
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1636043612
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1636043612
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1636043612
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1636043612
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1636043612
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1636043612
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1636043612
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1636043612
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1636043612
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1636043612
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1636043612
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1636043612
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1636043612
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1636043612
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1636043612
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1636043612
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1636043612
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1636043612
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1636043612
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1636043612
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1636043612
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1636043612
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1636043612
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1636043612
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1636043612
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1636043612
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1636043612
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1636043612
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1636043612
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1636043612
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1636043612
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1636043612
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1636043612
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1636043612
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1636043612
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1636043612
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1636043612
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1636043612
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1636043612
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1636043612
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1636043612
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1636043612
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1636043612
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1636043612
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1636043612
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1636043612
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1636043612
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1636043612
transform -1 0 47472 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1636043612
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_501
timestamp 1636043612
transform 1 0 47196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_504
timestamp 1636043612
transform 1 0 47472 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1636043612
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1636043612
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1636043612
transform -1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1636043612
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1636043612
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1636043612
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1636043612
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1636043612
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1636043612
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1636043612
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1636043612
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1636043612
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1636043612
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1636043612
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1636043612
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1636043612
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1636043612
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1636043612
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1636043612
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1636043612
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1636043612
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1636043612
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1636043612
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1636043612
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1636043612
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1636043612
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1636043612
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1636043612
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1636043612
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1636043612
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1636043612
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1636043612
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1636043612
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1636043612
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1636043612
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1636043612
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1636043612
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1636043612
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1636043612
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1636043612
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1636043612
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1636043612
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1636043612
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1636043612
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1636043612
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1636043612
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1636043612
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1636043612
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1636043612
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1636043612
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1636043612
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1636043612
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1636043612
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1636043612
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1636043612
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1636043612
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1636043612
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1636043612
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1636043612
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1636043612
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1636043612
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1636043612
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1636043612
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1636043612
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1636043612
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1636043612
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1636043612
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1636043612
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1636043612
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1636043612
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1636043612
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1636043612
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1636043612
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1636043612
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1636043612
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1636043612
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1636043612
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1636043612
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1636043612
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1636043612
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1636043612
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1636043612
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1636043612
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1636043612
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1636043612
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1636043612
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1636043612
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1636043612
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1636043612
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1636043612
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1636043612
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1636043612
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1636043612
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1636043612
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1636043612
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1636043612
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1636043612
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1636043612
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1636043612
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1636043612
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1636043612
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1636043612
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1636043612
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1636043612
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1636043612
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1636043612
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1636043612
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1636043612
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1636043612
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1636043612
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1636043612
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1636043612
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1636043612
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1636043612
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1636043612
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1636043612
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1636043612
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1636043612
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1636043612
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1636043612
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1636043612
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1636043612
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1636043612
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1636043612
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1636043612
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1636043612
transform -1 0 47472 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1636043612
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1636043612
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1636043612
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_501
timestamp 1636043612
transform 1 0 47196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1636043612
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1636043612
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_513
timestamp 1636043612
transform 1 0 48300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_504
timestamp 1636043612
transform 1 0 47472 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1636043612
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1636043612
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1636043612
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1636043612
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1636043612
transform -1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1636043612
transform 1 0 2576 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_12
timestamp 1636043612
transform 1 0 2208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_18
timestamp 1636043612
transform 1 0 2760 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_3
timestamp 1636043612
transform 1 0 1380 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1636043612
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _374_
timestamp 1636043612
transform 1 0 1932 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_30
timestamp 1636043612
transform 1 0 3864 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_42
timestamp 1636043612
transform 1 0 4968 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1636043612
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1636043612
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1636043612
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1636043612
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1636043612
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1636043612
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1636043612
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1636043612
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1636043612
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1636043612
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1636043612
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1636043612
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1636043612
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1636043612
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1636043612
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1636043612
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1636043612
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1636043612
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1636043612
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1636043612
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1636043612
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1636043612
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1636043612
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1636043612
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1636043612
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1636043612
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1636043612
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1636043612
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1636043612
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1636043612
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1636043612
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1636043612
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1636043612
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1636043612
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1636043612
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1636043612
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1636043612
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1636043612
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1636043612
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1636043612
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1636043612
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1636043612
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1636043612
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1636043612
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1636043612
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1636043612
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1636043612
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1636043612
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1636043612
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1636043612
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1636043612
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1636043612
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1636043612
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1636043612
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1636043612
transform -1 0 47104 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1636043612
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_497
timestamp 1636043612
transform 1 0 46828 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1636043612
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_505
timestamp 1636043612
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_512
timestamp 1636043612
transform 1 0 48208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1636043612
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1636043612
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1636043612
transform -1 0 48208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_19
timestamp 1636043612
transform 1 0 2852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_7
timestamp 1636043612
transform 1 0 1748 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1636043612
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1636043612
transform -1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1636043612
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1636043612
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1636043612
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1636043612
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1636043612
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1636043612
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1636043612
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1636043612
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1636043612
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1636043612
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1636043612
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1636043612
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1636043612
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1636043612
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1636043612
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1636043612
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1636043612
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1636043612
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1636043612
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1636043612
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1636043612
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1636043612
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1636043612
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_197
timestamp 1636043612
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_203
timestamp 1636043612
transform 1 0 19780 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform -1 0 21712 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1636043612
transform -1 0 22264 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_224
timestamp 1636043612
transform 1 0 21712 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1636043612
transform 1 0 22264 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_242
timestamp 1636043612
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1636043612
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1636043612
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1636043612
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1636043612
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1636043612
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1636043612
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1636043612
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1636043612
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1636043612
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1636043612
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1636043612
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1636043612
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1636043612
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1636043612
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1636043612
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1636043612
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1636043612
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1636043612
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1636043612
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1636043612
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1636043612
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1636043612
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1636043612
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1636043612
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1636043612
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1636043612
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1636043612
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1636043612
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1636043612
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1636043612
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1636043612
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1636043612
transform -1 0 47472 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1636043612
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_501
timestamp 1636043612
transform 1 0 47196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_504
timestamp 1636043612
transform 1 0 47472 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1636043612
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1636043612
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1636043612
transform -1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1636043612
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1636043612
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1636043612
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1636043612
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1636043612
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1636043612
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1636043612
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1636043612
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1636043612
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1636043612
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1636043612
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1636043612
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1636043612
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1636043612
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1636043612
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1636043612
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1636043612
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1636043612
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1636043612
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1636043612
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1636043612
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1636043612
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1636043612
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1636043612
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1636043612
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1636043612
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1636043612
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1636043612
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1636043612
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1636043612
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1636043612
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1636043612
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1636043612
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1636043612
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1636043612
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1636043612
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1636043612
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1636043612
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1636043612
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1636043612
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1636043612
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1636043612
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1636043612
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1636043612
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1636043612
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1636043612
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1636043612
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1636043612
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1636043612
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1636043612
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1636043612
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1636043612
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1636043612
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1636043612
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1636043612
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1636043612
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1636043612
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1636043612
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1636043612
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1636043612
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1636043612
transform -1 0 47104 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1636043612
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_497
timestamp 1636043612
transform 1 0 46828 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_500
timestamp 1636043612
transform 1 0 47104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_505
timestamp 1636043612
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_512
timestamp 1636043612
transform 1 0 48208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1636043612
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1636043612
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1636043612
transform -1 0 48208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1636043612
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1636043612
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1636043612
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1636043612
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1636043612
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1636043612
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1636043612
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1636043612
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1636043612
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1636043612
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1636043612
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1636043612
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1636043612
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1636043612
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1636043612
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1636043612
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1636043612
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1636043612
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1636043612
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1636043612
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1636043612
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1636043612
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1636043612
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1636043612
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1636043612
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1636043612
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1636043612
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1636043612
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1636043612
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1636043612
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1636043612
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1636043612
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1636043612
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1636043612
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1636043612
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1636043612
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1636043612
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1636043612
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1636043612
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1636043612
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1636043612
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1636043612
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1636043612
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1636043612
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1636043612
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1636043612
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1636043612
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1636043612
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1636043612
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1636043612
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1636043612
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1636043612
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1636043612
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1636043612
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1636043612
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1636043612
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1636043612
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1636043612
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1636043612
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1636043612
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1636043612
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1636043612
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1636043612
transform -1 0 47472 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1636043612
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_501
timestamp 1636043612
transform 1 0 47196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_504
timestamp 1636043612
transform 1 0 47472 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_512
timestamp 1636043612
transform 1 0 48208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1636043612
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1636043612
transform -1 0 48208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1636043612
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1636043612
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1636043612
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1636043612
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1636043612
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1636043612
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1636043612
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1636043612
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1636043612
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1636043612
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1636043612
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1636043612
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1636043612
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1636043612
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1636043612
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1636043612
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1636043612
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1636043612
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1636043612
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1636043612
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1636043612
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1636043612
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1636043612
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1636043612
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1636043612
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1636043612
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1636043612
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1636043612
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1636043612
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1636043612
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1636043612
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1636043612
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1636043612
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1636043612
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1636043612
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1636043612
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1636043612
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1636043612
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1636043612
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1636043612
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1636043612
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1636043612
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1636043612
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1636043612
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1636043612
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1636043612
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1636043612
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1636043612
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1636043612
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1636043612
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1636043612
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1636043612
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1636043612
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1636043612
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1636043612
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1636043612
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1636043612
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1636043612
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1636043612
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1636043612
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1636043612
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1636043612
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1636043612
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_505
timestamp 1636043612
transform 1 0 47564 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_512
timestamp 1636043612
transform 1 0 48208 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1636043612
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1636043612
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1636043612
transform -1 0 48208 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1636043612
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1636043612
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1636043612
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1636043612
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1636043612
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1636043612
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1636043612
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1636043612
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1636043612
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1636043612
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1636043612
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1636043612
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1636043612
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1636043612
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1636043612
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1636043612
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1636043612
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1636043612
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1636043612
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1636043612
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1636043612
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1636043612
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1636043612
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1636043612
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1636043612
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1636043612
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1636043612
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1636043612
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1636043612
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1636043612
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1636043612
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1636043612
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1636043612
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1636043612
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1636043612
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1636043612
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1636043612
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1636043612
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1636043612
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1636043612
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1636043612
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1636043612
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1636043612
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1636043612
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1636043612
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1636043612
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1636043612
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1636043612
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1636043612
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1636043612
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1636043612
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1636043612
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1636043612
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1636043612
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1636043612
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1636043612
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1636043612
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1636043612
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1636043612
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1636043612
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1636043612
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1636043612
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1636043612
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1636043612
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1636043612
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1636043612
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1636043612
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1636043612
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1636043612
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1636043612
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1636043612
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1636043612
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1636043612
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1636043612
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1636043612
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1636043612
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1636043612
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1636043612
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1636043612
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1636043612
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1636043612
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1636043612
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1636043612
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1636043612
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1636043612
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1636043612
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1636043612
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1636043612
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1636043612
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1636043612
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1636043612
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1636043612
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1636043612
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1636043612
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1636043612
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1636043612
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1636043612
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1636043612
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1636043612
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1636043612
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1636043612
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1636043612
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1636043612
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1636043612
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1636043612
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1636043612
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1636043612
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1636043612
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1636043612
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1636043612
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1636043612
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1636043612
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1636043612
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1636043612
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1636043612
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1636043612
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1636043612
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1636043612
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1636043612
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1636043612
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1636043612
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1636043612
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1636043612
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_501
timestamp 1636043612
transform 1 0 47196 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1636043612
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1636043612
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1636043612
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_505
timestamp 1636043612
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1636043612
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_506
timestamp 1636043612
transform 1 0 47656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1636043612
transform -1 0 47656 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1636043612
transform -1 0 48208 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1636043612
transform -1 0 48208 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1636043612
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1636043612
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_512
timestamp 1636043612
transform 1 0 48208 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1636043612
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1636043612
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1636043612
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1636043612
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1636043612
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1636043612
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1636043612
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1636043612
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1636043612
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1636043612
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1636043612
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1636043612
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1636043612
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1636043612
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1636043612
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1636043612
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1636043612
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1636043612
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1636043612
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1636043612
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1636043612
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1636043612
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1636043612
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1636043612
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1636043612
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1636043612
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1636043612
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1636043612
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1636043612
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1636043612
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1636043612
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1636043612
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1636043612
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1636043612
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1636043612
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1636043612
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1636043612
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1636043612
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1636043612
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1636043612
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1636043612
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1636043612
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1636043612
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1636043612
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1636043612
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1636043612
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1636043612
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1636043612
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1636043612
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1636043612
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1636043612
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1636043612
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1636043612
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1636043612
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1636043612
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1636043612
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1636043612
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1636043612
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1636043612
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1636043612
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1636043612
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1636043612
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1636043612
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1636043612
transform -1 0 47472 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1636043612
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_501
timestamp 1636043612
transform 1 0 47196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_504
timestamp 1636043612
transform 1 0 47472 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_512
timestamp 1636043612
transform 1 0 48208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1636043612
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1636043612
transform -1 0 48208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1636043612
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1636043612
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1636043612
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1636043612
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1636043612
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1636043612
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1636043612
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1636043612
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1636043612
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1636043612
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1636043612
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1636043612
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1636043612
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1636043612
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1636043612
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1636043612
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1636043612
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1636043612
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1636043612
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1636043612
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1636043612
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1636043612
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1636043612
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1636043612
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1636043612
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1636043612
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1636043612
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1636043612
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1636043612
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1636043612
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1636043612
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1636043612
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1636043612
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1636043612
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1636043612
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1636043612
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1636043612
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1636043612
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1636043612
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1636043612
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1636043612
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1636043612
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1636043612
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1636043612
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1636043612
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1636043612
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1636043612
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1636043612
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1636043612
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1636043612
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1636043612
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1636043612
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1636043612
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1636043612
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1636043612
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1636043612
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1636043612
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1636043612
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1636043612
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1636043612
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1636043612
transform -1 0 47104 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1636043612
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_497
timestamp 1636043612
transform 1 0 46828 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_500
timestamp 1636043612
transform 1 0 47104 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_505
timestamp 1636043612
transform 1 0 47564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_512
timestamp 1636043612
transform 1 0 48208 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1636043612
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1636043612
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1636043612
transform -1 0 48208 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1636043612
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1636043612
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1636043612
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1636043612
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1636043612
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1636043612
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1636043612
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1636043612
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1636043612
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1636043612
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1636043612
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1636043612
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1636043612
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1636043612
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1636043612
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1636043612
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1636043612
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1636043612
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1636043612
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1636043612
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1636043612
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1636043612
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1636043612
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1636043612
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1636043612
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1636043612
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1636043612
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1636043612
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1636043612
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1636043612
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1636043612
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1636043612
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1636043612
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1636043612
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1636043612
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1636043612
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1636043612
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1636043612
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1636043612
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1636043612
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1636043612
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1636043612
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1636043612
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1636043612
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1636043612
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1636043612
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1636043612
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1636043612
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1636043612
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1636043612
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1636043612
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1636043612
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1636043612
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1636043612
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1636043612
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1636043612
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1636043612
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1636043612
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1636043612
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1636043612
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1636043612
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1636043612
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1636043612
transform -1 0 47472 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1636043612
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1636043612
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_504
timestamp 1636043612
transform 1 0 47472 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1636043612
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1636043612
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1636043612
transform -1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1636043612
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1636043612
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1636043612
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1636043612
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1636043612
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1636043612
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1636043612
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1636043612
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1636043612
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1636043612
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1636043612
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1636043612
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1636043612
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1636043612
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1636043612
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1636043612
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1636043612
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1636043612
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1636043612
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1636043612
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1636043612
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1636043612
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1636043612
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1636043612
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1636043612
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1636043612
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1636043612
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1636043612
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1636043612
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1636043612
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1636043612
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1636043612
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1636043612
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1636043612
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1636043612
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1636043612
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1636043612
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1636043612
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1636043612
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1636043612
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1636043612
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1636043612
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1636043612
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1636043612
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1636043612
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1636043612
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1636043612
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1636043612
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1636043612
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1636043612
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1636043612
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1636043612
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1636043612
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1636043612
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1636043612
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1636043612
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1636043612
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1636043612
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1636043612
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1636043612
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1636043612
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1636043612
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1636043612
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_505
timestamp 1636043612
transform 1 0 47564 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_512
timestamp 1636043612
transform 1 0 48208 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1636043612
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1636043612
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1636043612
transform -1 0 48208 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1636043612
transform -1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1636043612
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1636043612
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_7
timestamp 1636043612
transform 1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _380_
timestamp 1636043612
transform 1 0 2116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_20
timestamp 1636043612
transform 1 0 2944 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_14
timestamp 1636043612
transform 1 0 2392 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A
timestamp 1636043612
transform 1 0 2760 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1636043612
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1636043612
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1636043612
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1636043612
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1636043612
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1636043612
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1636043612
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1636043612
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1636043612
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1636043612
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1636043612
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1636043612
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1636043612
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1636043612
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1636043612
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1636043612
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1636043612
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1636043612
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1636043612
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1636043612
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1636043612
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1636043612
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1636043612
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1636043612
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1636043612
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1636043612
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1636043612
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1636043612
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1636043612
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1636043612
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1636043612
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1636043612
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1636043612
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1636043612
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1636043612
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1636043612
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1636043612
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1636043612
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1636043612
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1636043612
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1636043612
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1636043612
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1636043612
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1636043612
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1636043612
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1636043612
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1636043612
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1636043612
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1636043612
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1636043612
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1636043612
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1636043612
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1636043612
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1636043612
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1636043612
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1636043612
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1636043612
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1636043612
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1636043612
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1636043612
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1636043612
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1636043612
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1636043612
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1636043612
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1636043612
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1636043612
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1636043612
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1636043612
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1636043612
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1636043612
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1636043612
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1636043612
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1636043612
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1636043612
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1636043612
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1636043612
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1636043612
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1636043612
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1636043612
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1636043612
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1636043612
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1636043612
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1636043612
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1636043612
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1636043612
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1636043612
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1636043612
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1636043612
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1636043612
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1636043612
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1636043612
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1636043612
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1636043612
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1636043612
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1636043612
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1636043612
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1636043612
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1636043612
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1636043612
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1636043612
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1636043612
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1636043612
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1636043612
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1636043612
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1636043612
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1636043612
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1636043612
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1636043612
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1636043612
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1636043612
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1636043612
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1636043612
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1636043612
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1636043612
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1636043612
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1636043612
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1636043612
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1636043612
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_501
timestamp 1636043612
transform 1 0 47196 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1636043612
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1636043612
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1636043612
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_505
timestamp 1636043612
transform 1 0 47564 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1636043612
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_506
timestamp 1636043612
transform 1 0 47656 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1636043612
transform -1 0 47656 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1636043612
transform -1 0 48208 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1636043612
transform -1 0 48208 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1636043612
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1636043612
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_512
timestamp 1636043612
transform 1 0 48208 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_512
timestamp 1636043612
transform 1 0 48208 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1636043612
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1636043612
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1636043612
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1636043612
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1636043612
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1636043612
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1636043612
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1636043612
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1636043612
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1636043612
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1636043612
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1636043612
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1636043612
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1636043612
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1636043612
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1636043612
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1636043612
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1636043612
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1636043612
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1636043612
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_153
timestamp 1636043612
transform 1 0 15180 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1636043612
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk
timestamp 1636043612
transform -1 0 16284 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1636043612
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1636043612
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1636043612
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1636043612
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1636043612
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1636043612
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1636043612
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1636043612
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1636043612
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1636043612
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1636043612
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1636043612
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1636043612
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1636043612
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1636043612
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1636043612
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1636043612
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1636043612
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1636043612
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1636043612
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1636043612
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1636043612
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1636043612
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1636043612
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1636043612
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1636043612
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1636043612
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1636043612
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1636043612
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1636043612
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1636043612
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1636043612
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1636043612
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1636043612
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1636043612
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1636043612
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1636043612
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1636043612
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1636043612
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1636043612
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1636043612
transform -1 0 47472 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1636043612
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_501
timestamp 1636043612
transform 1 0 47196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_504
timestamp 1636043612
transform 1 0 47472 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1636043612
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1636043612
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1636043612
transform -1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1636043612
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1636043612
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1636043612
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1636043612
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1636043612
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1636043612
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1636043612
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1636043612
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1636043612
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1636043612
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1636043612
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1636043612
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1636043612
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1636043612
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1636043612
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1636043612
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1636043612
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1636043612
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1636043612
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1636043612
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1636043612
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1636043612
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1636043612
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1636043612
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1636043612
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1636043612
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1636043612
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1636043612
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1636043612
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_237
timestamp 1636043612
transform 1 0 22908 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1636043612
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk
timestamp 1636043612
transform 1 0 23092 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_243
timestamp 1636043612
transform 1 0 23460 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_255
timestamp 1636043612
transform 1 0 24564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_267
timestamp 1636043612
transform 1 0 25668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1636043612
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1636043612
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1636043612
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1636043612
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1636043612
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1636043612
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1636043612
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1636043612
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1636043612
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1636043612
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1636043612
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1636043612
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1636043612
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1636043612
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1636043612
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1636043612
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1636043612
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1636043612
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1636043612
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1636043612
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1636043612
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1636043612
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1636043612
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1636043612
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1636043612
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1636043612
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1636043612
transform -1 0 47104 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1636043612
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_497
timestamp 1636043612
transform 1 0 46828 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1636043612
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_505
timestamp 1636043612
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_512
timestamp 1636043612
transform 1 0 48208 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1636043612
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1636043612
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1636043612
transform -1 0 48208 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1636043612
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1636043612
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1636043612
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1636043612
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1636043612
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1636043612
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1636043612
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1636043612
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1636043612
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1636043612
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1636043612
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1636043612
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1636043612
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1636043612
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1636043612
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1636043612
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1636043612
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1636043612
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1636043612
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1636043612
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1636043612
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1636043612
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1636043612
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1636043612
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1636043612
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1636043612
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1636043612
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1636043612
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1636043612
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1636043612
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1636043612
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1636043612
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1636043612
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1636043612
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1636043612
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1636043612
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1636043612
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1636043612
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1636043612
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1636043612
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1636043612
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1636043612
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1636043612
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1636043612
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1636043612
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1636043612
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1636043612
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1636043612
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1636043612
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1636043612
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1636043612
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1636043612
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1636043612
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1636043612
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1636043612
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1636043612
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1636043612
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1636043612
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1636043612
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1636043612
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1636043612
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1636043612
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1636043612
transform -1 0 47472 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_489
timestamp 1636043612
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_501
timestamp 1636043612
transform 1 0 47196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_504
timestamp 1636043612
transform 1 0 47472 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1636043612
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1636043612
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1636043612
transform -1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1636043612
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1636043612
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1636043612
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1636043612
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1636043612
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1636043612
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1636043612
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1636043612
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1636043612
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1636043612
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1636043612
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1636043612
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1636043612
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1636043612
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1636043612
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1636043612
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1636043612
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1636043612
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1636043612
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1636043612
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1636043612
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1636043612
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1636043612
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1636043612
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1636043612
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1636043612
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1636043612
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1636043612
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1636043612
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1636043612
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1636043612
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1636043612
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1636043612
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1636043612
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1636043612
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1636043612
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1636043612
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1636043612
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1636043612
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1636043612
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1636043612
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1636043612
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1636043612
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1636043612
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1636043612
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1636043612
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1636043612
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1636043612
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1636043612
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1636043612
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1636043612
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1636043612
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1636043612
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1636043612
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1636043612
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1636043612
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1636043612
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1636043612
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1636043612
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1636043612
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1636043612
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1636043612
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1636043612
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_505
timestamp 1636043612
transform 1 0 47564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_512
timestamp 1636043612
transform 1 0 48208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1636043612
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1636043612
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1636043612
transform -1 0 48208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1636043612
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1636043612
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1636043612
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1636043612
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1636043612
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1636043612
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1636043612
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1636043612
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1636043612
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1636043612
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1636043612
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1636043612
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1636043612
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1636043612
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1636043612
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1636043612
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1636043612
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1636043612
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1636043612
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1636043612
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1636043612
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1636043612
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1636043612
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1636043612
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1636043612
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1636043612
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1636043612
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1636043612
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1636043612
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1636043612
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1636043612
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1636043612
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1636043612
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1636043612
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1636043612
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1636043612
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1636043612
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1636043612
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1636043612
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1636043612
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1636043612
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1636043612
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1636043612
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1636043612
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1636043612
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1636043612
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1636043612
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1636043612
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1636043612
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1636043612
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1636043612
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1636043612
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1636043612
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1636043612
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1636043612
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1636043612
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1636043612
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1636043612
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1636043612
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1636043612
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1636043612
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1636043612
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1636043612
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_501
timestamp 1636043612
transform 1 0 47196 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1636043612
transform -1 0 48208 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1636043612
transform -1 0 47656 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_506
timestamp 1636043612
transform 1 0 47656 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1636043612
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1636043612
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1636043612
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1636043612
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1636043612
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1636043612
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1636043612
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1636043612
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1636043612
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1636043612
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1636043612
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1636043612
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1636043612
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1636043612
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1636043612
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1636043612
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1636043612
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1636043612
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1636043612
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1636043612
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1636043612
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1636043612
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1636043612
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1636043612
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1636043612
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1636043612
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1636043612
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1636043612
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1636043612
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1636043612
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1636043612
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1636043612
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1636043612
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1636043612
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1636043612
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1636043612
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1636043612
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1636043612
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1636043612
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1636043612
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1636043612
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1636043612
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1636043612
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1636043612
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1636043612
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1636043612
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1636043612
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1636043612
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1636043612
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1636043612
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1636043612
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1636043612
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1636043612
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1636043612
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1636043612
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1636043612
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1636043612
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1636043612
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1636043612
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1636043612
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1636043612
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1636043612
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1636043612
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1636043612
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1636043612
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1636043612
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1636043612
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1636043612
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1636043612
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1636043612
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1636043612
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1636043612
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1636043612
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1636043612
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1636043612
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1636043612
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1636043612
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1636043612
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1636043612
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1636043612
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1636043612
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1636043612
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1636043612
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1636043612
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1636043612
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1636043612
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1636043612
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1636043612
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1636043612
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1636043612
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1636043612
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1636043612
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1636043612
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1636043612
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1636043612
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1636043612
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1636043612
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1636043612
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1636043612
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1636043612
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1636043612
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1636043612
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1636043612
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1636043612
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1636043612
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1636043612
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1636043612
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1636043612
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1636043612
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1636043612
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1636043612
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1636043612
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1636043612
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1636043612
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1636043612
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1636043612
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1636043612
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1636043612
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1636043612
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1636043612
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1636043612
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1636043612
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1636043612
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1636043612
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1636043612
transform -1 0 47472 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1636043612
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1636043612
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1636043612
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_501
timestamp 1636043612
transform 1 0 47196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1636043612
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_504
timestamp 1636043612
transform 1 0 47472 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_505
timestamp 1636043612
transform 1 0 47564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1636043612
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1636043612
transform -1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1636043612
transform -1 0 48208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1636043612
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1636043612
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1636043612
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_512
timestamp 1636043612
transform 1 0 48208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1636043612
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1636043612
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1636043612
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1636043612
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1636043612
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1636043612
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1636043612
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1636043612
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1636043612
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1636043612
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1636043612
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1636043612
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1636043612
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1636043612
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1636043612
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1636043612
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1636043612
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1636043612
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1636043612
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1636043612
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1636043612
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1636043612
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1636043612
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1636043612
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1636043612
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1636043612
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1636043612
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1636043612
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1636043612
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1636043612
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1636043612
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1636043612
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1636043612
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1636043612
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1636043612
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1636043612
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1636043612
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1636043612
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1636043612
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1636043612
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1636043612
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1636043612
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1636043612
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1636043612
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1636043612
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1636043612
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1636043612
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1636043612
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1636043612
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1636043612
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1636043612
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1636043612
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1636043612
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1636043612
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1636043612
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1636043612
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1636043612
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1636043612
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1636043612
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1636043612
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1636043612
transform -1 0 47104 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1636043612
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_497
timestamp 1636043612
transform 1 0 46828 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_500
timestamp 1636043612
transform 1 0 47104 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_505
timestamp 1636043612
transform 1 0 47564 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_512
timestamp 1636043612
transform 1 0 48208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1636043612
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1636043612
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1636043612
transform -1 0 48208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A
timestamp 1636043612
transform 1 0 2760 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_14
timestamp 1636043612
transform 1 0 2392 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_20
timestamp 1636043612
transform 1 0 2944 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_7
timestamp 1636043612
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1636043612
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _388_
timestamp 1636043612
transform 1 0 2116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1636043612
transform -1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1636043612
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1636043612
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1636043612
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1636043612
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1636043612
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1636043612
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1636043612
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_85
timestamp 1636043612
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1636043612
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_93
timestamp 1636043612
transform 1 0 9660 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_99
timestamp 1636043612
transform 1 0 10212 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_clk
timestamp 1636043612
transform -1 0 10212 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_111
timestamp 1636043612
transform 1 0 11316 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_123
timestamp 1636043612
transform 1 0 12420 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_135
timestamp 1636043612
transform 1 0 13524 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1636043612
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1636043612
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1636043612
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1636043612
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1636043612
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1636043612
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1636043612
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1636043612
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1636043612
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1636043612
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1636043612
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1636043612
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1636043612
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1636043612
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1636043612
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1636043612
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1636043612
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1636043612
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1636043612
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1636043612
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1636043612
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1636043612
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1636043612
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1636043612
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1636043612
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1636043612
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1636043612
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1636043612
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1636043612
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1636043612
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1636043612
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1636043612
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1636043612
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1636043612
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1636043612
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1636043612
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1636043612
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1636043612
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1636043612
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1636043612
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1636043612
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1636043612
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1636043612
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1636043612
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1636043612
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1636043612
transform -1 0 47472 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1636043612
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_501
timestamp 1636043612
transform 1 0 47196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_504
timestamp 1636043612
transform 1 0 47472 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_512
timestamp 1636043612
transform 1 0 48208 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1636043612
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1636043612
transform -1 0 48208 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1636043612
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1636043612
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1636043612
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1636043612
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1636043612
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1636043612
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1636043612
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1636043612
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1636043612
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1636043612
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1636043612
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1636043612
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1636043612
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1636043612
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1636043612
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1636043612
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1636043612
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1636043612
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1636043612
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1636043612
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1636043612
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1636043612
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1636043612
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1636043612
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1636043612
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1636043612
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1636043612
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1636043612
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1636043612
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1636043612
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1636043612
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1636043612
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1636043612
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1636043612
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1636043612
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1636043612
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1636043612
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1636043612
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1636043612
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1636043612
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1636043612
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1636043612
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1636043612
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1636043612
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1636043612
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1636043612
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1636043612
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1636043612
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1636043612
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1636043612
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1636043612
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1636043612
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1636043612
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1636043612
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1636043612
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1636043612
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1636043612
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1636043612
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1636043612
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1636043612
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1636043612
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1636043612
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1636043612
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_505
timestamp 1636043612
transform 1 0 47564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_512
timestamp 1636043612
transform 1 0 48208 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1636043612
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1636043612
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1636043612
transform -1 0 48208 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1636043612
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1636043612
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1636043612
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1636043612
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1636043612
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1636043612
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1636043612
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1636043612
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1636043612
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1636043612
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1636043612
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1636043612
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1636043612
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1636043612
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1636043612
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1636043612
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1636043612
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1636043612
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1636043612
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1636043612
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1636043612
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1636043612
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1636043612
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1636043612
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1636043612
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1636043612
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1636043612
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1636043612
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1636043612
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1636043612
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1636043612
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1636043612
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1636043612
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1636043612
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1636043612
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1636043612
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1636043612
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1636043612
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1636043612
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1636043612
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1636043612
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1636043612
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1636043612
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1636043612
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1636043612
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1636043612
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1636043612
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1636043612
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1636043612
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1636043612
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1636043612
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1636043612
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1636043612
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1636043612
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1636043612
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1636043612
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1636043612
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1636043612
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1636043612
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1636043612
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1636043612
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1636043612
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1636043612
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_501
timestamp 1636043612
transform 1 0 47196 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1636043612
transform -1 0 48208 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1636043612
transform -1 0 47656 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_506
timestamp 1636043612
transform 1 0 47656 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_512
timestamp 1636043612
transform 1 0 48208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1636043612
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1636043612
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1636043612
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1636043612
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1636043612
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1636043612
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1636043612
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1636043612
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1636043612
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1636043612
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1636043612
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1636043612
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1636043612
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1636043612
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1636043612
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1636043612
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1636043612
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1636043612
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1636043612
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1636043612
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1636043612
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1636043612
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1636043612
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1636043612
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1636043612
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1636043612
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1636043612
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1636043612
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1636043612
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1636043612
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1636043612
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1636043612
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1636043612
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1636043612
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1636043612
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1636043612
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1636043612
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1636043612
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1636043612
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1636043612
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1636043612
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1636043612
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1636043612
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1636043612
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1636043612
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1636043612
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1636043612
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1636043612
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1636043612
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1636043612
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1636043612
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1636043612
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1636043612
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1636043612
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1636043612
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1636043612
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1636043612
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1636043612
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1636043612
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1636043612
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1636043612
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1636043612
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1636043612
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1636043612
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_505
timestamp 1636043612
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_512
timestamp 1636043612
transform 1 0 48208 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1636043612
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1636043612
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1636043612
transform -1 0 48208 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1636043612
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1636043612
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1636043612
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1636043612
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1636043612
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1636043612
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1636043612
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1636043612
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1636043612
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1636043612
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1636043612
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1636043612
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1636043612
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1636043612
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1636043612
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1636043612
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1636043612
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1636043612
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1636043612
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1636043612
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1636043612
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1636043612
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1636043612
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1636043612
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1636043612
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1636043612
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1636043612
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1636043612
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1636043612
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1636043612
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1636043612
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1636043612
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1636043612
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1636043612
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1636043612
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1636043612
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1636043612
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1636043612
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1636043612
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1636043612
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1636043612
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1636043612
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1636043612
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1636043612
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1636043612
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1636043612
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1636043612
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1636043612
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1636043612
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1636043612
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1636043612
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1636043612
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1636043612
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1636043612
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1636043612
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1636043612
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1636043612
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1636043612
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1636043612
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1636043612
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1636043612
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1636043612
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1636043612
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1636043612
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1636043612
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1636043612
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1636043612
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1636043612
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1636043612
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1636043612
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1636043612
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1636043612
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1636043612
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_293
timestamp 1636043612
transform 1 0 28060 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_305
timestamp 1636043612
transform 1 0 29164 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1636043612
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1636043612
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_clk
timestamp 1636043612
transform 1 0 27692 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1636043612
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1636043612
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1636043612
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1636043612
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1636043612
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1636043612
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1636043612
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1636043612
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1636043612
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1636043612
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1636043612
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1636043612
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1636043612
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1636043612
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1636043612
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1636043612
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1636043612
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1636043612
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1636043612
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1636043612
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1636043612
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1636043612
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1636043612
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1636043612
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1636043612
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1636043612
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1636043612
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1636043612
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1636043612
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1636043612
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1636043612
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1636043612
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1636043612
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1636043612
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1636043612
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1636043612
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1636043612
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1636043612
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1636043612
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1636043612
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1636043612
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1636043612
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1636043612
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1636043612
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1636043612
transform -1 0 47472 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1636043612
transform -1 0 47104 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_489
timestamp 1636043612
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_501
timestamp 1636043612
transform 1 0 47196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1636043612
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_497
timestamp 1636043612
transform 1 0 46828 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_500
timestamp 1636043612
transform 1 0 47104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_504
timestamp 1636043612
transform 1 0 47472 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1636043612
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_505
timestamp 1636043612
transform 1 0 47564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1636043612
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1636043612
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1636043612
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1636043612
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1636043612
transform -1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1636043612
transform -1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1636043612
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1636043612
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1636043612
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1636043612
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1636043612
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1636043612
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1636043612
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1636043612
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1636043612
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1636043612
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1636043612
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1636043612
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1636043612
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1636043612
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1636043612
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1636043612
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1636043612
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1636043612
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1636043612
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1636043612
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1636043612
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1636043612
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1636043612
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1636043612
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1636043612
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1636043612
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1636043612
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1636043612
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1636043612
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1636043612
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1636043612
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1636043612
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1636043612
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1636043612
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1636043612
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1636043612
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1636043612
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1636043612
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1636043612
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1636043612
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1636043612
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1636043612
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1636043612
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1636043612
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1636043612
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1636043612
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1636043612
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1636043612
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1636043612
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1636043612
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1636043612
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1636043612
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1636043612
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1636043612
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1636043612
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1636043612
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1636043612
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1636043612
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1636043612
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1636043612
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1636043612
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1636043612
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1636043612
transform -1 0 47472 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_489
timestamp 1636043612
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_501
timestamp 1636043612
transform 1 0 47196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_504
timestamp 1636043612
transform 1 0 47472 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1636043612
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1636043612
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1636043612
transform -1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1636043612
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1636043612
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1636043612
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1636043612
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1636043612
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1636043612
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1636043612
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1636043612
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1636043612
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1636043612
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1636043612
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1636043612
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1636043612
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1636043612
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1636043612
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_125
timestamp 1636043612
transform 1 0 12604 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1636043612
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_133
timestamp 1636043612
transform 1 0 13340 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_140
timestamp 1636043612
transform 1 0 13984 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_152
timestamp 1636043612
transform 1 0 15088 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_clk
timestamp 1636043612
transform -1 0 13984 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_164
timestamp 1636043612
transform 1 0 16192 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1636043612
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1636043612
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1636043612
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1636043612
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1636043612
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1636043612
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1636043612
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1636043612
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1636043612
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1636043612
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1636043612
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1636043612
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1636043612
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1636043612
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1636043612
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1636043612
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1636043612
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1636043612
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1636043612
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1636043612
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1636043612
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1636043612
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1636043612
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1636043612
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1636043612
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1636043612
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1636043612
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1636043612
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1636043612
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1636043612
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1636043612
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1636043612
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1636043612
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1636043612
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1636043612
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1636043612
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1636043612
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1636043612
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1636043612
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1636043612
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1636043612
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1636043612
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_505
timestamp 1636043612
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_512
timestamp 1636043612
transform 1 0 48208 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1636043612
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1636043612
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1636043612
transform -1 0 48208 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1636043612
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1636043612
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1636043612
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1636043612
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1636043612
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1636043612
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1636043612
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1636043612
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1636043612
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1636043612
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1636043612
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1636043612
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1636043612
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1636043612
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1636043612
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1636043612
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1636043612
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1636043612
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1636043612
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1636043612
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1636043612
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1636043612
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1636043612
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1636043612
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1636043612
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1636043612
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1636043612
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1636043612
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1636043612
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1636043612
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1636043612
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1636043612
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1636043612
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1636043612
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1636043612
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1636043612
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1636043612
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1636043612
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1636043612
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1636043612
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1636043612
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1636043612
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1636043612
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1636043612
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1636043612
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1636043612
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1636043612
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1636043612
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1636043612
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1636043612
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1636043612
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1636043612
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1636043612
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1636043612
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1636043612
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1636043612
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1636043612
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1636043612
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1636043612
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1636043612
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1636043612
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1636043612
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1636043612
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_501
timestamp 1636043612
transform 1 0 47196 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1636043612
transform -1 0 48208 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1636043612
transform -1 0 47656 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_506
timestamp 1636043612
transform 1 0 47656 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_512
timestamp 1636043612
transform 1 0 48208 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1636043612
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1636043612
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1636043612
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1636043612
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1636043612
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1636043612
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1636043612
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1636043612
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1636043612
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1636043612
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1636043612
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1636043612
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1636043612
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1636043612
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1636043612
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1636043612
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1636043612
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1636043612
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1636043612
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1636043612
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1636043612
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1636043612
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1636043612
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1636043612
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1636043612
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1636043612
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1636043612
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1636043612
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1636043612
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1636043612
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1636043612
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1636043612
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1636043612
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1636043612
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1636043612
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1636043612
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1636043612
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1636043612
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1636043612
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1636043612
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__B2
timestamp 1636043612
transform -1 0 30912 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_317
timestamp 1636043612
transform 1 0 30268 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_321
timestamp 1636043612
transform 1 0 30636 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_324
timestamp 1636043612
transform 1 0 30912 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1636043612
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1636043612
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1636043612
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1636043612
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1636043612
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1636043612
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1636043612
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1636043612
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1636043612
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1636043612
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1636043612
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1636043612
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1636043612
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1636043612
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1636043612
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1636043612
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1636043612
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1636043612
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_485
timestamp 1636043612
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1636043612
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1636043612
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1636043612
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_512
timestamp 1636043612
transform 1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1636043612
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1636043612
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1636043612
transform -1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1636043612
transform -1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _389_
timestamp 1636043612
transform 1 0 1932 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1636043612
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1636043612
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_73_7
timestamp 1636043612
transform 1 0 1748 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_72_3
timestamp 1636043612
transform 1 0 1380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_18
timestamp 1636043612
transform 1 0 2760 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_12
timestamp 1636043612
transform 1 0 2208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1636043612
transform 1 0 2576 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _444_
timestamp 1636043612
transform -1 0 3772 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1636043612
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_29
timestamp 1636043612
transform 1 0 3772 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1636043612
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__C1
timestamp 1636043612
transform -1 0 3956 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__B2
timestamp 1636043612
transform -1 0 3312 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_35
timestamp 1636043612
transform 1 0 4324 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__CLK
timestamp 1636043612
transform 1 0 4692 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A2
timestamp 1636043612
transform 1 0 4140 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_41
timestamp 1636043612
transform 1 0 4876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_43
timestamp 1636043612
transform 1 0 5060 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_31
timestamp 1636043612
transform 1 0 3956 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__B1
timestamp 1636043612
transform 1 0 6348 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_55
timestamp 1636043612
transform 1 0 6164 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_53
timestamp 1636043612
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_59
timestamp 1636043612
transform 1 0 6532 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1636043612
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1636043612
transform 1 0 9108 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__CLK
timestamp 1636043612
transform 1 0 8188 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_67
timestamp 1636043612
transform 1 0 7268 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_79
timestamp 1636043612
transform 1 0 8372 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1636043612
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1636043612
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_71
timestamp 1636043612
transform 1 0 7636 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_73_79
timestamp 1636043612
transform 1 0 8372 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1636043612
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1636043612
transform 1 0 10120 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1636043612
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1636043612
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_100
timestamp 1636043612
transform 1 0 10304 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_89
timestamp 1636043612
transform 1 0 9292 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_97
timestamp 1636043612
transform 1 0 10028 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1636043612
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1636043612
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1636043612
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1636043612
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1636043612
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1636043612
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1636043612
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1636043612
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1636043612
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1636043612
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1636043612
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1636043612
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1636043612
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1636043612
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1636043612
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1636043612
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1636043612
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1636043612
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1636043612
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1636043612
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1636043612
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1636043612
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__B1
timestamp 1636043612
transform 1 0 20148 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1636043612
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1636043612
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_205
timestamp 1636043612
transform 1 0 19964 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_209
timestamp 1636043612
transform 1 0 20332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1636043612
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1636043612
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_221
timestamp 1636043612
transform 1 0 21436 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1636043612
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1636043612
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1636043612
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__B1
timestamp 1636043612
transform 1 0 24196 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1636043612
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1636043612
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1636043612
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_249
timestamp 1636043612
transform 1 0 24012 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_253
timestamp 1636043612
transform 1 0 24380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1636043612
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1636043612
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1636043612
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_265
timestamp 1636043612
transform 1 0 25484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_277
timestamp 1636043612
transform 1 0 26588 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1636043612
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1636043612
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1636043612
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1636043612
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1636043612
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_305
timestamp 1636043612
transform 1 0 29164 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A2
timestamp 1636043612
transform -1 0 30728 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1636043612
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_309
timestamp 1636043612
transform 1 0 29532 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_317
timestamp 1636043612
transform 1 0 30268 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_322
timestamp 1636043612
transform 1 0 30728 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_313
timestamp 1636043612
transform 1 0 29900 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1636043612
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 31096 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _476_
timestamp 1636043612
transform 1 0 30176 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1636043612
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1636043612
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_332
timestamp 1636043612
transform 1 0 31648 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1636043612
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1636043612
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1636043612
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1636043612
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1636043612
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1636043612
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1636043612
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1636043612
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1636043612
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1636043612
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1636043612
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1636043612
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1636043612
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1636043612
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1636043612
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1636043612
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1636043612
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1636043612
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1636043612
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1636043612
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1636043612
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1636043612
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1636043612
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1636043612
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1636043612
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1636043612
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1636043612
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1636043612
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1636043612
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1636043612
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1636043612
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1636043612
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1636043612
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1636043612
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1636043612
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1636043612
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1636043612
transform -1 0 47472 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output137_A
timestamp 1636043612
transform 1 0 46920 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_489
timestamp 1636043612
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_501
timestamp 1636043612
transform 1 0 47196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1636043612
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_497
timestamp 1636043612
transform 1 0 46828 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_500
timestamp 1636043612
transform 1 0 47104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_504
timestamp 1636043612
transform 1 0 47472 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1636043612
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_505
timestamp 1636043612
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_512
timestamp 1636043612
transform 1 0 48208 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1636043612
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1636043612
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1636043612
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1636043612
transform -1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1636043612
transform 1 0 47840 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__B1
timestamp 1636043612
transform -1 0 1932 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_3
timestamp 1636043612
transform 1 0 1380 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_9
timestamp 1636043612
transform 1 0 1932 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1636043612
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform -1 0 3128 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__B1
timestamp 1636043612
transform -1 0 4416 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_22
timestamp 1636043612
transform 1 0 3128 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_29
timestamp 1636043612
transform 1 0 3772 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_33
timestamp 1636043612
transform 1 0 4140 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_36
timestamp 1636043612
transform 1 0 4416 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1636043612
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _173_
timestamp 1636043612
transform 1 0 4784 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_74_49
timestamp 1636043612
transform 1 0 5612 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _171_
timestamp 1636043612
transform 1 0 6348 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1636043612
transform -1 0 7820 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_66
timestamp 1636043612
transform 1 0 7176 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_70
timestamp 1636043612
transform 1 0 7544 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_73
timestamp 1636043612
transform 1 0 7820 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_80
timestamp 1636043612
transform 1 0 8464 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_85
timestamp 1636043612
transform 1 0 8924 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1636043612
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 1636043612
transform 1 0 8188 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_104
timestamp 1636043612
transform 1 0 10672 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_95
timestamp 1636043612
transform 1 0 9844 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_99
timestamp 1636043612
transform 1 0 10212 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _120_
timestamp 1636043612
transform 1 0 9292 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 10304 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__CLK
timestamp 1636043612
transform 1 0 11960 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_116
timestamp 1636043612
transform 1 0 11776 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_120
timestamp 1636043612
transform 1 0 12144 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_132
timestamp 1636043612
transform 1 0 13248 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1636043612
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1636043612
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__B1
timestamp 1636043612
transform -1 0 17204 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1636043612
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_165
timestamp 1636043612
transform 1 0 16284 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_175
timestamp 1636043612
transform 1 0 17204 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_188
timestamp 1636043612
transform 1 0 18400 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1636043612
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _157_
timestamp 1636043612
transform 1 0 17572 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_74_197
timestamp 1636043612
transform 1 0 19228 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_217
timestamp 1636043612
transform 1 0 21068 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _459_
timestamp 1636043612
transform 1 0 19596 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_74_225
timestamp 1636043612
transform 1 0 21804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_236
timestamp 1636043612
transform 1 0 22816 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _144_
timestamp 1636043612
transform 1 0 21896 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_clk
timestamp 1636043612
transform -1 0 23552 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_244
timestamp 1636043612
transform 1 0 23552 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_262
timestamp 1636043612
transform 1 0 25208 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1636043612
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _147_
timestamp 1636043612
transform 1 0 24380 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_74_274
timestamp 1636043612
transform 1 0 26312 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_286
timestamp 1636043612
transform 1 0 27416 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_298
timestamp 1636043612
transform 1 0 28520 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1636043612
transform -1 0 31372 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1636043612
transform 1 0 29808 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_306
timestamp 1636043612
transform 1 0 29256 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_74_309
timestamp 1636043612
transform 1 0 29532 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_74_314
timestamp 1636043612
transform 1 0 29992 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_323
timestamp 1636043612
transform 1 0 30820 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1636043612
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform -1 0 30820 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1636043612
transform 1 0 31924 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_329
timestamp 1636043612
transform 1 0 31372 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_74_337
timestamp 1636043612
transform 1 0 32108 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _475_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636043612
transform 1 0 32660 0 1 42432
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_74_360
timestamp 1636043612
transform 1 0 34224 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_365
timestamp 1636043612
transform 1 0 34684 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1636043612
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _471_
timestamp 1636043612
transform 1 0 34868 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_74_383
timestamp 1636043612
transform 1 0 36340 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_395
timestamp 1636043612
transform 1 0 37444 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_407
timestamp 1636043612
transform 1 0 38548 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1636043612
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1636043612
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1636043612
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1636043612
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1636043612
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1636043612
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1636043612
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1636043612
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1636043612
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1636043612
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output279_A
timestamp 1636043612
transform -1 0 47472 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_489
timestamp 1636043612
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_501
timestamp 1636043612
transform 1 0 47196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_504
timestamp 1636043612
transform 1 0 47472 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1636043612
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1636043612
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1636043612
transform 1 0 47840 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__B1
timestamp 1636043612
transform -1 0 1932 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_3
timestamp 1636043612
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_9
timestamp 1636043612
transform 1 0 1932 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1636043612
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _177_
timestamp 1636043612
transform 1 0 2300 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_75_22
timestamp 1636043612
transform 1 0 3128 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_30
timestamp 1636043612
transform 1 0 3864 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _367_
timestamp 1636043612
transform 1 0 3496 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _447_
timestamp 1636043612
transform 1 0 4416 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_52
timestamp 1636043612
transform 1 0 5888 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_57
timestamp 1636043612
transform 1 0 6348 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1636043612
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _449_
timestamp 1636043612
transform 1 0 6716 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_75_77
timestamp 1636043612
transform 1 0 8188 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_83
timestamp 1636043612
transform 1 0 8740 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _122_
timestamp 1636043612
transform 1 0 8832 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_75_106
timestamp 1636043612
transform 1 0 10856 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_90
timestamp 1636043612
transform 1 0 9384 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_98
timestamp 1636043612
transform 1 0 10120 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1636043612
transform 1 0 9752 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1636043612
transform -1 0 10856 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_113
timestamp 1636043612
transform 1 0 11500 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_121
timestamp 1636043612
transform 1 0 12236 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_129
timestamp 1636043612
transform 1 0 12972 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1636043612
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1636043612
transform 1 0 11868 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _453_
timestamp 1636043612
transform 1 0 13064 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__CLK
timestamp 1636043612
transform 1 0 14904 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_146
timestamp 1636043612
transform 1 0 14536 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_152
timestamp 1636043612
transform 1 0 15088 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__CLK
timestamp 1636043612
transform 1 0 16008 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_160
timestamp 1636043612
transform 1 0 15824 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_164
timestamp 1636043612
transform 1 0 16192 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1636043612
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _456_
timestamp 1636043612
transform 1 0 16652 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_185
timestamp 1636043612
transform 1 0 18124 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _457_
timestamp 1636043612
transform -1 0 19964 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_205
timestamp 1636043612
transform 1 0 19964 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_218
timestamp 1636043612
transform 1 0 21160 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _155_
timestamp 1636043612
transform 1 0 20332 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_75_229
timestamp 1636043612
transform 1 0 22172 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1636043612
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1636043612
transform 1 0 21804 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _462_
timestamp 1636043612
transform 1 0 22908 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_75_253
timestamp 1636043612
transform 1 0 24380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _464_
timestamp 1636043612
transform 1 0 24932 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_275
timestamp 1636043612
transform 1 0 26404 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1636043612
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1636043612
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1636043612
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_293
timestamp 1636043612
transform 1 0 28060 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _466_
timestamp 1636043612
transform 1 0 28152 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_310
timestamp 1636043612
transform 1 0 29624 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_318
timestamp 1636043612
transform 1 0 30360 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_326
timestamp 1636043612
transform 1 0 31096 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1636043612
transform 1 0 29992 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_332
timestamp 1636043612
transform 1 0 31648 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_347
timestamp 1636043612
transform 1 0 33028 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1636043612
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1636043612
transform -1 0 31648 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _123_
timestamp 1636043612
transform 1 0 32108 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__A
timestamp 1636043612
transform -1 0 34316 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__B1
timestamp 1636043612
transform 1 0 35052 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_355
timestamp 1636043612
transform 1 0 33764 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_361
timestamp 1636043612
transform 1 0 34316 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_371
timestamp 1636043612
transform 1 0 35236 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1636043612
transform 1 0 33396 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_384
timestamp 1636043612
transform 1 0 36432 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1636043612
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1636043612
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _129_
timestamp 1636043612
transform 1 0 35604 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1636043612
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1636043612
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1636043612
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1636043612
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1636043612
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1636043612
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1636043612
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1636043612
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1636043612
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output138_A
timestamp 1636043612
transform 1 0 46920 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1636043612
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_497
timestamp 1636043612
transform 1 0 46828 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1636043612
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_505
timestamp 1636043612
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_512
timestamp 1636043612
transform 1 0 48208 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1636043612
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1636043612
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1636043612
transform 1 0 47840 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_3
timestamp 1636043612
transform 1 0 1380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_7
timestamp 1636043612
transform 1 0 1748 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1636043612
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _443_
timestamp 1636043612
transform -1 0 3312 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A2
timestamp 1636043612
transform 1 0 3772 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__C1
timestamp 1636043612
transform 1 0 4324 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1636043612
transform -1 0 5060 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_24
timestamp 1636043612
transform 1 0 3312 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_31
timestamp 1636043612
transform 1 0 3956 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_37
timestamp 1636043612
transform 1 0 4508 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_43
timestamp 1636043612
transform 1 0 5060 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1636043612
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__CLK
timestamp 1636043612
transform 1 0 5888 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_51
timestamp 1636043612
transform 1 0 5796 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_54
timestamp 1636043612
transform 1 0 6072 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1636043612
transform -1 0 8464 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_66
timestamp 1636043612
transform 1 0 7176 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_74
timestamp 1636043612
transform 1 0 7912 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_80
timestamp 1636043612
transform 1 0 8464 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_85
timestamp 1636043612
transform 1 0 8924 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1636043612
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1636043612
transform -1 0 7912 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_101
timestamp 1636043612
transform 1 0 10396 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_93
timestamp 1636043612
transform 1 0 9660 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1636043612
transform 1 0 9292 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _451_
timestamp 1636043612
transform -1 0 11960 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_76_118
timestamp 1636043612
transform 1 0 11960 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_126
timestamp 1636043612
transform 1 0 12696 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _164_
timestamp 1636043612
transform 1 0 12788 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__CLK
timestamp 1636043612
transform 1 0 14076 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_136
timestamp 1636043612
transform 1 0 13616 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_143
timestamp 1636043612
transform 1 0 14260 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1636043612
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_155
timestamp 1636043612
transform 1 0 15364 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_161
timestamp 1636043612
transform 1 0 15916 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1636043612
transform -1 0 15916 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _158_
timestamp 1636043612
transform -1 0 17480 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_76_178
timestamp 1636043612
transform 1 0 17480 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_190
timestamp 1636043612
transform 1 0 18584 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1636043612
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__B1
timestamp 1636043612
transform 1 0 20516 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_207
timestamp 1636043612
transform 1 0 20148 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_213
timestamp 1636043612
transform 1 0 20700 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_217
timestamp 1636043612
transform 1 0 21068 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1636043612
transform -1 0 21528 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _152_
timestamp 1636043612
transform -1 0 20148 0 1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__B1
timestamp 1636043612
transform -1 0 22724 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_222
timestamp 1636043612
transform 1 0 21528 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_230
timestamp 1636043612
transform 1 0 22264 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_235
timestamp 1636043612
transform 1 0 22724 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _149_
timestamp 1636043612
transform -1 0 23920 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_76_248
timestamp 1636043612
transform 1 0 23920 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_262
timestamp 1636043612
transform 1 0 25208 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1636043612
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _145_
timestamp 1636043612
transform 1 0 24380 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_76_274
timestamp 1636043612
transform 1 0 26312 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_282
timestamp 1636043612
transform 1 0 27048 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1636043612
transform 1 0 27232 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_286
timestamp 1636043612
transform 1 0 27416 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_294
timestamp 1636043612
transform 1 0 28152 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_304
timestamp 1636043612
transform 1 0 29072 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _142_
timestamp 1636043612
transform -1 0 29072 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__B1
timestamp 1636043612
transform 1 0 30268 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__B1
timestamp 1636043612
transform -1 0 29716 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_311
timestamp 1636043612
transform 1 0 29716 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_319
timestamp 1636043612
transform 1 0 30452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1636043612
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A2
timestamp 1636043612
transform 1 0 31924 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_331
timestamp 1636043612
transform 1 0 31556 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_337
timestamp 1636043612
transform 1 0 32108 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _127_
timestamp 1636043612
transform -1 0 33304 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_76_350
timestamp 1636043612
transform 1 0 33304 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_362
timestamp 1636043612
transform 1 0 34408 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_76_365
timestamp 1636043612
transform 1 0 34684 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1636043612
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _132_
timestamp 1636043612
transform -1 0 35788 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_76_377
timestamp 1636043612
transform 1 0 35788 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _474_
timestamp 1636043612
transform 1 0 36340 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_399
timestamp 1636043612
transform 1 0 37812 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_411
timestamp 1636043612
transform 1 0 38916 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1636043612
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1636043612
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1636043612
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1636043612
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1636043612
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1636043612
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1636043612
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1636043612
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1636043612
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1636043612
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output145_A
timestamp 1636043612
transform -1 0 46920 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output151_A
timestamp 1636043612
transform -1 0 46368 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output169_A
timestamp 1636043612
transform -1 0 45816 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1636043612
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_486
timestamp 1636043612
transform 1 0 45816 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_492
timestamp 1636043612
transform 1 0 46368 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_498
timestamp 1636043612
transform 1 0 46920 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1636043612
transform 1 0 47288 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output141_A
timestamp 1636043612
transform -1 0 48208 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_506
timestamp 1636043612
transform 1 0 47656 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1636043612
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1636043612
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1636043612
transform 1 0 2576 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A
timestamp 1636043612
transform 1 0 2024 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_12
timestamp 1636043612
transform 1 0 2208 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_18
timestamp 1636043612
transform 1 0 2760 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_3
timestamp 1636043612
transform 1 0 1380 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_9
timestamp 1636043612
transform 1 0 1932 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1636043612
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__B1
timestamp 1636043612
transform -1 0 3864 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__C1
timestamp 1636043612
transform 1 0 4232 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__B2
timestamp 1636043612
transform -1 0 3312 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__CLK
timestamp 1636043612
transform 1 0 4784 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_24
timestamp 1636043612
transform 1 0 3312 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_30
timestamp 1636043612
transform 1 0 3864 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_36
timestamp 1636043612
transform 1 0 4416 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_42
timestamp 1636043612
transform 1 0 4968 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_54
timestamp 1636043612
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_57
timestamp 1636043612
transform 1 0 6348 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_65
timestamp 1636043612
transform 1 0 7084 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1636043612
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1636043612
transform 1 0 7360 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_70
timestamp 1636043612
transform 1 0 7544 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_78
timestamp 1636043612
transform 1 0 8280 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _167_
timestamp 1636043612
transform -1 0 9384 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _372_
timestamp 1636043612
transform 1 0 7912 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__B1
timestamp 1636043612
transform 1 0 10856 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_101
timestamp 1636043612
transform 1 0 10396 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_105
timestamp 1636043612
transform 1 0 10764 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_108
timestamp 1636043612
transform 1 0 11040 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_90
timestamp 1636043612
transform 1 0 9384 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_96
timestamp 1636043612
transform 1 0 9936 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1636043612
transform -1 0 10396 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__B1
timestamp 1636043612
transform -1 0 12880 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_122
timestamp 1636043612
transform 1 0 12328 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_128
timestamp 1636043612
transform 1 0 12880 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1636043612
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _166_
timestamp 1636043612
transform -1 0 12328 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1636043612
transform 1 0 13708 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A
timestamp 1636043612
transform 1 0 14996 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_136
timestamp 1636043612
transform 1 0 13616 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_139
timestamp 1636043612
transform 1 0 13892 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_147
timestamp 1636043612
transform 1 0 14628 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1636043612
transform 1 0 14260 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__B1
timestamp 1636043612
transform -1 0 16836 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__CLK
timestamp 1636043612
transform 1 0 15732 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_153
timestamp 1636043612
transform 1 0 15180 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1636043612
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1636043612
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_171
timestamp 1636043612
transform 1 0 16836 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1636043612
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1636043612
transform 1 0 18860 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A
timestamp 1636043612
transform 1 0 18032 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_183
timestamp 1636043612
transform 1 0 17940 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_186
timestamp 1636043612
transform 1 0 18216 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_192
timestamp 1636043612
transform 1 0 18768 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_195
timestamp 1636043612
transform 1 0 19044 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_203
timestamp 1636043612
transform 1 0 19780 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_216
timestamp 1636043612
transform 1 0 20976 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1636043612
transform 1 0 19412 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _153_
timestamp 1636043612
transform 1 0 20148 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1636043612
transform 1 0 22908 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_225
timestamp 1636043612
transform 1 0 21804 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_233
timestamp 1636043612
transform 1 0 22540 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_239
timestamp 1636043612
transform 1 0 23092 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1636043612
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1636043612
transform 1 0 22172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__B1
timestamp 1636043612
transform -1 0 24380 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_247
timestamp 1636043612
transform 1 0 23828 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_253
timestamp 1636043612
transform 1 0 24380 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_259
timestamp 1636043612
transform 1 0 24932 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1636043612
transform 1 0 23460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _465_
timestamp 1636043612
transform 1 0 25024 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_77_276
timestamp 1636043612
transform 1 0 26496 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_281
timestamp 1636043612
transform 1 0 26956 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1636043612
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_285
timestamp 1636043612
transform 1 0 27324 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_290
timestamp 1636043612
transform 1 0 27784 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1636043612
transform 1 0 27416 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _135_
timestamp 1636043612
transform 1 0 28336 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1636043612
transform 1 0 29624 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_306
timestamp 1636043612
transform 1 0 29256 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_312
timestamp 1636043612
transform 1 0 29808 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_318
timestamp 1636043612
transform 1 0 30360 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _140_
timestamp 1636043612
transform -1 0 31280 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_77_328
timestamp 1636043612
transform 1 0 31280 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1636043612
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_349
timestamp 1636043612
transform 1 0 33212 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1636043612
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__B1
timestamp 1636043612
transform -1 0 34960 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A
timestamp 1636043612
transform 1 0 34132 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_357
timestamp 1636043612
transform 1 0 33948 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_361
timestamp 1636043612
transform 1 0 34316 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_365
timestamp 1636043612
transform 1 0 34684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_368
timestamp 1636043612
transform 1 0 34960 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_380
timestamp 1636043612
transform 1 0 36064 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1636043612
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1636043612
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1636043612
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1636043612
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1636043612
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1636043612
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1636043612
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1636043612
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1636043612
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output161_A
timestamp 1636043612
transform -1 0 45448 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output170_A
timestamp 1636043612
transform -1 0 44896 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1636043612
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_473
timestamp 1636043612
transform 1 0 44620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_476
timestamp 1636043612
transform 1 0 44896 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output139_A
timestamp 1636043612
transform 1 0 46920 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output142_A
timestamp 1636043612
transform -1 0 46552 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output148_A
timestamp 1636043612
transform -1 0 46000 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_482
timestamp 1636043612
transform 1 0 45448 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_488
timestamp 1636043612
transform 1 0 46000 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_494
timestamp 1636043612
transform 1 0 46552 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1636043612
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_77_505
timestamp 1636043612
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_512
timestamp 1636043612
transform 1 0 48208 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1636043612
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1636043612
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1636043612
transform 1 0 47840 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1636043612
transform -1 0 2116 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_11
timestamp 1636043612
transform 1 0 2116 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_3
timestamp 1636043612
transform 1 0 1380 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1636043612
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _175_
timestamp 1636043612
transform -1 0 3312 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__B1
timestamp 1636043612
transform 1 0 4324 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A2
timestamp 1636043612
transform -1 0 3956 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1636043612
transform 1 0 4876 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_24
timestamp 1636043612
transform 1 0 3312 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_31
timestamp 1636043612
transform 1 0 3956 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_37
timestamp 1636043612
transform 1 0 4508 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_43
timestamp 1636043612
transform 1 0 5060 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1636043612
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__B1
timestamp 1636043612
transform 1 0 6256 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__CLK
timestamp 1636043612
transform 1 0 5428 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__CLK
timestamp 1636043612
transform 1 0 6808 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_49
timestamp 1636043612
transform 1 0 5612 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_55
timestamp 1636043612
transform 1 0 6164 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_58
timestamp 1636043612
transform 1 0 6440 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_64
timestamp 1636043612
transform 1 0 6992 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__B1
timestamp 1636043612
transform 1 0 8280 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1636043612
transform 1 0 7728 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_74
timestamp 1636043612
transform 1 0 7912 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_80
timestamp 1636043612
transform 1 0 8464 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_85
timestamp 1636043612
transform 1 0 8924 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1636043612
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A
timestamp 1636043612
transform -1 0 9568 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1636043612
transform -1 0 10856 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1636043612
transform 1 0 10028 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_103
timestamp 1636043612
transform 1 0 10580 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_106
timestamp 1636043612
transform 1 0 10856 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_89
timestamp 1636043612
transform 1 0 9292 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_92
timestamp 1636043612
transform 1 0 9568 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_96
timestamp 1636043612
transform 1 0 9936 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_99
timestamp 1636043612
transform 1 0 10212 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__B1
timestamp 1636043612
transform 1 0 11224 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__A
timestamp 1636043612
transform 1 0 12512 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_112
timestamp 1636043612
transform 1 0 11408 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_120
timestamp 1636043612
transform 1 0 12144 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_126
timestamp 1636043612
transform 1 0 12696 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _375_
timestamp 1636043612
transform 1 0 11776 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_135
timestamp 1636043612
transform 1 0 13524 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_132
timestamp 1636043612
transform 1 0 13248 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__B1
timestamp 1636043612
transform 1 0 13340 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1636043612
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1636043612
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _410_
timestamp 1636043612
transform -1 0 14444 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_145
timestamp 1636043612
transform 1 0 14444 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_141
timestamp 1636043612
transform 1 0 14076 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__B1
timestamp 1636043612
transform 1 0 14812 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_151
timestamp 1636043612
transform 1 0 14996 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1636043612
transform 1 0 16100 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_155
timestamp 1636043612
transform 1 0 15364 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_159
timestamp 1636043612
transform 1 0 15732 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1636043612
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1636043612
transform -1 0 15732 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__B1
timestamp 1636043612
transform 1 0 17388 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_179
timestamp 1636043612
transform 1 0 17572 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_192
timestamp 1636043612
transform 1 0 18768 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1636043612
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _156_
timestamp 1636043612
transform 1 0 17940 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1636043612
transform 1 0 19228 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__CLK
timestamp 1636043612
transform -1 0 19964 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_199
timestamp 1636043612
transform 1 0 19412 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_205
timestamp 1636043612
transform 1 0 19964 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _460_
timestamp 1636043612
transform 1 0 20332 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1636043612
transform 1 0 22172 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_225
timestamp 1636043612
transform 1 0 21804 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_231
timestamp 1636043612
transform 1 0 22356 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_238
timestamp 1636043612
transform 1 0 23000 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _417_
timestamp 1636043612
transform -1 0 23000 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__B1
timestamp 1636043612
transform 1 0 23736 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__A
timestamp 1636043612
transform 1 0 25024 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_248
timestamp 1636043612
transform 1 0 23920 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_256
timestamp 1636043612
transform 1 0 24656 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_262
timestamp 1636043612
transform 1 0 25208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1636043612
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _418_
timestamp 1636043612
transform 1 0 24380 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A
timestamp 1636043612
transform 1 0 25576 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A
timestamp 1636043612
transform 1 0 26956 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_268
timestamp 1636043612
transform 1 0 25760 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_280
timestamp 1636043612
transform 1 0 26864 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_283
timestamp 1636043612
transform 1 0 27140 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__B1
timestamp 1636043612
transform 1 0 27692 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_291
timestamp 1636043612
transform 1 0 27876 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_304
timestamp 1636043612
transform 1 0 29072 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _141_
timestamp 1636043612
transform -1 0 29072 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__A
timestamp 1636043612
transform 1 0 29532 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_311
timestamp 1636043612
transform 1 0 29716 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_317
timestamp 1636043612
transform 1 0 30268 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1636043612
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _468_
timestamp 1636043612
transform 1 0 30360 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__B1
timestamp 1636043612
transform 1 0 32200 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_334
timestamp 1636043612
transform 1 0 31832 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_340
timestamp 1636043612
transform 1 0 32384 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _136_
timestamp 1636043612
transform 1 0 32752 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__B1
timestamp 1636043612
transform 1 0 35144 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__A
timestamp 1636043612
transform 1 0 33948 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_353
timestamp 1636043612
transform 1 0 33580 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_359
timestamp 1636043612
transform 1 0 34132 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1636043612
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_365
timestamp 1636043612
transform 1 0 34684 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_369
timestamp 1636043612
transform 1 0 35052 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1636043612
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_372
timestamp 1636043612
transform 1 0 35328 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_385
timestamp 1636043612
transform 1 0 36524 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _131_
timestamp 1636043612
transform 1 0 35696 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A
timestamp 1636043612
transform 1 0 38916 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_397
timestamp 1636043612
transform 1 0 37628 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_409
timestamp 1636043612
transform 1 0 38732 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1636043612
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1636043612
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1636043612
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1636043612
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1636043612
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_445
timestamp 1636043612
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_457
timestamp 1636043612
transform 1 0 43148 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__A
timestamp 1636043612
transform 1 0 44988 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output166_A
timestamp 1636043612
transform -1 0 44528 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output200_A
timestamp 1636043612
transform 1 0 43792 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_463
timestamp 1636043612
transform 1 0 43700 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_466
timestamp 1636043612
transform 1 0 43976 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1636043612
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_479
timestamp 1636043612
transform 1 0 45172 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1636043612
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_485
timestamp 1636043612
transform 1 0 45724 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_489
timestamp 1636043612
transform 1 0 46092 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_497
timestamp 1636043612
transform 1 0 46828 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_502
timestamp 1636043612
transform 1 0 47288 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _439_
timestamp 1636043612
transform -1 0 46092 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1636043612
transform 1 0 46920 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_510
timestamp 1636043612
transform 1 0 48024 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1636043612
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1636043612
transform 1 0 47656 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _400_
timestamp 1636043612
transform -1 0 2024 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _398_
timestamp 1636043612
transform 1 0 1932 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1636043612
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1636043612
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_5
timestamp 1636043612
transform 1 0 1564 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1636043612
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_10
timestamp 1636043612
transform 1 0 2024 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1636043612
transform -1 0 1564 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _399_
timestamp 1636043612
transform 1 0 2576 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_19
timestamp 1636043612
transform 1 0 2852 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_12
timestamp 1636043612
transform 1 0 2208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _445_
timestamp 1636043612
transform -1 0 3864 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_79_30
timestamp 1636043612
transform 1 0 3864 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_36
timestamp 1636043612
transform 1 0 4416 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1636043612
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_32
timestamp 1636043612
transform 1 0 4048 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1636043612
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _174_
timestamp 1636043612
transform 1 0 4508 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _401_
timestamp 1636043612
transform 1 0 3772 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _446_
timestamp 1636043612
transform 1 0 4416 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A
timestamp 1636043612
transform 1 0 5704 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_46
timestamp 1636043612
transform 1 0 5336 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_52
timestamp 1636043612
transform 1 0 5888 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_57
timestamp 1636043612
transform 1 0 6348 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_52
timestamp 1636043612
transform 1 0 5888 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_56
timestamp 1636043612
transform 1 0 6256 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1636043612
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _172_
timestamp 1636043612
transform -1 0 7268 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _448_
timestamp 1636043612
transform 1 0 6348 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _405_
timestamp 1636043612
transform -1 0 8096 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_73
timestamp 1636043612
transform 1 0 7820 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_76
timestamp 1636043612
transform 1 0 8096 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_67
timestamp 1636043612
transform 1 0 7268 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _404_
timestamp 1636043612
transform 1 0 8188 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _169_
timestamp 1636043612
transform 1 0 8556 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1636043612
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_80
timestamp 1636043612
transform 1 0 8464 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_80
timestamp 1636043612
transform 1 0 8464 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _450_
timestamp 1636043612
transform 1 0 8924 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_79_104
timestamp 1636043612
transform 1 0 10672 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_90
timestamp 1636043612
transform 1 0 9384 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_97
timestamp 1636043612
transform 1 0 10028 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_101
timestamp 1636043612
transform 1 0 10396 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_107
timestamp 1636043612
transform 1 0 10948 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _406_
timestamp 1636043612
transform 1 0 9752 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _407_
timestamp 1636043612
transform -1 0 10672 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _452_
timestamp 1636043612
transform 1 0 11040 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_79_122
timestamp 1636043612
transform 1 0 12328 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_131
timestamp 1636043612
transform 1 0 13156 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_124
timestamp 1636043612
transform 1 0 12512 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_131
timestamp 1636043612
transform 1 0 13156 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1636043612
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _165_
timestamp 1636043612
transform -1 0 12328 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _408_
timestamp 1636043612
transform 1 0 12880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp 1636043612
transform -1 0 13156 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_144
timestamp 1636043612
transform 1 0 14352 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_148
timestamp 1636043612
transform 1 0 14720 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1636043612
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1636043612
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _161_
timestamp 1636043612
transform 1 0 14812 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _163_
timestamp 1636043612
transform 1 0 13524 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _454_
timestamp 1636043612
transform 1 0 14076 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1636043612
transform 1 0 16652 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A
timestamp 1636043612
transform 1 0 16008 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_158
timestamp 1636043612
transform 1 0 15640 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_164
timestamp 1636043612
transform 1 0 16192 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_171
timestamp 1636043612
transform 1 0 16836 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_157
timestamp 1636043612
transform 1 0 15548 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1636043612
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _455_
timestamp 1636043612
transform -1 0 17388 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _412_
timestamp 1636043612
transform 1 0 17756 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _379_
timestamp 1636043612
transform 1 0 17204 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_184
timestamp 1636043612
transform 1 0 18032 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_177
timestamp 1636043612
transform 1 0 17388 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_179
timestamp 1636043612
transform 1 0 17572 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _413_
timestamp 1636043612
transform 1 0 18400 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1636043612
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1636043612
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_191
timestamp 1636043612
transform 1 0 18676 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _458_
timestamp 1636043612
transform 1 0 18308 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  _382_
timestamp 1636043612
transform 1 0 19596 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_205
timestamp 1636043612
transform 1 0 19964 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_197
timestamp 1636043612
transform 1 0 19228 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_203
timestamp 1636043612
transform 1 0 19780 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _415_
timestamp 1636043612
transform -1 0 20608 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_212
timestamp 1636043612
transform 1 0 20608 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_209
timestamp 1636043612
transform 1 0 20332 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A
timestamp 1636043612
transform 1 0 20700 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1636043612
transform -1 0 20332 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_218
timestamp 1636043612
transform 1 0 21160 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_215
timestamp 1636043612
transform 1 0 20884 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A
timestamp 1636043612
transform 1 0 20976 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__B1
timestamp 1636043612
transform 1 0 22172 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1636043612
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_225
timestamp 1636043612
transform 1 0 21804 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_231
timestamp 1636043612
transform 1 0 22356 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_225
timestamp 1636043612
transform 1 0 21804 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1636043612
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _150_
timestamp 1636043612
transform -1 0 23552 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _416_
timestamp 1636043612
transform -1 0 21804 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _461_
timestamp 1636043612
transform 1 0 22356 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_79_244
timestamp 1636043612
transform 1 0 23552 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_261
timestamp 1636043612
transform 1 0 25116 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_247
timestamp 1636043612
transform 1 0 23828 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1636043612
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_253
timestamp 1636043612
transform 1 0 24380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_257
timestamp 1636043612
transform 1 0 24748 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1636043612
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _148_
timestamp 1636043612
transform 1 0 24288 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _463_
timestamp 1636043612
transform 1 0 24840 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _419_
timestamp 1636043612
transform -1 0 25760 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_268
timestamp 1636043612
transform 1 0 25760 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _420_
timestamp 1636043612
transform -1 0 26956 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_274
timestamp 1636043612
transform 1 0 26312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_274
timestamp 1636043612
transform 1 0 26312 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1636043612
transform 1 0 26128 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1636043612
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_281
timestamp 1636043612
transform 1 0 26956 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_281
timestamp 1636043612
transform 1 0 26956 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__A
timestamp 1636043612
transform 1 0 27140 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_285
timestamp 1636043612
transform 1 0 27324 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_293
timestamp 1636043612
transform 1 0 28060 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_289
timestamp 1636043612
transform 1 0 27692 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_293
timestamp 1636043612
transform 1 0 28060 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_297
timestamp 1636043612
transform 1 0 28428 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_302
timestamp 1636043612
transform 1 0 28888 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _421_
timestamp 1636043612
transform -1 0 28060 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _467_
timestamp 1636043612
transform 1 0 28152 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1636043612
transform 1 0 28520 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _422_
timestamp 1636043612
transform 1 0 29532 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1636043612
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_312
timestamp 1636043612
transform 1 0 29808 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_79_310
timestamp 1636043612
transform 1 0 29624 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1636043612
transform 1 0 31004 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _423_
timestamp 1636043612
transform -1 0 30636 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _139_
timestamp 1636043612
transform 1 0 30820 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_80_321
timestamp 1636043612
transform 1 0 30636 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_319
timestamp 1636043612
transform 1 0 30452 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_316
timestamp 1636043612
transform 1 0 30176 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__B1
timestamp 1636043612
transform 1 0 30268 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1636043612
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_333
timestamp 1636043612
transform 1 0 31740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_329
timestamp 1636043612
transform 1 0 31372 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_332
timestamp 1636043612
transform 1 0 31648 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A
timestamp 1636043612
transform 1 0 32108 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_345
timestamp 1636043612
transform 1 0 32844 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_339
timestamp 1636043612
transform 1 0 32292 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1636043612
transform 1 0 32660 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _470_
timestamp 1636043612
transform 1 0 33212 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _469_
timestamp 1636043612
transform 1 0 31832 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1636043612
transform 1 0 34776 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A
timestamp 1636043612
transform 1 0 33672 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_365
timestamp 1636043612
transform 1 0 34684 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_371
timestamp 1636043612
transform 1 0 35236 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_350
timestamp 1636043612
transform 1 0 33304 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_356
timestamp 1636043612
transform 1 0 33856 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_365
timestamp 1636043612
transform 1 0 34684 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_368
timestamp 1636043612
transform 1 0 34960 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1636043612
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _427_
timestamp 1636043612
transform -1 0 35604 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _130_
timestamp 1636043612
transform 1 0 35880 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_80_375
timestamp 1636043612
transform 1 0 35604 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_374
timestamp 1636043612
transform 1 0 35512 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__B1
timestamp 1636043612
transform 1 0 35328 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1636043612
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1636043612
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_387
timestamp 1636043612
transform 1 0 36708 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _473_
timestamp 1636043612
transform 1 0 37260 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _472_
timestamp 1636043612
transform 1 0 35972 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A
timestamp 1636043612
transform 1 0 37812 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A
timestamp 1636043612
transform 1 0 38364 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__A
timestamp 1636043612
transform 1 0 39100 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_409
timestamp 1636043612
transform 1 0 38732 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_395
timestamp 1636043612
transform 1 0 37444 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_401
timestamp 1636043612
transform 1 0 37996 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_407
timestamp 1636043612
transform 1 0 38548 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _430_
timestamp 1636043612
transform -1 0 39376 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _397_
timestamp 1636043612
transform -1 0 40112 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1636043612
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_424
timestamp 1636043612
transform 1 0 40112 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_416
timestamp 1636043612
transform 1 0 39376 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_415
timestamp 1636043612
transform 1 0 39284 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1636043612
transform 1 0 39652 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _435_
timestamp 1636043612
transform -1 0 41032 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_80_434
timestamp 1636043612
transform 1 0 41032 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_430
timestamp 1636043612
transform 1 0 40664 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1636043612
transform 1 0 40940 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_435
timestamp 1636043612
transform 1 0 41124 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_421
timestamp 1636043612
transform 1 0 39836 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _432_
timestamp 1636043612
transform -1 0 41952 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_440
timestamp 1636043612
transform 1 0 41584 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _436_
timestamp 1636043612
transform 1 0 42412 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1636043612
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_450
timestamp 1636043612
transform 1 0 42504 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_444
timestamp 1636043612
transform 1 0 41952 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1636043612
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A
timestamp 1636043612
transform 1 0 42320 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _433_
timestamp 1636043612
transform -1 0 43148 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_457
timestamp 1636043612
transform 1 0 43148 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_452
timestamp 1636043612
transform 1 0 42688 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _437_
timestamp 1636043612
transform -1 0 43516 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_463
timestamp 1636043612
transform 1 0 43700 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_461
timestamp 1636043612
transform 1 0 43516 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A
timestamp 1636043612
transform 1 0 43884 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A
timestamp 1636043612
transform 1 0 43516 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _438_
timestamp 1636043612
transform -1 0 44712 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _434_
timestamp 1636043612
transform -1 0 44344 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_80_470
timestamp 1636043612
transform 1 0 44344 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_467
timestamp 1636043612
transform 1 0 44068 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _393_
timestamp 1636043612
transform -1 0 45356 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _235_
timestamp 1636043612
transform 1 0 44988 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1636043612
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_474
timestamp 1636043612
transform 1 0 44712 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_480
timestamp 1636043612
transform 1 0 45264 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1636043612
transform 1 0 45632 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_487
timestamp 1636043612
transform 1 0 45908 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_481
timestamp 1636043612
transform 1 0 45356 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1636043612
transform 1 0 46000 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1636043612
transform 1 0 46368 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_488
timestamp 1636043612
transform 1 0 46000 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_492
timestamp 1636043612
transform 1 0 46368 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1636043612
transform 1 0 46736 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1636043612
transform 1 0 47104 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_496
timestamp 1636043612
transform 1 0 46736 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_500
timestamp 1636043612
transform 1 0 47104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_505
timestamp 1636043612
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_512
timestamp 1636043612
transform 1 0 48208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_504
timestamp 1636043612
transform 1 0 47472 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1636043612
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1636043612
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1636043612
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1636043612
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1636043612
transform 1 0 47840 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1636043612
transform 1 0 47840 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_17
timestamp 1636043612
transform 1 0 2668 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_81_7
timestamp 1636043612
transform 1 0 1748 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1636043612
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1636043612
transform -1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1636043612
transform -1 0 2668 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_29
timestamp 1636043612
transform 1 0 3772 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_37
timestamp 1636043612
transform 1 0 4508 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _369_
timestamp 1636043612
transform 1 0 3404 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _402_
timestamp 1636043612
transform 1 0 4876 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1636043612
transform 1 0 4140 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_44
timestamp 1636043612
transform 1 0 5152 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1636043612
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1636043612
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_61
timestamp 1636043612
transform 1 0 6716 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1636043612
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _403_
timestamp 1636043612
transform -1 0 5796 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1636043612
transform 1 0 6348 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__A
timestamp 1636043612
transform 1 0 8004 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_71
timestamp 1636043612
transform 1 0 7636 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_77
timestamp 1636043612
transform 1 0 8188 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_85
timestamp 1636043612
transform 1 0 8924 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1636043612
transform -1 0 7636 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1636043612
transform 1 0 8556 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1636043612
transform 1 0 9292 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_103
timestamp 1636043612
transform 1 0 10580 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1636043612
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_91
timestamp 1636043612
transform 1 0 9476 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_99
timestamp 1636043612
transform 1 0 10212 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1636043612
transform -1 0 10212 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1636043612
transform -1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A
timestamp 1636043612
transform 1 0 11500 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_115
timestamp 1636043612
transform 1 0 11684 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_123
timestamp 1636043612
transform 1 0 12420 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_131
timestamp 1636043612
transform 1 0 13156 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1636043612
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _376_
timestamp 1636043612
transform 1 0 12052 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1636043612
transform 1 0 12788 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1636043612
transform 1 0 14260 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_139
timestamp 1636043612
transform 1 0 13892 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_145
timestamp 1636043612
transform 1 0 14444 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1636043612
transform -1 0 13892 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1636043612
transform -1 0 15180 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1636043612
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_153
timestamp 1636043612
transform 1 0 15180 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_159
timestamp 1636043612
transform 1 0 15732 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_164
timestamp 1636043612
transform 1 0 16192 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_171
timestamp 1636043612
transform 1 0 16836 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1636043612
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1636043612
transform -1 0 16192 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_179
timestamp 1636043612
transform 1 0 17572 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_187
timestamp 1636043612
transform 1 0 18308 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_195
timestamp 1636043612
transform 1 0 19044 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _378_
timestamp 1636043612
transform 1 0 17204 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1636043612
transform 1 0 17940 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1636043612
transform 1 0 18676 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A
timestamp 1636043612
transform 1 0 21160 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_207
timestamp 1636043612
transform 1 0 20148 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_214
timestamp 1636043612
transform 1 0 20792 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _414_
timestamp 1636043612
transform 1 0 20516 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1636043612
transform 1 0 19780 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1636043612
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_229
timestamp 1636043612
transform 1 0 22172 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_237
timestamp 1636043612
transform 1 0 22908 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1636043612
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1636043612
transform 1 0 21804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1636043612
transform 1 0 22540 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_241
timestamp 1636043612
transform 1 0 23276 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_246
timestamp 1636043612
transform 1 0 23736 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_254
timestamp 1636043612
transform 1 0 24472 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_262
timestamp 1636043612
transform 1 0 25208 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _385_
timestamp 1636043612
transform 1 0 23368 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1636043612
transform 1 0 24104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1636043612
transform 1 0 24840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_270
timestamp 1636043612
transform 1 0 25944 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_275
timestamp 1636043612
transform 1 0 26404 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1636043612
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_281
timestamp 1636043612
transform 1 0 26956 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1636043612
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1636043612
transform -1 0 26404 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_289
timestamp 1636043612
transform 1 0 27692 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_297
timestamp 1636043612
transform 1 0 28428 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_305
timestamp 1636043612
transform 1 0 29164 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _387_
timestamp 1636043612
transform 1 0 27324 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _391_
timestamp 1636043612
transform 1 0 28796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1636043612
transform 1 0 28060 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_311
timestamp 1636043612
transform 1 0 29716 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_316
timestamp 1636043612
transform 1 0 30176 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_324
timestamp 1636043612
transform 1 0 30912 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _392_
timestamp 1636043612
transform 1 0 31004 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1636043612
transform 1 0 29808 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1636043612
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1636043612
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_337
timestamp 1636043612
transform 1 0 32108 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_343
timestamp 1636043612
transform 1 0 32660 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1636043612
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _424_
timestamp 1636043612
transform 1 0 33028 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1636043612
transform 1 0 32292 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_350
timestamp 1636043612
transform 1 0 33304 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_357
timestamp 1636043612
transform 1 0 33948 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_364
timestamp 1636043612
transform 1 0 34592 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _394_
timestamp 1636043612
transform 1 0 34960 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _425_
timestamp 1636043612
transform 1 0 33672 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _426_
timestamp 1636043612
transform -1 0 34592 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_372
timestamp 1636043612
transform 1 0 35328 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_81_384
timestamp 1636043612
transform 1 0 36432 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1636043612
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1636043612
transform -1 0 36432 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1636043612
transform 1 0 37260 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_397
timestamp 1636043612
transform 1 0 37628 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_404
timestamp 1636043612
transform 1 0 38272 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_411
timestamp 1636043612
transform 1 0 38916 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _428_
timestamp 1636043612
transform 1 0 37996 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _429_
timestamp 1636043612
transform 1 0 38640 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_81_419
timestamp 1636043612
transform 1 0 39652 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_424
timestamp 1636043612
transform 1 0 40112 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_431
timestamp 1636043612
transform 1 0 40756 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _396_
timestamp 1636043612
transform -1 0 40756 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _431_
timestamp 1636043612
transform 1 0 41124 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1636043612
transform 1 0 39744 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1636043612
transform -1 0 41952 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_438
timestamp 1636043612
transform 1 0 41400 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1636043612
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_453
timestamp 1636043612
transform 1 0 42780 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1636043612
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1636043612
transform 1 0 42412 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_465
timestamp 1636043612
transform 1 0 43884 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_471
timestamp 1636043612
transform 1 0 44436 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_476
timestamp 1636043612
transform 1 0 44896 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1636043612
transform 1 0 45264 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1636043612
transform 1 0 43516 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1636043612
transform 1 0 44528 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_484
timestamp 1636043612
transform 1 0 45632 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_492
timestamp 1636043612
transform 1 0 46368 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1636043612
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1636043612
transform 1 0 46736 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1636043612
transform 1 0 46000 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1636043612
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1636043612
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1636043612
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1636043612
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1636043612
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_15
timestamp 1636043612
transform 1 0 2484 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_7
timestamp 1636043612
transform 1 0 1748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1636043612
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1636043612
transform -1 0 1748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1636043612
transform 1 0 2116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1636043612
transform 1 0 2852 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_23
timestamp 1636043612
transform 1 0 3220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1636043612
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_33
timestamp 1636043612
transform 1 0 4140 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_41
timestamp 1636043612
transform 1 0 4876 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1636043612
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1636043612
transform 1 0 3772 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1636043612
transform -1 0 4876 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_49
timestamp 1636043612
transform 1 0 5612 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_55
timestamp 1636043612
transform 1 0 6164 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_61
timestamp 1636043612
transform 1 0 6716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1636043612
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1636043612
transform 1 0 6348 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1636043612
transform -1 0 7452 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1636043612
transform -1 0 5612 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_69
timestamp 1636043612
transform 1 0 7452 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_75
timestamp 1636043612
transform 1 0 8004 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_80
timestamp 1636043612
transform 1 0 8464 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1636043612
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1636043612
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1636043612
transform 1 0 8096 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__CLK
timestamp 1636043612
transform -1 0 10304 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_100
timestamp 1636043612
transform 1 0 10304 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_108
timestamp 1636043612
transform 1 0 11040 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_89
timestamp 1636043612
transform 1 0 9292 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_94
timestamp 1636043612
transform 1 0 9752 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1636043612
transform -1 0 9752 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1636043612
transform 1 0 10672 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__CLK
timestamp 1636043612
transform -1 0 12788 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_113
timestamp 1636043612
transform 1 0 11500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_121
timestamp 1636043612
transform 1 0 12236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_127
timestamp 1636043612
transform 1 0 12788 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1636043612
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1636043612
transform 1 0 13156 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1636043612
transform -1 0 12236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__CLK
timestamp 1636043612
transform -1 0 15272 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1636043612
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1636043612
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_141
timestamp 1636043612
transform 1 0 14076 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_148
timestamp 1636043612
transform 1 0 14720 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1636043612
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1636043612
transform 1 0 14352 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_154
timestamp 1636043612
transform 1 0 15272 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_162
timestamp 1636043612
transform 1 0 16008 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_82_169
timestamp 1636043612
transform 1 0 16652 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1636043612
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1636043612
transform 1 0 15640 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1636043612
transform -1 0 17296 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_176
timestamp 1636043612
transform 1 0 17296 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_184
timestamp 1636043612
transform 1 0 18032 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1636043612
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1636043612
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1636043612
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1636043612
transform -1 0 18492 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_197
timestamp 1636043612
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_203
timestamp 1636043612
transform 1 0 19780 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_211
timestamp 1636043612
transform 1 0 20516 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_216
timestamp 1636043612
transform 1 0 20976 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1636043612
transform -1 0 19780 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1636043612
transform 1 0 20608 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_225
timestamp 1636043612
transform 1 0 21804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_230
timestamp 1636043612
transform 1 0 22264 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_238
timestamp 1636043612
transform 1 0 23000 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1636043612
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1636043612
transform 1 0 21896 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1636043612
transform 1 0 23092 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_243
timestamp 1636043612
transform 1 0 23460 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1636043612
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_257
timestamp 1636043612
transform 1 0 24748 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1636043612
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1636043612
transform 1 0 24380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_265
timestamp 1636043612
transform 1 0 25484 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_271
timestamp 1636043612
transform 1 0 26036 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_279
timestamp 1636043612
transform 1 0 26772 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1636043612
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1636043612
transform 1 0 25668 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1636043612
transform 1 0 26956 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A
timestamp 1636043612
transform -1 0 29072 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_285
timestamp 1636043612
transform 1 0 27324 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_293
timestamp 1636043612
transform 1 0 28060 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_298
timestamp 1636043612
transform 1 0 28520 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_304
timestamp 1636043612
transform 1 0 29072 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1636043612
transform 1 0 28152 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_313
timestamp 1636043612
transform 1 0 29900 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_325
timestamp 1636043612
transform 1 0 31004 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1636043612
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1636043612
transform 1 0 29532 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1636043612
transform 1 0 30636 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__A
timestamp 1636043612
transform -1 0 31556 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_331
timestamp 1636043612
transform 1 0 31556 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_335
timestamp 1636043612
transform 1 0 31924 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_341
timestamp 1636043612
transform 1 0 32476 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_347
timestamp 1636043612
transform 1 0 33028 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1636043612
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1636043612
transform -1 0 32476 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1636043612
transform -1 0 33488 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_352
timestamp 1636043612
transform 1 0 33488 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_360
timestamp 1636043612
transform 1 0 34224 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_369
timestamp 1636043612
transform 1 0 35052 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1636043612
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1636043612
transform 1 0 34684 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1636043612
transform 1 0 33856 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_379
timestamp 1636043612
transform 1 0 35972 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_387
timestamp 1636043612
transform 1 0 36708 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_391
timestamp 1636043612
transform 1 0 37076 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1636043612
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1636043612
transform 1 0 35604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1636043612
transform -1 0 37628 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1636043612
transform 1 0 36340 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_397
timestamp 1636043612
transform 1 0 37628 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_401
timestamp 1636043612
transform 1 0 37996 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_406
timestamp 1636043612
transform 1 0 38456 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_414
timestamp 1636043612
transform 1 0 39192 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1636043612
transform -1 0 38456 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1636043612
transform 1 0 38824 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_425
timestamp 1636043612
transform 1 0 40204 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_433
timestamp 1636043612
transform 1 0 40940 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1636043612
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1636043612
transform 1 0 39836 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1636043612
transform -1 0 40940 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_441
timestamp 1636043612
transform 1 0 41676 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_447
timestamp 1636043612
transform 1 0 42228 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_453
timestamp 1636043612
transform 1 0 42780 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1636043612
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1636043612
transform 1 0 42412 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1636043612
transform 1 0 43148 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1636043612
transform 1 0 41308 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_461
timestamp 1636043612
transform 1 0 43516 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_467
timestamp 1636043612
transform 1 0 44068 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1636043612
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_477
timestamp 1636043612
transform 1 0 44988 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1636043612
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1636043612
transform 1 0 45264 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1636043612
transform 1 0 44160 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_484
timestamp 1636043612
transform 1 0 45632 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_492
timestamp 1636043612
transform 1 0 46368 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1636043612
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1636043612
transform 1 0 46736 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1636043612
transform 1 0 46000 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_505
timestamp 1636043612
transform 1 0 47564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_512
timestamp 1636043612
transform 1 0 48208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1636043612
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1636043612
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1636043612
transform 1 0 47840 0 1 46784
box -38 -48 406 592
<< labels >>
rlabel metal3 s 49200 41760 50000 41880 6 csb0
port 0 nsew signal tristate
rlabel metal3 s 49200 43120 50000 43240 6 csb1
port 1 nsew signal tristate
rlabel metal3 s 49200 43800 50000 43920 6 din0[0]
port 2 nsew signal tristate
rlabel metal2 s 49238 0 49294 800 6 din0[10]
port 3 nsew signal tristate
rlabel metal2 s 48410 49200 48466 50000 6 din0[11]
port 4 nsew signal tristate
rlabel metal3 s 49200 45704 50000 45824 6 din0[12]
port 5 nsew signal tristate
rlabel metal3 s 0 30472 800 30592 6 din0[13]
port 6 nsew signal tristate
rlabel metal2 s 49330 0 49386 800 6 din0[14]
port 7 nsew signal tristate
rlabel metal3 s 49200 46384 50000 46504 6 din0[15]
port 8 nsew signal tristate
rlabel metal2 s 49422 0 49478 800 6 din0[16]
port 9 nsew signal tristate
rlabel metal2 s 49514 0 49570 800 6 din0[17]
port 10 nsew signal tristate
rlabel metal3 s 49200 47064 50000 47184 6 din0[18]
port 11 nsew signal tristate
rlabel metal2 s 49606 0 49662 800 6 din0[19]
port 12 nsew signal tristate
rlabel metal3 s 0 2728 800 2848 6 din0[1]
port 13 nsew signal tristate
rlabel metal2 s 48870 49200 48926 50000 6 din0[20]
port 14 nsew signal tristate
rlabel metal3 s 0 36048 800 36168 6 din0[21]
port 15 nsew signal tristate
rlabel metal3 s 0 41624 800 41744 6 din0[22]
port 16 nsew signal tristate
rlabel metal2 s 49698 0 49754 800 6 din0[23]
port 17 nsew signal tristate
rlabel metal2 s 49238 49200 49294 50000 6 din0[24]
port 18 nsew signal tristate
rlabel metal2 s 49698 49200 49754 50000 6 din0[25]
port 19 nsew signal tristate
rlabel metal3 s 49200 47608 50000 47728 6 din0[26]
port 20 nsew signal tristate
rlabel metal3 s 49200 48288 50000 48408 6 din0[27]
port 21 nsew signal tristate
rlabel metal2 s 49790 0 49846 800 6 din0[28]
port 22 nsew signal tristate
rlabel metal3 s 49200 48968 50000 49088 6 din0[29]
port 23 nsew signal tristate
rlabel metal2 s 47582 49200 47638 50000 6 din0[2]
port 24 nsew signal tristate
rlabel metal3 s 49200 49648 50000 49768 6 din0[30]
port 25 nsew signal tristate
rlabel metal3 s 0 47200 800 47320 6 din0[31]
port 26 nsew signal tristate
rlabel metal3 s 0 8168 800 8288 6 din0[3]
port 27 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 din0[4]
port 28 nsew signal tristate
rlabel metal3 s 49200 44344 50000 44464 6 din0[5]
port 29 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 din0[6]
port 30 nsew signal tristate
rlabel metal3 s 0 24896 800 25016 6 din0[7]
port 31 nsew signal tristate
rlabel metal3 s 49200 45024 50000 45144 6 din0[8]
port 32 nsew signal tristate
rlabel metal2 s 48042 49200 48098 50000 6 din0[9]
port 33 nsew signal tristate
rlabel metal3 s 49200 280 50000 400 6 dout0[0]
port 34 nsew signal input
rlabel metal3 s 49200 6672 50000 6792 6 dout0[10]
port 35 nsew signal input
rlabel metal3 s 49200 7352 50000 7472 6 dout0[11]
port 36 nsew signal input
rlabel metal3 s 49200 8032 50000 8152 6 dout0[12]
port 37 nsew signal input
rlabel metal3 s 49200 8712 50000 8832 6 dout0[13]
port 38 nsew signal input
rlabel metal3 s 49200 9256 50000 9376 6 dout0[14]
port 39 nsew signal input
rlabel metal3 s 49200 9936 50000 10056 6 dout0[15]
port 40 nsew signal input
rlabel metal3 s 49200 10616 50000 10736 6 dout0[16]
port 41 nsew signal input
rlabel metal3 s 49200 11296 50000 11416 6 dout0[17]
port 42 nsew signal input
rlabel metal3 s 49200 11976 50000 12096 6 dout0[18]
port 43 nsew signal input
rlabel metal3 s 49200 12520 50000 12640 6 dout0[19]
port 44 nsew signal input
rlabel metal3 s 49200 824 50000 944 6 dout0[1]
port 45 nsew signal input
rlabel metal3 s 49200 13200 50000 13320 6 dout0[20]
port 46 nsew signal input
rlabel metal3 s 49200 13880 50000 14000 6 dout0[21]
port 47 nsew signal input
rlabel metal3 s 49200 14560 50000 14680 6 dout0[22]
port 48 nsew signal input
rlabel metal3 s 49200 15104 50000 15224 6 dout0[23]
port 49 nsew signal input
rlabel metal3 s 49200 15784 50000 15904 6 dout0[24]
port 50 nsew signal input
rlabel metal3 s 49200 16464 50000 16584 6 dout0[25]
port 51 nsew signal input
rlabel metal3 s 49200 17144 50000 17264 6 dout0[26]
port 52 nsew signal input
rlabel metal3 s 49200 17824 50000 17944 6 dout0[27]
port 53 nsew signal input
rlabel metal3 s 49200 18368 50000 18488 6 dout0[28]
port 54 nsew signal input
rlabel metal3 s 49200 19048 50000 19168 6 dout0[29]
port 55 nsew signal input
rlabel metal3 s 49200 1504 50000 1624 6 dout0[2]
port 56 nsew signal input
rlabel metal3 s 49200 19728 50000 19848 6 dout0[30]
port 57 nsew signal input
rlabel metal3 s 49200 20408 50000 20528 6 dout0[31]
port 58 nsew signal input
rlabel metal3 s 49200 2184 50000 2304 6 dout0[3]
port 59 nsew signal input
rlabel metal3 s 49200 2864 50000 2984 6 dout0[4]
port 60 nsew signal input
rlabel metal3 s 49200 3408 50000 3528 6 dout0[5]
port 61 nsew signal input
rlabel metal3 s 49200 4088 50000 4208 6 dout0[6]
port 62 nsew signal input
rlabel metal3 s 49200 4768 50000 4888 6 dout0[7]
port 63 nsew signal input
rlabel metal3 s 49200 5448 50000 5568 6 dout0[8]
port 64 nsew signal input
rlabel metal3 s 49200 6128 50000 6248 6 dout0[9]
port 65 nsew signal input
rlabel metal3 s 49200 20952 50000 21072 6 dout1[0]
port 66 nsew signal input
rlabel metal3 s 49200 27480 50000 27600 6 dout1[10]
port 67 nsew signal input
rlabel metal3 s 49200 28160 50000 28280 6 dout1[11]
port 68 nsew signal input
rlabel metal3 s 49200 28840 50000 28960 6 dout1[12]
port 69 nsew signal input
rlabel metal3 s 49200 29520 50000 29640 6 dout1[13]
port 70 nsew signal input
rlabel metal3 s 49200 30064 50000 30184 6 dout1[14]
port 71 nsew signal input
rlabel metal3 s 49200 30744 50000 30864 6 dout1[15]
port 72 nsew signal input
rlabel metal3 s 49200 31424 50000 31544 6 dout1[16]
port 73 nsew signal input
rlabel metal3 s 49200 32104 50000 32224 6 dout1[17]
port 74 nsew signal input
rlabel metal3 s 49200 32648 50000 32768 6 dout1[18]
port 75 nsew signal input
rlabel metal3 s 49200 33328 50000 33448 6 dout1[19]
port 76 nsew signal input
rlabel metal3 s 49200 21632 50000 21752 6 dout1[1]
port 77 nsew signal input
rlabel metal3 s 49200 34008 50000 34128 6 dout1[20]
port 78 nsew signal input
rlabel metal3 s 49200 34688 50000 34808 6 dout1[21]
port 79 nsew signal input
rlabel metal3 s 49200 35368 50000 35488 6 dout1[22]
port 80 nsew signal input
rlabel metal3 s 49200 35912 50000 36032 6 dout1[23]
port 81 nsew signal input
rlabel metal3 s 49200 36592 50000 36712 6 dout1[24]
port 82 nsew signal input
rlabel metal3 s 49200 37272 50000 37392 6 dout1[25]
port 83 nsew signal input
rlabel metal3 s 49200 37952 50000 38072 6 dout1[26]
port 84 nsew signal input
rlabel metal3 s 49200 38496 50000 38616 6 dout1[27]
port 85 nsew signal input
rlabel metal3 s 49200 39176 50000 39296 6 dout1[28]
port 86 nsew signal input
rlabel metal3 s 49200 39856 50000 39976 6 dout1[29]
port 87 nsew signal input
rlabel metal3 s 49200 22312 50000 22432 6 dout1[2]
port 88 nsew signal input
rlabel metal3 s 49200 40536 50000 40656 6 dout1[30]
port 89 nsew signal input
rlabel metal3 s 49200 41216 50000 41336 6 dout1[31]
port 90 nsew signal input
rlabel metal3 s 49200 22992 50000 23112 6 dout1[3]
port 91 nsew signal input
rlabel metal3 s 49200 23672 50000 23792 6 dout1[4]
port 92 nsew signal input
rlabel metal3 s 49200 24216 50000 24336 6 dout1[5]
port 93 nsew signal input
rlabel metal3 s 49200 24896 50000 25016 6 dout1[6]
port 94 nsew signal input
rlabel metal3 s 49200 25576 50000 25696 6 dout1[7]
port 95 nsew signal input
rlabel metal3 s 49200 26256 50000 26376 6 dout1[8]
port 96 nsew signal input
rlabel metal3 s 49200 26800 50000 26920 6 dout1[9]
port 97 nsew signal input
rlabel metal2 s 202 49200 258 50000 6 io_in[0]
port 98 nsew signal input
rlabel metal2 s 12622 49200 12678 50000 6 io_in[10]
port 99 nsew signal input
rlabel metal2 s 13910 49200 13966 50000 6 io_in[11]
port 100 nsew signal input
rlabel metal2 s 15106 49200 15162 50000 6 io_in[12]
port 101 nsew signal input
rlabel metal2 s 16394 49200 16450 50000 6 io_in[13]
port 102 nsew signal input
rlabel metal2 s 17682 49200 17738 50000 6 io_in[14]
port 103 nsew signal input
rlabel metal2 s 18878 49200 18934 50000 6 io_in[15]
port 104 nsew signal input
rlabel metal2 s 20166 49200 20222 50000 6 io_in[16]
port 105 nsew signal input
rlabel metal2 s 21362 49200 21418 50000 6 io_in[17]
port 106 nsew signal input
rlabel metal2 s 22650 49200 22706 50000 6 io_in[18]
port 107 nsew signal input
rlabel metal2 s 23846 49200 23902 50000 6 io_in[19]
port 108 nsew signal input
rlabel metal2 s 1398 49200 1454 50000 6 io_in[1]
port 109 nsew signal input
rlabel metal2 s 25134 49200 25190 50000 6 io_in[20]
port 110 nsew signal input
rlabel metal2 s 26422 49200 26478 50000 6 io_in[21]
port 111 nsew signal input
rlabel metal2 s 27618 49200 27674 50000 6 io_in[22]
port 112 nsew signal input
rlabel metal2 s 28906 49200 28962 50000 6 io_in[23]
port 113 nsew signal input
rlabel metal2 s 30102 49200 30158 50000 6 io_in[24]
port 114 nsew signal input
rlabel metal2 s 31390 49200 31446 50000 6 io_in[25]
port 115 nsew signal input
rlabel metal2 s 32586 49200 32642 50000 6 io_in[26]
port 116 nsew signal input
rlabel metal2 s 33874 49200 33930 50000 6 io_in[27]
port 117 nsew signal input
rlabel metal2 s 35162 49200 35218 50000 6 io_in[28]
port 118 nsew signal input
rlabel metal2 s 36358 49200 36414 50000 6 io_in[29]
port 119 nsew signal input
rlabel metal2 s 2686 49200 2742 50000 6 io_in[2]
port 120 nsew signal input
rlabel metal2 s 37646 49200 37702 50000 6 io_in[30]
port 121 nsew signal input
rlabel metal2 s 38842 49200 38898 50000 6 io_in[31]
port 122 nsew signal input
rlabel metal2 s 40130 49200 40186 50000 6 io_in[32]
port 123 nsew signal input
rlabel metal2 s 41326 49200 41382 50000 6 io_in[33]
port 124 nsew signal input
rlabel metal2 s 42614 49200 42670 50000 6 io_in[34]
port 125 nsew signal input
rlabel metal2 s 43902 49200 43958 50000 6 io_in[35]
port 126 nsew signal input
rlabel metal2 s 45098 49200 45154 50000 6 io_in[36]
port 127 nsew signal input
rlabel metal2 s 46386 49200 46442 50000 6 io_in[37]
port 128 nsew signal input
rlabel metal2 s 3882 49200 3938 50000 6 io_in[3]
port 129 nsew signal input
rlabel metal2 s 5170 49200 5226 50000 6 io_in[4]
port 130 nsew signal input
rlabel metal2 s 6366 49200 6422 50000 6 io_in[5]
port 131 nsew signal input
rlabel metal2 s 7654 49200 7710 50000 6 io_in[6]
port 132 nsew signal input
rlabel metal2 s 8942 49200 8998 50000 6 io_in[7]
port 133 nsew signal input
rlabel metal2 s 10138 49200 10194 50000 6 io_in[8]
port 134 nsew signal input
rlabel metal2 s 11426 49200 11482 50000 6 io_in[9]
port 135 nsew signal input
rlabel metal2 s 570 49200 626 50000 6 io_oeb[0]
port 136 nsew signal tristate
rlabel metal2 s 13082 49200 13138 50000 6 io_oeb[10]
port 137 nsew signal tristate
rlabel metal2 s 14278 49200 14334 50000 6 io_oeb[11]
port 138 nsew signal tristate
rlabel metal2 s 15566 49200 15622 50000 6 io_oeb[12]
port 139 nsew signal tristate
rlabel metal2 s 16854 49200 16910 50000 6 io_oeb[13]
port 140 nsew signal tristate
rlabel metal2 s 18050 49200 18106 50000 6 io_oeb[14]
port 141 nsew signal tristate
rlabel metal2 s 19338 49200 19394 50000 6 io_oeb[15]
port 142 nsew signal tristate
rlabel metal2 s 20534 49200 20590 50000 6 io_oeb[16]
port 143 nsew signal tristate
rlabel metal2 s 21822 49200 21878 50000 6 io_oeb[17]
port 144 nsew signal tristate
rlabel metal2 s 23018 49200 23074 50000 6 io_oeb[18]
port 145 nsew signal tristate
rlabel metal2 s 24306 49200 24362 50000 6 io_oeb[19]
port 146 nsew signal tristate
rlabel metal2 s 1858 49200 1914 50000 6 io_oeb[1]
port 147 nsew signal tristate
rlabel metal2 s 25594 49200 25650 50000 6 io_oeb[20]
port 148 nsew signal tristate
rlabel metal2 s 26790 49200 26846 50000 6 io_oeb[21]
port 149 nsew signal tristate
rlabel metal2 s 28078 49200 28134 50000 6 io_oeb[22]
port 150 nsew signal tristate
rlabel metal2 s 29274 49200 29330 50000 6 io_oeb[23]
port 151 nsew signal tristate
rlabel metal2 s 30562 49200 30618 50000 6 io_oeb[24]
port 152 nsew signal tristate
rlabel metal2 s 31758 49200 31814 50000 6 io_oeb[25]
port 153 nsew signal tristate
rlabel metal2 s 33046 49200 33102 50000 6 io_oeb[26]
port 154 nsew signal tristate
rlabel metal2 s 34334 49200 34390 50000 6 io_oeb[27]
port 155 nsew signal tristate
rlabel metal2 s 35530 49200 35586 50000 6 io_oeb[28]
port 156 nsew signal tristate
rlabel metal2 s 36818 49200 36874 50000 6 io_oeb[29]
port 157 nsew signal tristate
rlabel metal2 s 3054 49200 3110 50000 6 io_oeb[2]
port 158 nsew signal tristate
rlabel metal2 s 38014 49200 38070 50000 6 io_oeb[30]
port 159 nsew signal tristate
rlabel metal2 s 39302 49200 39358 50000 6 io_oeb[31]
port 160 nsew signal tristate
rlabel metal2 s 40498 49200 40554 50000 6 io_oeb[32]
port 161 nsew signal tristate
rlabel metal2 s 41786 49200 41842 50000 6 io_oeb[33]
port 162 nsew signal tristate
rlabel metal2 s 43074 49200 43130 50000 6 io_oeb[34]
port 163 nsew signal tristate
rlabel metal2 s 44270 49200 44326 50000 6 io_oeb[35]
port 164 nsew signal tristate
rlabel metal2 s 45558 49200 45614 50000 6 io_oeb[36]
port 165 nsew signal tristate
rlabel metal2 s 46754 49200 46810 50000 6 io_oeb[37]
port 166 nsew signal tristate
rlabel metal2 s 4342 49200 4398 50000 6 io_oeb[3]
port 167 nsew signal tristate
rlabel metal2 s 5538 49200 5594 50000 6 io_oeb[4]
port 168 nsew signal tristate
rlabel metal2 s 6826 49200 6882 50000 6 io_oeb[5]
port 169 nsew signal tristate
rlabel metal2 s 8022 49200 8078 50000 6 io_oeb[6]
port 170 nsew signal tristate
rlabel metal2 s 9310 49200 9366 50000 6 io_oeb[7]
port 171 nsew signal tristate
rlabel metal2 s 10598 49200 10654 50000 6 io_oeb[8]
port 172 nsew signal tristate
rlabel metal2 s 11794 49200 11850 50000 6 io_oeb[9]
port 173 nsew signal tristate
rlabel metal2 s 1030 49200 1086 50000 6 io_out[0]
port 174 nsew signal tristate
rlabel metal2 s 13450 49200 13506 50000 6 io_out[10]
port 175 nsew signal tristate
rlabel metal2 s 14738 49200 14794 50000 6 io_out[11]
port 176 nsew signal tristate
rlabel metal2 s 15934 49200 15990 50000 6 io_out[12]
port 177 nsew signal tristate
rlabel metal2 s 17222 49200 17278 50000 6 io_out[13]
port 178 nsew signal tristate
rlabel metal2 s 18510 49200 18566 50000 6 io_out[14]
port 179 nsew signal tristate
rlabel metal2 s 19706 49200 19762 50000 6 io_out[15]
port 180 nsew signal tristate
rlabel metal2 s 20994 49200 21050 50000 6 io_out[16]
port 181 nsew signal tristate
rlabel metal2 s 22190 49200 22246 50000 6 io_out[17]
port 182 nsew signal tristate
rlabel metal2 s 23478 49200 23534 50000 6 io_out[18]
port 183 nsew signal tristate
rlabel metal2 s 24674 49200 24730 50000 6 io_out[19]
port 184 nsew signal tristate
rlabel metal2 s 2226 49200 2282 50000 6 io_out[1]
port 185 nsew signal tristate
rlabel metal2 s 25962 49200 26018 50000 6 io_out[20]
port 186 nsew signal tristate
rlabel metal2 s 27250 49200 27306 50000 6 io_out[21]
port 187 nsew signal tristate
rlabel metal2 s 28446 49200 28502 50000 6 io_out[22]
port 188 nsew signal tristate
rlabel metal2 s 29734 49200 29790 50000 6 io_out[23]
port 189 nsew signal tristate
rlabel metal2 s 30930 49200 30986 50000 6 io_out[24]
port 190 nsew signal tristate
rlabel metal2 s 32218 49200 32274 50000 6 io_out[25]
port 191 nsew signal tristate
rlabel metal2 s 33506 49200 33562 50000 6 io_out[26]
port 192 nsew signal tristate
rlabel metal2 s 34702 49200 34758 50000 6 io_out[27]
port 193 nsew signal tristate
rlabel metal2 s 35990 49200 36046 50000 6 io_out[28]
port 194 nsew signal tristate
rlabel metal2 s 37186 49200 37242 50000 6 io_out[29]
port 195 nsew signal tristate
rlabel metal2 s 3514 49200 3570 50000 6 io_out[2]
port 196 nsew signal tristate
rlabel metal2 s 38474 49200 38530 50000 6 io_out[30]
port 197 nsew signal tristate
rlabel metal2 s 39670 49200 39726 50000 6 io_out[31]
port 198 nsew signal tristate
rlabel metal2 s 40958 49200 41014 50000 6 io_out[32]
port 199 nsew signal tristate
rlabel metal2 s 42246 49200 42302 50000 6 io_out[33]
port 200 nsew signal tristate
rlabel metal2 s 43442 49200 43498 50000 6 io_out[34]
port 201 nsew signal tristate
rlabel metal2 s 44730 49200 44786 50000 6 io_out[35]
port 202 nsew signal tristate
rlabel metal2 s 45926 49200 45982 50000 6 io_out[36]
port 203 nsew signal tristate
rlabel metal2 s 47214 49200 47270 50000 6 io_out[37]
port 204 nsew signal tristate
rlabel metal2 s 4710 49200 4766 50000 6 io_out[3]
port 205 nsew signal tristate
rlabel metal2 s 5998 49200 6054 50000 6 io_out[4]
port 206 nsew signal tristate
rlabel metal2 s 7194 49200 7250 50000 6 io_out[5]
port 207 nsew signal tristate
rlabel metal2 s 8482 49200 8538 50000 6 io_out[6]
port 208 nsew signal tristate
rlabel metal2 s 9770 49200 9826 50000 6 io_out[7]
port 209 nsew signal tristate
rlabel metal2 s 10966 49200 11022 50000 6 io_out[8]
port 210 nsew signal tristate
rlabel metal2 s 12254 49200 12310 50000 6 io_out[9]
port 211 nsew signal tristate
rlabel metal2 s 48962 0 49018 800 6 irq[0]
port 212 nsew signal tristate
rlabel metal2 s 49054 0 49110 800 6 irq[1]
port 213 nsew signal tristate
rlabel metal2 s 49146 0 49202 800 6 irq[2]
port 214 nsew signal tristate
rlabel metal2 s 10598 0 10654 800 6 la_data_in[0]
port 215 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[100]
port 216 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[101]
port 217 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[102]
port 218 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[103]
port 219 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[104]
port 220 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_data_in[105]
port 221 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[106]
port 222 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_data_in[107]
port 223 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_data_in[108]
port 224 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_data_in[109]
port 225 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 la_data_in[10]
port 226 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[110]
port 227 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_data_in[111]
port 228 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[112]
port 229 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[113]
port 230 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[114]
port 231 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[115]
port 232 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_data_in[116]
port 233 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[117]
port 234 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_data_in[118]
port 235 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_data_in[119]
port 236 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 la_data_in[11]
port 237 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[120]
port 238 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[121]
port 239 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_data_in[122]
port 240 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_data_in[123]
port 241 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[124]
port 242 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[125]
port 243 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[126]
port 244 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[127]
port 245 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 la_data_in[12]
port 246 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 la_data_in[13]
port 247 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 la_data_in[14]
port 248 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 la_data_in[15]
port 249 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 la_data_in[16]
port 250 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 la_data_in[17]
port 251 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 la_data_in[18]
port 252 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 la_data_in[19]
port 253 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 la_data_in[1]
port 254 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 la_data_in[20]
port 255 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 la_data_in[21]
port 256 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 la_data_in[22]
port 257 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 la_data_in[23]
port 258 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 la_data_in[24]
port 259 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 la_data_in[25]
port 260 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 la_data_in[26]
port 261 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 la_data_in[27]
port 262 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 la_data_in[28]
port 263 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 la_data_in[29]
port 264 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 la_data_in[2]
port 265 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 la_data_in[30]
port 266 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 la_data_in[31]
port 267 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 la_data_in[32]
port 268 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 la_data_in[33]
port 269 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 la_data_in[34]
port 270 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 la_data_in[35]
port 271 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 la_data_in[36]
port 272 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_data_in[37]
port 273 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 la_data_in[38]
port 274 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 la_data_in[39]
port 275 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 la_data_in[3]
port 276 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_data_in[40]
port 277 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 la_data_in[41]
port 278 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 la_data_in[42]
port 279 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[43]
port 280 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 la_data_in[44]
port 281 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_data_in[45]
port 282 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 la_data_in[46]
port 283 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 la_data_in[47]
port 284 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 la_data_in[48]
port 285 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[49]
port 286 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 la_data_in[4]
port 287 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 la_data_in[50]
port 288 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_data_in[51]
port 289 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 la_data_in[52]
port 290 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_data_in[53]
port 291 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_data_in[54]
port 292 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[55]
port 293 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_data_in[56]
port 294 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[57]
port 295 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 la_data_in[58]
port 296 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 la_data_in[59]
port 297 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 la_data_in[5]
port 298 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 la_data_in[60]
port 299 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 la_data_in[61]
port 300 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 la_data_in[62]
port 301 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 la_data_in[63]
port 302 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_data_in[64]
port 303 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_data_in[65]
port 304 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 la_data_in[66]
port 305 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_data_in[67]
port 306 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_data_in[68]
port 307 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_data_in[69]
port 308 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 la_data_in[6]
port 309 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_data_in[70]
port 310 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_data_in[71]
port 311 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_data_in[72]
port 312 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_data_in[73]
port 313 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 la_data_in[74]
port 314 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 la_data_in[75]
port 315 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_data_in[76]
port 316 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in[77]
port 317 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_data_in[78]
port 318 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_data_in[79]
port 319 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 la_data_in[7]
port 320 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[80]
port 321 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_data_in[81]
port 322 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 la_data_in[82]
port 323 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[83]
port 324 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 la_data_in[84]
port 325 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_data_in[85]
port 326 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_data_in[86]
port 327 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_data_in[87]
port 328 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_data_in[88]
port 329 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_data_in[89]
port 330 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 la_data_in[8]
port 331 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_data_in[90]
port 332 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_data_in[91]
port 333 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[92]
port 334 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_data_in[93]
port 335 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_data_in[94]
port 336 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_data_in[95]
port 337 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_in[96]
port 338 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[97]
port 339 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[98]
port 340 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[99]
port 341 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 la_data_in[9]
port 342 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 la_data_out[0]
port 343 nsew signal tristate
rlabel metal2 s 40682 0 40738 800 6 la_data_out[100]
port 344 nsew signal tristate
rlabel metal2 s 40958 0 41014 800 6 la_data_out[101]
port 345 nsew signal tristate
rlabel metal2 s 41234 0 41290 800 6 la_data_out[102]
port 346 nsew signal tristate
rlabel metal2 s 41510 0 41566 800 6 la_data_out[103]
port 347 nsew signal tristate
rlabel metal2 s 41878 0 41934 800 6 la_data_out[104]
port 348 nsew signal tristate
rlabel metal2 s 42154 0 42210 800 6 la_data_out[105]
port 349 nsew signal tristate
rlabel metal2 s 42430 0 42486 800 6 la_data_out[106]
port 350 nsew signal tristate
rlabel metal2 s 42706 0 42762 800 6 la_data_out[107]
port 351 nsew signal tristate
rlabel metal2 s 43074 0 43130 800 6 la_data_out[108]
port 352 nsew signal tristate
rlabel metal2 s 43350 0 43406 800 6 la_data_out[109]
port 353 nsew signal tristate
rlabel metal2 s 13634 0 13690 800 6 la_data_out[10]
port 354 nsew signal tristate
rlabel metal2 s 43626 0 43682 800 6 la_data_out[110]
port 355 nsew signal tristate
rlabel metal2 s 43902 0 43958 800 6 la_data_out[111]
port 356 nsew signal tristate
rlabel metal2 s 44270 0 44326 800 6 la_data_out[112]
port 357 nsew signal tristate
rlabel metal2 s 44546 0 44602 800 6 la_data_out[113]
port 358 nsew signal tristate
rlabel metal2 s 44822 0 44878 800 6 la_data_out[114]
port 359 nsew signal tristate
rlabel metal2 s 45098 0 45154 800 6 la_data_out[115]
port 360 nsew signal tristate
rlabel metal2 s 45466 0 45522 800 6 la_data_out[116]
port 361 nsew signal tristate
rlabel metal2 s 45742 0 45798 800 6 la_data_out[117]
port 362 nsew signal tristate
rlabel metal2 s 46018 0 46074 800 6 la_data_out[118]
port 363 nsew signal tristate
rlabel metal2 s 46294 0 46350 800 6 la_data_out[119]
port 364 nsew signal tristate
rlabel metal2 s 14002 0 14058 800 6 la_data_out[11]
port 365 nsew signal tristate
rlabel metal2 s 46662 0 46718 800 6 la_data_out[120]
port 366 nsew signal tristate
rlabel metal2 s 46938 0 46994 800 6 la_data_out[121]
port 367 nsew signal tristate
rlabel metal2 s 47214 0 47270 800 6 la_data_out[122]
port 368 nsew signal tristate
rlabel metal2 s 47490 0 47546 800 6 la_data_out[123]
port 369 nsew signal tristate
rlabel metal2 s 47858 0 47914 800 6 la_data_out[124]
port 370 nsew signal tristate
rlabel metal2 s 48134 0 48190 800 6 la_data_out[125]
port 371 nsew signal tristate
rlabel metal2 s 48410 0 48466 800 6 la_data_out[126]
port 372 nsew signal tristate
rlabel metal2 s 48686 0 48742 800 6 la_data_out[127]
port 373 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 la_data_out[12]
port 374 nsew signal tristate
rlabel metal2 s 14554 0 14610 800 6 la_data_out[13]
port 375 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 la_data_out[14]
port 376 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 la_data_out[15]
port 377 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 la_data_out[16]
port 378 nsew signal tristate
rlabel metal2 s 15750 0 15806 800 6 la_data_out[17]
port 379 nsew signal tristate
rlabel metal2 s 16026 0 16082 800 6 la_data_out[18]
port 380 nsew signal tristate
rlabel metal2 s 16394 0 16450 800 6 la_data_out[19]
port 381 nsew signal tristate
rlabel metal2 s 10966 0 11022 800 6 la_data_out[1]
port 382 nsew signal tristate
rlabel metal2 s 16670 0 16726 800 6 la_data_out[20]
port 383 nsew signal tristate
rlabel metal2 s 16946 0 17002 800 6 la_data_out[21]
port 384 nsew signal tristate
rlabel metal2 s 17222 0 17278 800 6 la_data_out[22]
port 385 nsew signal tristate
rlabel metal2 s 17590 0 17646 800 6 la_data_out[23]
port 386 nsew signal tristate
rlabel metal2 s 17866 0 17922 800 6 la_data_out[24]
port 387 nsew signal tristate
rlabel metal2 s 18142 0 18198 800 6 la_data_out[25]
port 388 nsew signal tristate
rlabel metal2 s 18418 0 18474 800 6 la_data_out[26]
port 389 nsew signal tristate
rlabel metal2 s 18786 0 18842 800 6 la_data_out[27]
port 390 nsew signal tristate
rlabel metal2 s 19062 0 19118 800 6 la_data_out[28]
port 391 nsew signal tristate
rlabel metal2 s 19338 0 19394 800 6 la_data_out[29]
port 392 nsew signal tristate
rlabel metal2 s 11242 0 11298 800 6 la_data_out[2]
port 393 nsew signal tristate
rlabel metal2 s 19614 0 19670 800 6 la_data_out[30]
port 394 nsew signal tristate
rlabel metal2 s 19982 0 20038 800 6 la_data_out[31]
port 395 nsew signal tristate
rlabel metal2 s 20258 0 20314 800 6 la_data_out[32]
port 396 nsew signal tristate
rlabel metal2 s 20534 0 20590 800 6 la_data_out[33]
port 397 nsew signal tristate
rlabel metal2 s 20810 0 20866 800 6 la_data_out[34]
port 398 nsew signal tristate
rlabel metal2 s 21178 0 21234 800 6 la_data_out[35]
port 399 nsew signal tristate
rlabel metal2 s 21454 0 21510 800 6 la_data_out[36]
port 400 nsew signal tristate
rlabel metal2 s 21730 0 21786 800 6 la_data_out[37]
port 401 nsew signal tristate
rlabel metal2 s 22098 0 22154 800 6 la_data_out[38]
port 402 nsew signal tristate
rlabel metal2 s 22374 0 22430 800 6 la_data_out[39]
port 403 nsew signal tristate
rlabel metal2 s 11518 0 11574 800 6 la_data_out[3]
port 404 nsew signal tristate
rlabel metal2 s 22650 0 22706 800 6 la_data_out[40]
port 405 nsew signal tristate
rlabel metal2 s 22926 0 22982 800 6 la_data_out[41]
port 406 nsew signal tristate
rlabel metal2 s 23294 0 23350 800 6 la_data_out[42]
port 407 nsew signal tristate
rlabel metal2 s 23570 0 23626 800 6 la_data_out[43]
port 408 nsew signal tristate
rlabel metal2 s 23846 0 23902 800 6 la_data_out[44]
port 409 nsew signal tristate
rlabel metal2 s 24122 0 24178 800 6 la_data_out[45]
port 410 nsew signal tristate
rlabel metal2 s 24490 0 24546 800 6 la_data_out[46]
port 411 nsew signal tristate
rlabel metal2 s 24766 0 24822 800 6 la_data_out[47]
port 412 nsew signal tristate
rlabel metal2 s 25042 0 25098 800 6 la_data_out[48]
port 413 nsew signal tristate
rlabel metal2 s 25318 0 25374 800 6 la_data_out[49]
port 414 nsew signal tristate
rlabel metal2 s 11886 0 11942 800 6 la_data_out[4]
port 415 nsew signal tristate
rlabel metal2 s 25686 0 25742 800 6 la_data_out[50]
port 416 nsew signal tristate
rlabel metal2 s 25962 0 26018 800 6 la_data_out[51]
port 417 nsew signal tristate
rlabel metal2 s 26238 0 26294 800 6 la_data_out[52]
port 418 nsew signal tristate
rlabel metal2 s 26514 0 26570 800 6 la_data_out[53]
port 419 nsew signal tristate
rlabel metal2 s 26882 0 26938 800 6 la_data_out[54]
port 420 nsew signal tristate
rlabel metal2 s 27158 0 27214 800 6 la_data_out[55]
port 421 nsew signal tristate
rlabel metal2 s 27434 0 27490 800 6 la_data_out[56]
port 422 nsew signal tristate
rlabel metal2 s 27710 0 27766 800 6 la_data_out[57]
port 423 nsew signal tristate
rlabel metal2 s 28078 0 28134 800 6 la_data_out[58]
port 424 nsew signal tristate
rlabel metal2 s 28354 0 28410 800 6 la_data_out[59]
port 425 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 la_data_out[5]
port 426 nsew signal tristate
rlabel metal2 s 28630 0 28686 800 6 la_data_out[60]
port 427 nsew signal tristate
rlabel metal2 s 28906 0 28962 800 6 la_data_out[61]
port 428 nsew signal tristate
rlabel metal2 s 29274 0 29330 800 6 la_data_out[62]
port 429 nsew signal tristate
rlabel metal2 s 29550 0 29606 800 6 la_data_out[63]
port 430 nsew signal tristate
rlabel metal2 s 29826 0 29882 800 6 la_data_out[64]
port 431 nsew signal tristate
rlabel metal2 s 30102 0 30158 800 6 la_data_out[65]
port 432 nsew signal tristate
rlabel metal2 s 30470 0 30526 800 6 la_data_out[66]
port 433 nsew signal tristate
rlabel metal2 s 30746 0 30802 800 6 la_data_out[67]
port 434 nsew signal tristate
rlabel metal2 s 31022 0 31078 800 6 la_data_out[68]
port 435 nsew signal tristate
rlabel metal2 s 31390 0 31446 800 6 la_data_out[69]
port 436 nsew signal tristate
rlabel metal2 s 12438 0 12494 800 6 la_data_out[6]
port 437 nsew signal tristate
rlabel metal2 s 31666 0 31722 800 6 la_data_out[70]
port 438 nsew signal tristate
rlabel metal2 s 31942 0 31998 800 6 la_data_out[71]
port 439 nsew signal tristate
rlabel metal2 s 32218 0 32274 800 6 la_data_out[72]
port 440 nsew signal tristate
rlabel metal2 s 32586 0 32642 800 6 la_data_out[73]
port 441 nsew signal tristate
rlabel metal2 s 32862 0 32918 800 6 la_data_out[74]
port 442 nsew signal tristate
rlabel metal2 s 33138 0 33194 800 6 la_data_out[75]
port 443 nsew signal tristate
rlabel metal2 s 33414 0 33470 800 6 la_data_out[76]
port 444 nsew signal tristate
rlabel metal2 s 33782 0 33838 800 6 la_data_out[77]
port 445 nsew signal tristate
rlabel metal2 s 34058 0 34114 800 6 la_data_out[78]
port 446 nsew signal tristate
rlabel metal2 s 34334 0 34390 800 6 la_data_out[79]
port 447 nsew signal tristate
rlabel metal2 s 12806 0 12862 800 6 la_data_out[7]
port 448 nsew signal tristate
rlabel metal2 s 34610 0 34666 800 6 la_data_out[80]
port 449 nsew signal tristate
rlabel metal2 s 34978 0 35034 800 6 la_data_out[81]
port 450 nsew signal tristate
rlabel metal2 s 35254 0 35310 800 6 la_data_out[82]
port 451 nsew signal tristate
rlabel metal2 s 35530 0 35586 800 6 la_data_out[83]
port 452 nsew signal tristate
rlabel metal2 s 35806 0 35862 800 6 la_data_out[84]
port 453 nsew signal tristate
rlabel metal2 s 36174 0 36230 800 6 la_data_out[85]
port 454 nsew signal tristate
rlabel metal2 s 36450 0 36506 800 6 la_data_out[86]
port 455 nsew signal tristate
rlabel metal2 s 36726 0 36782 800 6 la_data_out[87]
port 456 nsew signal tristate
rlabel metal2 s 37002 0 37058 800 6 la_data_out[88]
port 457 nsew signal tristate
rlabel metal2 s 37370 0 37426 800 6 la_data_out[89]
port 458 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 la_data_out[8]
port 459 nsew signal tristate
rlabel metal2 s 37646 0 37702 800 6 la_data_out[90]
port 460 nsew signal tristate
rlabel metal2 s 37922 0 37978 800 6 la_data_out[91]
port 461 nsew signal tristate
rlabel metal2 s 38198 0 38254 800 6 la_data_out[92]
port 462 nsew signal tristate
rlabel metal2 s 38566 0 38622 800 6 la_data_out[93]
port 463 nsew signal tristate
rlabel metal2 s 38842 0 38898 800 6 la_data_out[94]
port 464 nsew signal tristate
rlabel metal2 s 39118 0 39174 800 6 la_data_out[95]
port 465 nsew signal tristate
rlabel metal2 s 39394 0 39450 800 6 la_data_out[96]
port 466 nsew signal tristate
rlabel metal2 s 39762 0 39818 800 6 la_data_out[97]
port 467 nsew signal tristate
rlabel metal2 s 40038 0 40094 800 6 la_data_out[98]
port 468 nsew signal tristate
rlabel metal2 s 40314 0 40370 800 6 la_data_out[99]
port 469 nsew signal tristate
rlabel metal2 s 13358 0 13414 800 6 la_data_out[9]
port 470 nsew signal tristate
rlabel metal2 s 10782 0 10838 800 6 la_oenb[0]
port 471 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_oenb[100]
port 472 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_oenb[101]
port 473 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_oenb[102]
port 474 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_oenb[103]
port 475 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_oenb[104]
port 476 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_oenb[105]
port 477 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_oenb[106]
port 478 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_oenb[107]
port 479 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[108]
port 480 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_oenb[109]
port 481 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 la_oenb[10]
port 482 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_oenb[110]
port 483 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_oenb[111]
port 484 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_oenb[112]
port 485 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_oenb[113]
port 486 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_oenb[114]
port 487 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[115]
port 488 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_oenb[116]
port 489 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[117]
port 490 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_oenb[118]
port 491 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[119]
port 492 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 la_oenb[11]
port 493 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_oenb[120]
port 494 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[121]
port 495 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_oenb[122]
port 496 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_oenb[123]
port 497 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_oenb[124]
port 498 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[125]
port 499 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[126]
port 500 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[127]
port 501 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 la_oenb[12]
port 502 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 la_oenb[13]
port 503 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 la_oenb[14]
port 504 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 la_oenb[15]
port 505 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 la_oenb[16]
port 506 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 la_oenb[17]
port 507 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_oenb[18]
port 508 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 la_oenb[19]
port 509 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 la_oenb[1]
port 510 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 la_oenb[20]
port 511 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 la_oenb[21]
port 512 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 la_oenb[22]
port 513 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 la_oenb[23]
port 514 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 la_oenb[24]
port 515 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 la_oenb[25]
port 516 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 la_oenb[26]
port 517 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 la_oenb[27]
port 518 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 la_oenb[28]
port 519 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 la_oenb[29]
port 520 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 la_oenb[2]
port 521 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 la_oenb[30]
port 522 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 la_oenb[31]
port 523 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 la_oenb[32]
port 524 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 la_oenb[33]
port 525 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 la_oenb[34]
port 526 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_oenb[35]
port 527 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 la_oenb[36]
port 528 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_oenb[37]
port 529 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_oenb[38]
port 530 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 la_oenb[39]
port 531 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 la_oenb[3]
port 532 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 la_oenb[40]
port 533 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 la_oenb[41]
port 534 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 la_oenb[42]
port 535 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 la_oenb[43]
port 536 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_oenb[44]
port 537 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 la_oenb[45]
port 538 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_oenb[46]
port 539 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 la_oenb[47]
port 540 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_oenb[48]
port 541 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 la_oenb[49]
port 542 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 la_oenb[4]
port 543 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_oenb[50]
port 544 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 la_oenb[51]
port 545 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_oenb[52]
port 546 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 la_oenb[53]
port 547 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_oenb[54]
port 548 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 la_oenb[55]
port 549 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_oenb[56]
port 550 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 la_oenb[57]
port 551 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_oenb[58]
port 552 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_oenb[59]
port 553 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_oenb[5]
port 554 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_oenb[60]
port 555 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 la_oenb[61]
port 556 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_oenb[62]
port 557 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la_oenb[63]
port 558 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[64]
port 559 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_oenb[65]
port 560 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_oenb[66]
port 561 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 la_oenb[67]
port 562 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_oenb[68]
port 563 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 la_oenb[69]
port 564 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 la_oenb[6]
port 565 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_oenb[70]
port 566 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 la_oenb[71]
port 567 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_oenb[72]
port 568 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_oenb[73]
port 569 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_oenb[74]
port 570 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_oenb[75]
port 571 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_oenb[76]
port 572 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 la_oenb[77]
port 573 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_oenb[78]
port 574 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_oenb[79]
port 575 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 la_oenb[7]
port 576 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_oenb[80]
port 577 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_oenb[81]
port 578 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_oenb[82]
port 579 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_oenb[83]
port 580 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_oenb[84]
port 581 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_oenb[85]
port 582 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[86]
port 583 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_oenb[87]
port 584 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_oenb[88]
port 585 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_oenb[89]
port 586 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 la_oenb[8]
port 587 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_oenb[90]
port 588 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_oenb[91]
port 589 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_oenb[92]
port 590 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_oenb[93]
port 591 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_oenb[94]
port 592 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_oenb[95]
port 593 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_oenb[96]
port 594 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_oenb[97]
port 595 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 la_oenb[98]
port 596 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[99]
port 597 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 la_oenb[9]
port 598 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 599 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 599 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 600 nsew ground input
rlabel metal2 s 18 0 74 800 6 wb_clk_i
port 601 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_rst_i
port 602 nsew signal input
rlabel metal2 s 202 0 258 800 6 wbs_ack_o
port 603 nsew signal tristate
rlabel metal2 s 570 0 626 800 6 wbs_adr_i[0]
port 604 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_adr_i[10]
port 605 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[11]
port 606 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[12]
port 607 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_adr_i[13]
port 608 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[14]
port 609 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[15]
port 610 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[16]
port 611 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_adr_i[17]
port 612 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[18]
port 613 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[19]
port 614 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_adr_i[1]
port 615 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_adr_i[20]
port 616 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wbs_adr_i[21]
port 617 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[22]
port 618 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_adr_i[23]
port 619 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[24]
port 620 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[25]
port 621 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[26]
port 622 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[27]
port 623 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[28]
port 624 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_adr_i[29]
port 625 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_adr_i[2]
port 626 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[30]
port 627 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[31]
port 628 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_adr_i[3]
port 629 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[4]
port 630 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_adr_i[5]
port 631 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_adr_i[6]
port 632 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_adr_i[7]
port 633 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_adr_i[8]
port 634 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[9]
port 635 nsew signal input
rlabel metal2 s 294 0 350 800 6 wbs_cyc_i
port 636 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_dat_i[0]
port 637 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[10]
port 638 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_i[11]
port 639 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[12]
port 640 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_i[13]
port 641 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_i[14]
port 642 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[15]
port 643 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[16]
port 644 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_i[17]
port 645 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_i[18]
port 646 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[19]
port 647 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_dat_i[1]
port 648 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[20]
port 649 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_i[21]
port 650 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_i[22]
port 651 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_i[23]
port 652 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[24]
port 653 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_i[25]
port 654 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_i[26]
port 655 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_i[27]
port 656 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[28]
port 657 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_i[29]
port 658 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[2]
port 659 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_i[30]
port 660 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_i[31]
port 661 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_dat_i[3]
port 662 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_dat_i[4]
port 663 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[5]
port 664 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_dat_i[6]
port 665 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_i[7]
port 666 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_dat_i[8]
port 667 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_dat_i[9]
port 668 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_dat_o[0]
port 669 nsew signal tristate
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_o[10]
port 670 nsew signal tristate
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[11]
port 671 nsew signal tristate
rlabel metal2 s 4802 0 4858 800 6 wbs_dat_o[12]
port 672 nsew signal tristate
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[13]
port 673 nsew signal tristate
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_o[14]
port 674 nsew signal tristate
rlabel metal2 s 5630 0 5686 800 6 wbs_dat_o[15]
port 675 nsew signal tristate
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_o[16]
port 676 nsew signal tristate
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_o[17]
port 677 nsew signal tristate
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[18]
port 678 nsew signal tristate
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_o[19]
port 679 nsew signal tristate
rlabel metal2 s 1214 0 1270 800 6 wbs_dat_o[1]
port 680 nsew signal tristate
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[20]
port 681 nsew signal tristate
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_o[21]
port 682 nsew signal tristate
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_o[22]
port 683 nsew signal tristate
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[23]
port 684 nsew signal tristate
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_o[24]
port 685 nsew signal tristate
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[25]
port 686 nsew signal tristate
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_o[26]
port 687 nsew signal tristate
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[27]
port 688 nsew signal tristate
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[28]
port 689 nsew signal tristate
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[29]
port 690 nsew signal tristate
rlabel metal2 s 1582 0 1638 800 6 wbs_dat_o[2]
port 691 nsew signal tristate
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[30]
port 692 nsew signal tristate
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_o[31]
port 693 nsew signal tristate
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_o[3]
port 694 nsew signal tristate
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_o[4]
port 695 nsew signal tristate
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_o[5]
port 696 nsew signal tristate
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[6]
port 697 nsew signal tristate
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_o[7]
port 698 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_o[8]
port 699 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[9]
port 700 nsew signal tristate
rlabel metal2 s 846 0 902 800 6 wbs_sel_i[0]
port 701 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_sel_i[1]
port 702 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_sel_i[2]
port 703 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_sel_i[3]
port 704 nsew signal input
rlabel metal2 s 386 0 442 800 6 wbs_stb_i
port 705 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_we_i
port 706 nsew signal input
rlabel metal3 s 49200 42440 50000 42560 6 web0
port 707 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
